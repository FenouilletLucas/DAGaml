// Benchmark "dalu" written by ABC on Tue May 16 16:07:48 2017

module dalu ( 
    inA0, inA1, inA2, inA3, inA4, inA5, inA6, inA7, inA8, inA9, inB0, inB1,
    inB2, inB3, inB4, inB5, inB6, inB7, inB8, inB9, inC0, inC1, inC2, inC3,
    inC4, inC5, inC6, inC7, inC8, inC9, inD0, inD1, inD2, inD3, inD4, inD5,
    inD6, inD7, inD8, inD9, inA10, inA11, inA12, inA13, inA14, inA15,
    inB10, inB11, inB12, inB13, inB14, inB15, inC10, inC11, inC12, inC13,
    inC14, inC15, inD10, inD11, inD12, inD13, inD14, inD15, musel1, musel2,
    musel3, musel4, sh0, sh1, sh2, opsel0, opsel1, opsel2, opsel3,
    O10, O11, O12, O13, O14, O15, O0, O1, O2, O3, O4, O5, O6, O7, O8, O9  );
  input  inA0, inA1, inA2, inA3, inA4, inA5, inA6, inA7, inA8, inA9,
    inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7, inB8, inB9, inC0, inC1,
    inC2, inC3, inC4, inC5, inC6, inC7, inC8, inC9, inD0, inD1, inD2, inD3,
    inD4, inD5, inD6, inD7, inD8, inD9, inA10, inA11, inA12, inA13, inA14,
    inA15, inB10, inB11, inB12, inB13, inB14, inB15, inC10, inC11, inC12,
    inC13, inC14, inC15, inD10, inD11, inD12, inD13, inD14, inD15, musel1,
    musel2, musel3, musel4, sh0, sh1, sh2, opsel0, opsel1, opsel2, opsel3;
  output O10, O11, O12, O13, O14, O15, O0, O1, O2, O3, O4, O5, O6, O7, O8, O9;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
  assign n92 = ~sh0 & sh2;
  assign n93 = ~sh1 & n92;
  assign n94 = ~opsel0 & ~opsel1;
  assign n95 = ~opsel2 & opsel3;
  assign n96 = ~opsel1 & n95;
  assign n97 = opsel2 & ~opsel3;
  assign n98 = ~n94 & n97;
  assign n99 = n94 & n96;
  assign n100 = ~n98 & ~n99;
  assign n101 = musel1 & ~musel2;
  assign n102 = musel3 & ~musel4;
  assign n103 = ~musel1 & musel2;
  assign n104 = n102 & n103;
  assign n105 = n101 & n102;
  assign n106 = ~n104 & ~n105;
  assign n107 = musel2 & n102;
  assign n108 = ~musel1 & ~musel2;
  assign n109 = ~musel3 & musel4;
  assign n110 = n108 & n109;
  assign n111 = musel1 & n107;
  assign n112 = ~n110 & ~n111;
  assign n113 = inB14 & ~n106;
  assign n114 = inD14 & ~n112;
  assign n115 = ~n113 & ~n114;
  assign n116 = sh0 & sh2;
  assign n117 = sh1 & ~sh2;
  assign n118 = sh0 & ~sh1;
  assign n119 = ~n92 & ~n117;
  assign n120 = ~n118 & n119;
  assign n121 = n116 & ~n120;
  assign n122 = inB15 & ~n106;
  assign n123 = inD15 & ~n112;
  assign n124 = ~n122 & ~n123;
  assign n125 = sh0 & sh1;
  assign n126 = ~n120 & n125;
  assign n127 = inB13 & ~n106;
  assign n128 = inD13 & ~n112;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~sh0 & n117;
  assign n131 = inB12 & ~n106;
  assign n132 = inD12 & ~n112;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~sh1 & ~sh2;
  assign n135 = ~n120 & n134;
  assign n136 = inB11 & ~n106;
  assign n137 = inD11 & ~n112;
  assign n138 = ~n136 & ~n137;
  assign n139 = inB10 & ~n106;
  assign n140 = inD10 & ~n112;
  assign n141 = ~n139 & ~n140;
  assign n142 = sh2 & ~n125;
  assign n143 = sh1 & n142;
  assign n144 = ~n124 & n143;
  assign n145 = ~opsel2 & ~opsel3;
  assign n146 = ~n94 & n145;
  assign n147 = n94 & n97;
  assign n148 = ~n146 & ~n147;
  assign n149 = inA15 & n101;
  assign n150 = inC15 & n103;
  assign n151 = ~n149 & ~n150;
  assign n152 = n109 & ~n151;
  assign n153 = n109 & ~n152;
  assign n154 = inA0 & n101;
  assign n155 = inC0 & n103;
  assign n156 = ~n154 & ~n155;
  assign n157 = n153 & ~n156;
  assign n158 = n152 & n156;
  assign n159 = ~n157 & ~n158;
  assign n160 = n152 & ~n159;
  assign n161 = inA1 & n101;
  assign n162 = inC1 & n103;
  assign n163 = ~n161 & ~n162;
  assign n164 = n153 & ~n163;
  assign n165 = n152 & n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = n160 & ~n166;
  assign n168 = inA2 & n101;
  assign n169 = inC2 & n103;
  assign n170 = ~n168 & ~n169;
  assign n171 = n153 & ~n170;
  assign n172 = n152 & n170;
  assign n173 = ~n171 & ~n172;
  assign n174 = inA3 & n101;
  assign n175 = inC3 & n103;
  assign n176 = ~n174 & ~n175;
  assign n177 = n153 & ~n176;
  assign n178 = n152 & n176;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n173 & ~n179;
  assign n181 = n167 & n180;
  assign n182 = inA8 & n101;
  assign n183 = inC8 & n103;
  assign n184 = ~n182 & ~n183;
  assign n185 = n153 & ~n184;
  assign n186 = n152 & n184;
  assign n187 = ~n185 & ~n186;
  assign n188 = inA9 & n101;
  assign n189 = inC9 & n103;
  assign n190 = ~n188 & ~n189;
  assign n191 = n153 & ~n190;
  assign n192 = n152 & n190;
  assign n193 = ~n191 & ~n192;
  assign n194 = inA10 & n101;
  assign n195 = inC10 & n103;
  assign n196 = ~n194 & ~n195;
  assign n197 = n153 & ~n196;
  assign n198 = n152 & n196;
  assign n199 = ~n197 & ~n198;
  assign n200 = inA11 & n101;
  assign n201 = inC11 & n103;
  assign n202 = ~n200 & ~n201;
  assign n203 = n153 & ~n202;
  assign n204 = n152 & n202;
  assign n205 = ~n203 & ~n204;
  assign n206 = ~n199 & ~n205;
  assign n207 = ~n193 & n206;
  assign n208 = ~n187 & n207;
  assign n209 = n181 & n208;
  assign n210 = ~n199 & ~n209;
  assign n211 = ~n94 & n96;
  assign n212 = ~opsel0 & ~n94;
  assign n213 = n95 & n212;
  assign n214 = ~n211 & ~n213;
  assign n215 = musel1 & n102;
  assign n216 = inC10 & n196;
  assign n217 = n107 & n216;
  assign n218 = inA10 & n104;
  assign n219 = ~n196 & n215;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~n217 & n220;
  assign n222 = inC10 & n110;
  assign n223 = n221 & ~n222;
  assign n224 = musel3 & n108;
  assign n225 = ~musel3 & n103;
  assign n226 = musel1 & ~musel3;
  assign n227 = ~inA10 & ~musel2;
  assign n228 = ~n225 & n227;
  assign n229 = ~n224 & n228;
  assign n230 = ~inC10 & musel2;
  assign n231 = ~n225 & n230;
  assign n232 = ~n224 & n231;
  assign n233 = ~inA10 & ~inB10;
  assign n234 = ~musel2 & n233;
  assign n235 = ~n224 & n234;
  assign n236 = ~inB10 & ~inC10;
  assign n237 = musel2 & n236;
  assign n238 = ~n224 & n237;
  assign n239 = ~inA10 & ~inD10;
  assign n240 = ~musel2 & n239;
  assign n241 = ~n225 & n240;
  assign n242 = ~inC10 & ~inD10;
  assign n243 = musel2 & n242;
  assign n244 = ~n225 & n243;
  assign n245 = ~inD10 & n233;
  assign n246 = ~musel2 & n245;
  assign n247 = ~inD10 & n236;
  assign n248 = musel2 & n247;
  assign n249 = ~n225 & ~n226;
  assign n250 = ~n224 & n249;
  assign n251 = ~inB10 & ~n226;
  assign n252 = ~n224 & n251;
  assign n253 = ~inD10 & ~n226;
  assign n254 = ~n225 & n253;
  assign n255 = ~inB10 & ~inD10;
  assign n256 = ~n226 & n255;
  assign n257 = ~musel4 & ~n256;
  assign n258 = ~n254 & n257;
  assign n259 = ~n252 & n258;
  assign n260 = ~n250 & n259;
  assign n261 = ~n248 & n260;
  assign n262 = ~n246 & n261;
  assign n263 = ~n244 & n262;
  assign n264 = ~n241 & n263;
  assign n265 = ~n238 & n264;
  assign n266 = ~n235 & n265;
  assign n267 = ~n232 & n266;
  assign n268 = ~n229 & n267;
  assign n269 = n223 & ~n268;
  assign n270 = ~n100 & ~n115;
  assign n271 = n93 & n270;
  assign n272 = ~n100 & ~n124;
  assign n273 = n121 & n272;
  assign n274 = ~n100 & ~n129;
  assign n275 = n126 & n274;
  assign n276 = ~n100 & ~n133;
  assign n277 = n130 & n276;
  assign n278 = ~n100 & ~n138;
  assign n279 = n135 & n278;
  assign n280 = n120 & ~n141;
  assign n281 = ~n100 & n280;
  assign n282 = ~n100 & n144;
  assign n283 = ~n148 & n210;
  assign n284 = ~n214 & ~n269;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n282 & n285;
  assign n287 = ~n281 & n286;
  assign n288 = ~n279 & n287;
  assign n289 = ~n277 & n288;
  assign n290 = ~n275 & n289;
  assign n291 = ~n273 & n290;
  assign O10 = n271 | ~n291;
  assign n293 = ~n199 & ~n210;
  assign n294 = inC11 & n202;
  assign n295 = n107 & n294;
  assign n296 = inA11 & n104;
  assign n297 = ~n202 & n215;
  assign n298 = ~n296 & ~n297;
  assign n299 = ~n295 & n298;
  assign n300 = inC11 & n110;
  assign n301 = n299 & ~n300;
  assign n302 = ~inA11 & ~musel2;
  assign n303 = ~n225 & n302;
  assign n304 = ~n224 & n303;
  assign n305 = ~inC11 & musel2;
  assign n306 = ~n225 & n305;
  assign n307 = ~n224 & n306;
  assign n308 = ~inA11 & ~inB11;
  assign n309 = ~musel2 & n308;
  assign n310 = ~n224 & n309;
  assign n311 = ~inB11 & ~inC11;
  assign n312 = musel2 & n311;
  assign n313 = ~n224 & n312;
  assign n314 = ~inA11 & ~inD11;
  assign n315 = ~musel2 & n314;
  assign n316 = ~n225 & n315;
  assign n317 = ~inC11 & ~inD11;
  assign n318 = musel2 & n317;
  assign n319 = ~n225 & n318;
  assign n320 = ~inD11 & n308;
  assign n321 = ~musel2 & n320;
  assign n322 = ~inD11 & n311;
  assign n323 = musel2 & n322;
  assign n324 = ~inB11 & ~n226;
  assign n325 = ~n224 & n324;
  assign n326 = ~inD11 & ~n226;
  assign n327 = ~n225 & n326;
  assign n328 = ~inB11 & ~inD11;
  assign n329 = ~n226 & n328;
  assign n330 = ~musel4 & ~n329;
  assign n331 = ~n327 & n330;
  assign n332 = ~n325 & n331;
  assign n333 = ~n250 & n332;
  assign n334 = ~n323 & n333;
  assign n335 = ~n321 & n334;
  assign n336 = ~n319 & n335;
  assign n337 = ~n316 & n336;
  assign n338 = ~n313 & n337;
  assign n339 = ~n310 & n338;
  assign n340 = ~n307 & n339;
  assign n341 = ~n304 & n340;
  assign n342 = n301 & ~n341;
  assign n343 = ~n148 & ~n205;
  assign n344 = ~n293 & n343;
  assign n345 = n126 & n270;
  assign n346 = n130 & n274;
  assign n347 = n135 & n276;
  assign n348 = n142 & n272;
  assign n349 = n120 & ~n138;
  assign n350 = ~n100 & n349;
  assign n351 = ~n214 & ~n342;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~n348 & n352;
  assign n354 = ~n347 & n353;
  assign n355 = ~n346 & n354;
  assign n356 = ~n345 & n355;
  assign O11 = n344 | ~n356;
  assign n358 = ~n98 & n100;
  assign n359 = n135 & ~n358;
  assign n360 = n120 & ~n358;
  assign n361 = n130 & ~n358;
  assign n362 = inA4 & n101;
  assign n363 = inC4 & n103;
  assign n364 = ~n362 & ~n363;
  assign n365 = n153 & ~n364;
  assign n366 = n152 & n364;
  assign n367 = ~n365 & ~n366;
  assign n368 = inA5 & n101;
  assign n369 = inC5 & n103;
  assign n370 = ~n368 & ~n369;
  assign n371 = n153 & ~n370;
  assign n372 = n152 & n370;
  assign n373 = ~n371 & ~n372;
  assign n374 = inA6 & n101;
  assign n375 = inC6 & n103;
  assign n376 = ~n374 & ~n375;
  assign n377 = n153 & ~n376;
  assign n378 = n152 & n376;
  assign n379 = ~n377 & ~n378;
  assign n380 = inA7 & n101;
  assign n381 = inC7 & n103;
  assign n382 = ~n380 & ~n381;
  assign n383 = n153 & ~n382;
  assign n384 = n152 & n382;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n379 & ~n385;
  assign n387 = ~n373 & n386;
  assign n388 = ~n367 & n387;
  assign n389 = n209 & n388;
  assign n390 = inA12 & n101;
  assign n391 = inC12 & n103;
  assign n392 = ~n390 & ~n391;
  assign n393 = n153 & ~n392;
  assign n394 = n152 & n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = n389 & ~n395;
  assign n397 = ~inA12 & ~musel2;
  assign n398 = ~n225 & n397;
  assign n399 = ~n224 & n398;
  assign n400 = ~inC12 & musel2;
  assign n401 = ~n225 & n400;
  assign n402 = ~n224 & n401;
  assign n403 = ~inA12 & ~inB12;
  assign n404 = ~musel2 & n403;
  assign n405 = ~n224 & n404;
  assign n406 = ~inB12 & ~inC12;
  assign n407 = musel2 & n406;
  assign n408 = ~n224 & n407;
  assign n409 = ~inA12 & ~inD12;
  assign n410 = ~musel2 & n409;
  assign n411 = ~n225 & n410;
  assign n412 = ~inC12 & ~inD12;
  assign n413 = musel2 & n412;
  assign n414 = ~n225 & n413;
  assign n415 = ~inD12 & n403;
  assign n416 = ~musel2 & n415;
  assign n417 = ~inD12 & n406;
  assign n418 = musel2 & n417;
  assign n419 = ~inB12 & ~n226;
  assign n420 = ~n224 & n419;
  assign n421 = ~inD12 & ~n226;
  assign n422 = ~n225 & n421;
  assign n423 = ~inB12 & ~inD12;
  assign n424 = ~n226 & n423;
  assign n425 = ~musel4 & ~n424;
  assign n426 = ~n422 & n425;
  assign n427 = ~n420 & n426;
  assign n428 = ~n250 & n427;
  assign n429 = ~n418 & n428;
  assign n430 = ~n416 & n429;
  assign n431 = ~n414 & n430;
  assign n432 = ~n411 & n431;
  assign n433 = ~n408 & n432;
  assign n434 = ~n405 & n433;
  assign n435 = ~n402 & n434;
  assign n436 = ~n399 & n435;
  assign n437 = inC12 & n392;
  assign n438 = n107 & n437;
  assign n439 = inA12 & n104;
  assign n440 = n215 & ~n392;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n438 & n441;
  assign n443 = inC12 & n110;
  assign n444 = n442 & ~n443;
  assign n445 = ~n124 & ~n358;
  assign n446 = ~n361 & n445;
  assign n447 = ~n360 & n446;
  assign n448 = ~n359 & n447;
  assign n449 = ~n148 & n389;
  assign n450 = ~n396 & n449;
  assign n451 = ~n148 & ~n395;
  assign n452 = ~n396 & n451;
  assign n453 = ~n129 & n359;
  assign n454 = ~n133 & n360;
  assign n455 = ~n115 & n361;
  assign n456 = ~n214 & n436;
  assign n457 = ~n214 & ~n444;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~n455 & n458;
  assign n460 = ~n454 & n459;
  assign n461 = ~n453 & n460;
  assign n462 = ~n452 & n461;
  assign n463 = ~n450 & n462;
  assign O12 = n448 | ~n463;
  assign n465 = ~n100 & n135;
  assign n466 = ~n100 & n120;
  assign n467 = inA13 & n101;
  assign n468 = inC13 & n103;
  assign n469 = ~n467 & ~n468;
  assign n470 = n153 & ~n469;
  assign n471 = n152 & n469;
  assign n472 = ~n470 & ~n471;
  assign n473 = n396 & ~n472;
  assign n474 = ~inA13 & ~musel2;
  assign n475 = ~n225 & n474;
  assign n476 = ~n224 & n475;
  assign n477 = ~inC13 & musel2;
  assign n478 = ~n225 & n477;
  assign n479 = ~n224 & n478;
  assign n480 = ~inA13 & ~inB13;
  assign n481 = ~musel2 & n480;
  assign n482 = ~n224 & n481;
  assign n483 = ~inB13 & ~inC13;
  assign n484 = musel2 & n483;
  assign n485 = ~n224 & n484;
  assign n486 = ~inA13 & ~inD13;
  assign n487 = ~musel2 & n486;
  assign n488 = ~n225 & n487;
  assign n489 = ~inC13 & ~inD13;
  assign n490 = musel2 & n489;
  assign n491 = ~n225 & n490;
  assign n492 = ~inD13 & n480;
  assign n493 = ~musel2 & n492;
  assign n494 = ~inD13 & n483;
  assign n495 = musel2 & n494;
  assign n496 = ~inB13 & ~n226;
  assign n497 = ~n224 & n496;
  assign n498 = ~inD13 & ~n226;
  assign n499 = ~n225 & n498;
  assign n500 = ~inB13 & ~inD13;
  assign n501 = ~n226 & n500;
  assign n502 = ~musel4 & ~n501;
  assign n503 = ~n499 & n502;
  assign n504 = ~n497 & n503;
  assign n505 = ~n250 & n504;
  assign n506 = ~n495 & n505;
  assign n507 = ~n493 & n506;
  assign n508 = ~n491 & n507;
  assign n509 = ~n488 & n508;
  assign n510 = ~n485 & n509;
  assign n511 = ~n482 & n510;
  assign n512 = ~n479 & n511;
  assign n513 = ~n476 & n512;
  assign n514 = inC13 & n469;
  assign n515 = n107 & n514;
  assign n516 = inA13 & n104;
  assign n517 = n215 & ~n469;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n515 & n518;
  assign n520 = inC13 & n110;
  assign n521 = n519 & ~n520;
  assign n522 = ~n513 & n521;
  assign n523 = n272 & ~n466;
  assign n524 = ~n465 & n523;
  assign n525 = ~n148 & n396;
  assign n526 = ~n473 & n525;
  assign n527 = ~n148 & ~n472;
  assign n528 = ~n473 & n527;
  assign n529 = ~n115 & n465;
  assign n530 = ~n129 & n466;
  assign n531 = ~n214 & ~n522;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~n529 & n532;
  assign n534 = ~n528 & n533;
  assign n535 = ~n526 & n534;
  assign O13 = n524 | ~n535;
  assign n537 = inA14 & n101;
  assign n538 = inC14 & n103;
  assign n539 = ~n537 & ~n538;
  assign n540 = n153 & ~n539;
  assign n541 = n152 & n539;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~n473 & ~n542;
  assign n544 = n473 & n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~inA14 & ~musel2;
  assign n547 = ~n225 & n546;
  assign n548 = ~n224 & n547;
  assign n549 = ~inC14 & musel2;
  assign n550 = ~n225 & n549;
  assign n551 = ~n224 & n550;
  assign n552 = ~inA14 & ~inB14;
  assign n553 = ~musel2 & n552;
  assign n554 = ~n224 & n553;
  assign n555 = ~inB14 & ~inC14;
  assign n556 = musel2 & n555;
  assign n557 = ~n224 & n556;
  assign n558 = ~inA14 & ~inD14;
  assign n559 = ~musel2 & n558;
  assign n560 = ~n225 & n559;
  assign n561 = ~inC14 & ~inD14;
  assign n562 = musel2 & n561;
  assign n563 = ~n225 & n562;
  assign n564 = ~inD14 & n552;
  assign n565 = ~musel2 & n564;
  assign n566 = ~inD14 & n555;
  assign n567 = musel2 & n566;
  assign n568 = ~inB14 & ~n226;
  assign n569 = ~n224 & n568;
  assign n570 = ~inD14 & ~n226;
  assign n571 = ~n225 & n570;
  assign n572 = ~inB14 & ~inD14;
  assign n573 = ~n226 & n572;
  assign n574 = ~musel4 & ~n573;
  assign n575 = ~n571 & n574;
  assign n576 = ~n569 & n575;
  assign n577 = ~n250 & n576;
  assign n578 = ~n567 & n577;
  assign n579 = ~n565 & n578;
  assign n580 = ~n563 & n579;
  assign n581 = ~n560 & n580;
  assign n582 = ~n557 & n581;
  assign n583 = ~n554 & n582;
  assign n584 = ~n551 & n583;
  assign n585 = ~n548 & n584;
  assign n586 = inC14 & n539;
  assign n587 = n107 & n586;
  assign n588 = inA14 & n104;
  assign n589 = n215 & ~n539;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n587 & n590;
  assign n592 = inC14 & n110;
  assign n593 = n591 & ~n592;
  assign n594 = ~n585 & n593;
  assign n595 = ~n115 & n466;
  assign n596 = ~n120 & n272;
  assign n597 = ~n148 & ~n545;
  assign n598 = ~n214 & ~n594;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n596 & n599;
  assign O14 = n595 | ~n600;
  assign n602 = inC15 & n151;
  assign n603 = n107 & n602;
  assign n604 = inA15 & n104;
  assign n605 = ~n151 & n215;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n603 & n606;
  assign n608 = inC15 & n110;
  assign n609 = n607 & ~n608;
  assign n610 = ~inA15 & ~musel2;
  assign n611 = ~n225 & n610;
  assign n612 = ~n224 & n611;
  assign n613 = ~inC15 & musel2;
  assign n614 = ~n225 & n613;
  assign n615 = ~n224 & n614;
  assign n616 = ~inA15 & ~inB15;
  assign n617 = ~musel2 & n616;
  assign n618 = ~n224 & n617;
  assign n619 = ~inB15 & ~inC15;
  assign n620 = musel2 & n619;
  assign n621 = ~n224 & n620;
  assign n622 = ~inA15 & ~inD15;
  assign n623 = ~musel2 & n622;
  assign n624 = ~n225 & n623;
  assign n625 = ~inC15 & ~inD15;
  assign n626 = musel2 & n625;
  assign n627 = ~n225 & n626;
  assign n628 = ~inD15 & n616;
  assign n629 = ~musel2 & n628;
  assign n630 = ~inD15 & n619;
  assign n631 = musel2 & n630;
  assign n632 = ~inB15 & ~n226;
  assign n633 = ~n224 & n632;
  assign n634 = ~inD15 & ~n226;
  assign n635 = ~n225 & n634;
  assign n636 = ~inB15 & ~inD15;
  assign n637 = ~n226 & n636;
  assign n638 = ~musel4 & ~n637;
  assign n639 = ~n635 & n638;
  assign n640 = ~n633 & n639;
  assign n641 = ~n250 & n640;
  assign n642 = ~n631 & n641;
  assign n643 = ~n629 & n642;
  assign n644 = ~n627 & n643;
  assign n645 = ~n624 & n644;
  assign n646 = ~n621 & n645;
  assign n647 = ~n618 & n646;
  assign n648 = ~n615 & n647;
  assign n649 = ~n612 & n648;
  assign n650 = n609 & ~n649;
  assign n651 = ~n542 & n545;
  assign n652 = ~n148 & n651;
  assign n653 = ~n214 & ~n650;
  assign n654 = ~n272 & ~n653;
  assign O15 = n652 | ~n654;
  assign n656 = inB4 & ~n106;
  assign n657 = inD4 & ~n112;
  assign n658 = ~n656 & ~n657;
  assign n659 = inB8 & ~n106;
  assign n660 = inD8 & ~n112;
  assign n661 = ~n659 & ~n660;
  assign n662 = inB5 & ~n106;
  assign n663 = inD5 & ~n112;
  assign n664 = ~n662 & ~n663;
  assign n665 = inB3 & ~n106;
  assign n666 = inD3 & ~n112;
  assign n667 = ~n665 & ~n666;
  assign n668 = inB2 & ~n106;
  assign n669 = inD2 & ~n112;
  assign n670 = ~n668 & ~n669;
  assign n671 = inB1 & ~n106;
  assign n672 = inD1 & ~n112;
  assign n673 = ~n671 & ~n672;
  assign n674 = inC0 & n156;
  assign n675 = n107 & n674;
  assign n676 = inA0 & n104;
  assign n677 = ~n156 & n215;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n675 & n678;
  assign n680 = inC0 & n110;
  assign n681 = n679 & ~n680;
  assign n682 = ~inA0 & ~musel2;
  assign n683 = ~n225 & n682;
  assign n684 = ~n224 & n683;
  assign n685 = ~inC0 & musel2;
  assign n686 = ~n225 & n685;
  assign n687 = ~n224 & n686;
  assign n688 = ~inA0 & ~inB0;
  assign n689 = ~musel2 & n688;
  assign n690 = ~n224 & n689;
  assign n691 = ~inB0 & ~inC0;
  assign n692 = musel2 & n691;
  assign n693 = ~n224 & n692;
  assign n694 = ~inA0 & ~inD0;
  assign n695 = ~musel2 & n694;
  assign n696 = ~n225 & n695;
  assign n697 = ~inC0 & ~inD0;
  assign n698 = musel2 & n697;
  assign n699 = ~n225 & n698;
  assign n700 = ~inD0 & n688;
  assign n701 = ~musel2 & n700;
  assign n702 = ~inD0 & n691;
  assign n703 = musel2 & n702;
  assign n704 = ~inB0 & ~n226;
  assign n705 = ~n224 & n704;
  assign n706 = ~inD0 & ~n226;
  assign n707 = ~n225 & n706;
  assign n708 = ~inB0 & ~inD0;
  assign n709 = ~n226 & n708;
  assign n710 = ~musel4 & ~n709;
  assign n711 = ~n707 & n710;
  assign n712 = ~n705 & n711;
  assign n713 = ~n250 & n712;
  assign n714 = ~n703 & n713;
  assign n715 = ~n701 & n714;
  assign n716 = ~n699 & n715;
  assign n717 = ~n696 & n716;
  assign n718 = ~n693 & n717;
  assign n719 = ~n690 & n718;
  assign n720 = ~n687 & n719;
  assign n721 = ~n684 & n720;
  assign n722 = n681 & ~n721;
  assign n723 = inB0 & ~n106;
  assign n724 = n466 & n723;
  assign n725 = inD0 & ~n112;
  assign n726 = n466 & n725;
  assign n727 = ~n148 & ~n159;
  assign n728 = ~n160 & n727;
  assign n729 = ~n148 & n152;
  assign n730 = ~n160 & n729;
  assign n731 = ~n100 & ~n658;
  assign n732 = n93 & n731;
  assign n733 = ~n100 & ~n661;
  assign n734 = n143 & n733;
  assign n735 = ~n100 & ~n664;
  assign n736 = n121 & n735;
  assign n737 = ~n100 & ~n667;
  assign n738 = n126 & n737;
  assign n739 = ~n100 & ~n670;
  assign n740 = n130 & n739;
  assign n741 = n465 & ~n673;
  assign n742 = ~n214 & ~n722;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n740 & n743;
  assign n745 = ~n738 & n744;
  assign n746 = ~n736 & n745;
  assign n747 = ~n734 & n746;
  assign n748 = ~n732 & n747;
  assign n749 = ~n730 & n748;
  assign n750 = ~n728 & n749;
  assign n751 = ~n726 & n750;
  assign O0 = n724 | ~n751;
  assign n753 = inB9 & ~n106;
  assign n754 = inD9 & ~n112;
  assign n755 = ~n753 & ~n754;
  assign n756 = inB6 & ~n106;
  assign n757 = inD6 & ~n112;
  assign n758 = ~n756 & ~n757;
  assign n759 = inC1 & n163;
  assign n760 = n107 & n759;
  assign n761 = inA1 & n104;
  assign n762 = ~n163 & n215;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n760 & n763;
  assign n765 = inC1 & n110;
  assign n766 = n764 & ~n765;
  assign n767 = ~inA1 & ~musel2;
  assign n768 = ~n225 & n767;
  assign n769 = ~n224 & n768;
  assign n770 = ~inC1 & musel2;
  assign n771 = ~n225 & n770;
  assign n772 = ~n224 & n771;
  assign n773 = ~inA1 & ~inB1;
  assign n774 = ~musel2 & n773;
  assign n775 = ~n224 & n774;
  assign n776 = ~inB1 & ~inC1;
  assign n777 = musel2 & n776;
  assign n778 = ~n224 & n777;
  assign n779 = ~inA1 & ~inD1;
  assign n780 = ~musel2 & n779;
  assign n781 = ~n225 & n780;
  assign n782 = ~inC1 & ~inD1;
  assign n783 = musel2 & n782;
  assign n784 = ~n225 & n783;
  assign n785 = ~inD1 & n773;
  assign n786 = ~musel2 & n785;
  assign n787 = ~inD1 & n776;
  assign n788 = musel2 & n787;
  assign n789 = ~inB1 & ~n226;
  assign n790 = ~n224 & n789;
  assign n791 = ~inD1 & ~n226;
  assign n792 = ~n225 & n791;
  assign n793 = ~inB1 & ~inD1;
  assign n794 = ~n226 & n793;
  assign n795 = ~musel4 & ~n794;
  assign n796 = ~n792 & n795;
  assign n797 = ~n790 & n796;
  assign n798 = ~n250 & n797;
  assign n799 = ~n788 & n798;
  assign n800 = ~n786 & n799;
  assign n801 = ~n784 & n800;
  assign n802 = ~n781 & n801;
  assign n803 = ~n778 & n802;
  assign n804 = ~n775 & n803;
  assign n805 = ~n772 & n804;
  assign n806 = ~n769 & n805;
  assign n807 = n766 & ~n806;
  assign n808 = ~n148 & n166;
  assign n809 = n160 & n808;
  assign n810 = ~n148 & ~n166;
  assign n811 = ~n160 & n810;
  assign n812 = n93 & n735;
  assign n813 = ~n100 & ~n755;
  assign n814 = n143 & n813;
  assign n815 = ~n100 & ~n758;
  assign n816 = n121 & n815;
  assign n817 = n126 & n731;
  assign n818 = n130 & n737;
  assign n819 = n465 & ~n670;
  assign n820 = n466 & ~n673;
  assign n821 = ~n214 & ~n807;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~n819 & n822;
  assign n824 = ~n818 & n823;
  assign n825 = ~n817 & n824;
  assign n826 = ~n816 & n825;
  assign n827 = ~n814 & n826;
  assign n828 = ~n812 & n827;
  assign n829 = ~n811 & n828;
  assign O1 = n809 | ~n829;
  assign n831 = inB7 & ~n106;
  assign n832 = inD7 & ~n112;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n167 & ~n173;
  assign n835 = n167 & n173;
  assign n836 = ~n834 & ~n835;
  assign n837 = inC2 & n170;
  assign n838 = n107 & n837;
  assign n839 = inA2 & n104;
  assign n840 = ~n170 & n215;
  assign n841 = ~n839 & ~n840;
  assign n842 = ~n838 & n841;
  assign n843 = inC2 & n110;
  assign n844 = n842 & ~n843;
  assign n845 = ~inA2 & ~musel2;
  assign n846 = ~n225 & n845;
  assign n847 = ~n224 & n846;
  assign n848 = ~inC2 & musel2;
  assign n849 = ~n225 & n848;
  assign n850 = ~n224 & n849;
  assign n851 = ~inA2 & ~inB2;
  assign n852 = ~musel2 & n851;
  assign n853 = ~n224 & n852;
  assign n854 = ~inB2 & ~inC2;
  assign n855 = musel2 & n854;
  assign n856 = ~n224 & n855;
  assign n857 = ~inA2 & ~inD2;
  assign n858 = ~musel2 & n857;
  assign n859 = ~n225 & n858;
  assign n860 = ~inC2 & ~inD2;
  assign n861 = musel2 & n860;
  assign n862 = ~n225 & n861;
  assign n863 = ~inD2 & n851;
  assign n864 = ~musel2 & n863;
  assign n865 = ~inD2 & n854;
  assign n866 = musel2 & n865;
  assign n867 = ~inB2 & ~n226;
  assign n868 = ~n224 & n867;
  assign n869 = ~inD2 & ~n226;
  assign n870 = ~n225 & n869;
  assign n871 = ~inB2 & ~inD2;
  assign n872 = ~n226 & n871;
  assign n873 = ~musel4 & ~n872;
  assign n874 = ~n870 & n873;
  assign n875 = ~n868 & n874;
  assign n876 = ~n250 & n875;
  assign n877 = ~n866 & n876;
  assign n878 = ~n864 & n877;
  assign n879 = ~n862 & n878;
  assign n880 = ~n859 & n879;
  assign n881 = ~n856 & n880;
  assign n882 = ~n853 & n881;
  assign n883 = ~n850 & n882;
  assign n884 = ~n847 & n883;
  assign n885 = n844 & ~n884;
  assign n886 = n93 & n815;
  assign n887 = ~n100 & ~n141;
  assign n888 = n143 & n887;
  assign n889 = ~n100 & ~n833;
  assign n890 = n121 & n889;
  assign n891 = n126 & n735;
  assign n892 = n130 & n731;
  assign n893 = n465 & ~n667;
  assign n894 = n466 & ~n670;
  assign n895 = ~n214 & ~n885;
  assign n896 = ~n148 & ~n836;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n894 & n897;
  assign n899 = ~n893 & n898;
  assign n900 = ~n892 & n899;
  assign n901 = ~n891 & n900;
  assign n902 = ~n890 & n901;
  assign n903 = ~n888 & n902;
  assign O2 = n886 | ~n903;
  assign n905 = inC3 & n176;
  assign n906 = n107 & n905;
  assign n907 = inA3 & n104;
  assign n908 = ~n176 & n215;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n906 & n909;
  assign n911 = inC3 & n110;
  assign n912 = n910 & ~n911;
  assign n913 = ~inA3 & ~musel2;
  assign n914 = ~n225 & n913;
  assign n915 = ~n224 & n914;
  assign n916 = ~inC3 & musel2;
  assign n917 = ~n225 & n916;
  assign n918 = ~n224 & n917;
  assign n919 = ~inA3 & ~inB3;
  assign n920 = ~musel2 & n919;
  assign n921 = ~n224 & n920;
  assign n922 = ~inB3 & ~inC3;
  assign n923 = musel2 & n922;
  assign n924 = ~n224 & n923;
  assign n925 = ~inA3 & ~inD3;
  assign n926 = ~musel2 & n925;
  assign n927 = ~n225 & n926;
  assign n928 = ~inC3 & ~inD3;
  assign n929 = musel2 & n928;
  assign n930 = ~n225 & n929;
  assign n931 = ~inD3 & n919;
  assign n932 = ~musel2 & n931;
  assign n933 = ~inD3 & n922;
  assign n934 = musel2 & n933;
  assign n935 = ~inB3 & ~n226;
  assign n936 = ~n224 & n935;
  assign n937 = ~inD3 & ~n226;
  assign n938 = ~n225 & n937;
  assign n939 = ~inB3 & ~inD3;
  assign n940 = ~n226 & n939;
  assign n941 = ~musel4 & ~n940;
  assign n942 = ~n938 & n941;
  assign n943 = ~n936 & n942;
  assign n944 = ~n250 & n943;
  assign n945 = ~n934 & n944;
  assign n946 = ~n932 & n945;
  assign n947 = ~n930 & n946;
  assign n948 = ~n927 & n947;
  assign n949 = ~n924 & n948;
  assign n950 = ~n921 & n949;
  assign n951 = ~n918 & n950;
  assign n952 = ~n915 & n951;
  assign n953 = n912 & ~n952;
  assign n954 = ~n173 & ~n181;
  assign n955 = n836 & n954;
  assign n956 = ~n148 & n955;
  assign n957 = n93 & n889;
  assign n958 = n143 & n278;
  assign n959 = n121 & n733;
  assign n960 = n126 & n815;
  assign n961 = n130 & n735;
  assign n962 = n135 & n731;
  assign n963 = ~n179 & ~n181;
  assign n964 = ~n148 & n963;
  assign n965 = n120 & ~n667;
  assign n966 = ~n100 & n965;
  assign n967 = ~n214 & ~n953;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~n964 & n968;
  assign n970 = ~n962 & n969;
  assign n971 = ~n961 & n970;
  assign n972 = ~n960 & n971;
  assign n973 = ~n959 & n972;
  assign n974 = ~n958 & n973;
  assign n975 = ~n957 & n974;
  assign O3 = n956 | ~n975;
  assign n977 = inC4 & n364;
  assign n978 = n107 & n977;
  assign n979 = inA4 & n104;
  assign n980 = n215 & ~n364;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n978 & n981;
  assign n983 = inC4 & n110;
  assign n984 = n982 & ~n983;
  assign n985 = ~inA4 & ~musel2;
  assign n986 = ~n225 & n985;
  assign n987 = ~n224 & n986;
  assign n988 = ~inC4 & musel2;
  assign n989 = ~n225 & n988;
  assign n990 = ~n224 & n989;
  assign n991 = ~inA4 & ~inB4;
  assign n992 = ~musel2 & n991;
  assign n993 = ~n224 & n992;
  assign n994 = ~inB4 & ~inC4;
  assign n995 = musel2 & n994;
  assign n996 = ~n224 & n995;
  assign n997 = ~inA4 & ~inD4;
  assign n998 = ~musel2 & n997;
  assign n999 = ~n225 & n998;
  assign n1000 = ~inC4 & ~inD4;
  assign n1001 = musel2 & n1000;
  assign n1002 = ~n225 & n1001;
  assign n1003 = ~inD4 & n991;
  assign n1004 = ~musel2 & n1003;
  assign n1005 = ~inD4 & n994;
  assign n1006 = musel2 & n1005;
  assign n1007 = ~inB4 & ~n226;
  assign n1008 = ~n224 & n1007;
  assign n1009 = ~inD4 & ~n226;
  assign n1010 = ~n225 & n1009;
  assign n1011 = ~inB4 & ~inD4;
  assign n1012 = ~n226 & n1011;
  assign n1013 = ~musel4 & ~n1012;
  assign n1014 = ~n1010 & n1013;
  assign n1015 = ~n1008 & n1014;
  assign n1016 = ~n250 & n1015;
  assign n1017 = ~n1006 & n1016;
  assign n1018 = ~n1004 & n1017;
  assign n1019 = ~n1002 & n1018;
  assign n1020 = ~n999 & n1019;
  assign n1021 = ~n996 & n1020;
  assign n1022 = ~n993 & n1021;
  assign n1023 = ~n990 & n1022;
  assign n1024 = ~n987 & n1023;
  assign n1025 = n984 & ~n1024;
  assign n1026 = ~n358 & ~n661;
  assign n1027 = n93 & n1026;
  assign n1028 = ~n133 & ~n358;
  assign n1029 = n143 & n1028;
  assign n1030 = ~n358 & ~n755;
  assign n1031 = n121 & n1030;
  assign n1032 = ~n358 & ~n833;
  assign n1033 = n126 & n1032;
  assign n1034 = ~n181 & ~n367;
  assign n1035 = ~n148 & n1034;
  assign n1036 = n181 & n367;
  assign n1037 = ~n148 & n1036;
  assign n1038 = n359 & ~n664;
  assign n1039 = n360 & ~n658;
  assign n1040 = n361 & ~n758;
  assign n1041 = ~n214 & ~n1025;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n1039 & n1042;
  assign n1044 = ~n1038 & n1043;
  assign n1045 = ~n1037 & n1044;
  assign n1046 = ~n1035 & n1045;
  assign n1047 = ~n1033 & n1046;
  assign n1048 = ~n1031 & n1047;
  assign n1049 = ~n1029 & n1048;
  assign O4 = n1027 | ~n1049;
  assign n1051 = n181 & ~n367;
  assign n1052 = inC5 & n370;
  assign n1053 = n107 & n1052;
  assign n1054 = inA5 & n104;
  assign n1055 = n215 & ~n370;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1053 & n1056;
  assign n1058 = inC5 & n110;
  assign n1059 = n1057 & ~n1058;
  assign n1060 = ~inA5 & ~musel2;
  assign n1061 = ~n225 & n1060;
  assign n1062 = ~n224 & n1061;
  assign n1063 = ~inC5 & musel2;
  assign n1064 = ~n225 & n1063;
  assign n1065 = ~n224 & n1064;
  assign n1066 = ~inA5 & ~inB5;
  assign n1067 = ~musel2 & n1066;
  assign n1068 = ~n224 & n1067;
  assign n1069 = ~inB5 & ~inC5;
  assign n1070 = musel2 & n1069;
  assign n1071 = ~n224 & n1070;
  assign n1072 = ~inA5 & ~inD5;
  assign n1073 = ~musel2 & n1072;
  assign n1074 = ~n225 & n1073;
  assign n1075 = ~inC5 & ~inD5;
  assign n1076 = musel2 & n1075;
  assign n1077 = ~n225 & n1076;
  assign n1078 = ~inD5 & n1066;
  assign n1079 = ~musel2 & n1078;
  assign n1080 = ~inD5 & n1069;
  assign n1081 = musel2 & n1080;
  assign n1082 = ~inB5 & ~n226;
  assign n1083 = ~n224 & n1082;
  assign n1084 = ~inD5 & ~n226;
  assign n1085 = ~n225 & n1084;
  assign n1086 = ~inB5 & ~inD5;
  assign n1087 = ~n226 & n1086;
  assign n1088 = ~musel4 & ~n1087;
  assign n1089 = ~n1085 & n1088;
  assign n1090 = ~n1083 & n1089;
  assign n1091 = ~n250 & n1090;
  assign n1092 = ~n1081 & n1091;
  assign n1093 = ~n1079 & n1092;
  assign n1094 = ~n1077 & n1093;
  assign n1095 = ~n1074 & n1094;
  assign n1096 = ~n1071 & n1095;
  assign n1097 = ~n1068 & n1096;
  assign n1098 = ~n1065 & n1097;
  assign n1099 = ~n1062 & n1098;
  assign n1100 = n1059 & ~n1099;
  assign n1101 = ~n148 & n373;
  assign n1102 = n1051 & n1101;
  assign n1103 = ~n148 & ~n373;
  assign n1104 = ~n1051 & n1103;
  assign n1105 = n93 & n813;
  assign n1106 = n143 & n274;
  assign n1107 = n121 & n887;
  assign n1108 = n126 & n733;
  assign n1109 = n130 & n889;
  assign n1110 = n465 & ~n758;
  assign n1111 = n466 & ~n664;
  assign n1112 = ~n214 & ~n1100;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1110 & n1113;
  assign n1115 = ~n1109 & n1114;
  assign n1116 = ~n1108 & n1115;
  assign n1117 = ~n1107 & n1116;
  assign n1118 = ~n1106 & n1117;
  assign n1119 = ~n1105 & n1118;
  assign n1120 = ~n1104 & n1119;
  assign O5 = n1102 | ~n1120;
  assign n1122 = ~n373 & n1051;
  assign n1123 = ~n379 & ~n1122;
  assign n1124 = n379 & n1122;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = inC6 & n376;
  assign n1127 = n107 & n1126;
  assign n1128 = inA6 & n104;
  assign n1129 = n215 & ~n376;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1127 & n1130;
  assign n1132 = inC6 & n110;
  assign n1133 = n1131 & ~n1132;
  assign n1134 = ~inA6 & ~musel2;
  assign n1135 = ~n225 & n1134;
  assign n1136 = ~n224 & n1135;
  assign n1137 = ~inC6 & musel2;
  assign n1138 = ~n225 & n1137;
  assign n1139 = ~n224 & n1138;
  assign n1140 = ~inA6 & ~inB6;
  assign n1141 = ~musel2 & n1140;
  assign n1142 = ~n224 & n1141;
  assign n1143 = ~inB6 & ~inC6;
  assign n1144 = musel2 & n1143;
  assign n1145 = ~n224 & n1144;
  assign n1146 = ~inA6 & ~inD6;
  assign n1147 = ~musel2 & n1146;
  assign n1148 = ~n225 & n1147;
  assign n1149 = ~inC6 & ~inD6;
  assign n1150 = musel2 & n1149;
  assign n1151 = ~n225 & n1150;
  assign n1152 = ~inD6 & n1140;
  assign n1153 = ~musel2 & n1152;
  assign n1154 = ~inD6 & n1143;
  assign n1155 = musel2 & n1154;
  assign n1156 = ~inB6 & ~n226;
  assign n1157 = ~n224 & n1156;
  assign n1158 = ~inD6 & ~n226;
  assign n1159 = ~n225 & n1158;
  assign n1160 = ~inB6 & ~inD6;
  assign n1161 = ~n226 & n1160;
  assign n1162 = ~musel4 & ~n1161;
  assign n1163 = ~n1159 & n1162;
  assign n1164 = ~n1157 & n1163;
  assign n1165 = ~n250 & n1164;
  assign n1166 = ~n1155 & n1165;
  assign n1167 = ~n1153 & n1166;
  assign n1168 = ~n1151 & n1167;
  assign n1169 = ~n1148 & n1168;
  assign n1170 = ~n1145 & n1169;
  assign n1171 = ~n1142 & n1170;
  assign n1172 = ~n1139 & n1171;
  assign n1173 = ~n1136 & n1172;
  assign n1174 = n1133 & ~n1173;
  assign n1175 = n93 & n887;
  assign n1176 = n143 & n270;
  assign n1177 = n121 & n278;
  assign n1178 = n126 & n813;
  assign n1179 = n130 & n733;
  assign n1180 = n465 & ~n833;
  assign n1181 = n466 & ~n758;
  assign n1182 = ~n214 & ~n1174;
  assign n1183 = ~n148 & ~n1125;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1181 & n1184;
  assign n1186 = ~n1180 & n1185;
  assign n1187 = ~n1179 & n1186;
  assign n1188 = ~n1178 & n1187;
  assign n1189 = ~n1177 & n1188;
  assign n1190 = ~n1176 & n1189;
  assign O6 = n1175 | ~n1190;
  assign n1192 = ~n379 & n1125;
  assign n1193 = inC7 & n382;
  assign n1194 = n107 & n1193;
  assign n1195 = inA7 & n104;
  assign n1196 = n215 & ~n382;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1194 & n1197;
  assign n1199 = inC7 & n110;
  assign n1200 = n1198 & ~n1199;
  assign n1201 = ~inA7 & ~musel2;
  assign n1202 = ~n225 & n1201;
  assign n1203 = ~n224 & n1202;
  assign n1204 = ~inC7 & musel2;
  assign n1205 = ~n225 & n1204;
  assign n1206 = ~n224 & n1205;
  assign n1207 = ~inA7 & ~inB7;
  assign n1208 = ~musel2 & n1207;
  assign n1209 = ~n224 & n1208;
  assign n1210 = ~inB7 & ~inC7;
  assign n1211 = musel2 & n1210;
  assign n1212 = ~n224 & n1211;
  assign n1213 = ~inA7 & ~inD7;
  assign n1214 = ~musel2 & n1213;
  assign n1215 = ~n225 & n1214;
  assign n1216 = ~inC7 & ~inD7;
  assign n1217 = musel2 & n1216;
  assign n1218 = ~n225 & n1217;
  assign n1219 = ~inD7 & n1207;
  assign n1220 = ~musel2 & n1219;
  assign n1221 = ~inD7 & n1210;
  assign n1222 = musel2 & n1221;
  assign n1223 = ~inB7 & ~n226;
  assign n1224 = ~n224 & n1223;
  assign n1225 = ~inD7 & ~n226;
  assign n1226 = ~n225 & n1225;
  assign n1227 = ~inB7 & ~inD7;
  assign n1228 = ~n226 & n1227;
  assign n1229 = ~musel4 & ~n1228;
  assign n1230 = ~n1226 & n1229;
  assign n1231 = ~n1224 & n1230;
  assign n1232 = ~n250 & n1231;
  assign n1233 = ~n1222 & n1232;
  assign n1234 = ~n1220 & n1233;
  assign n1235 = ~n1218 & n1234;
  assign n1236 = ~n1215 & n1235;
  assign n1237 = ~n1212 & n1236;
  assign n1238 = ~n1209 & n1237;
  assign n1239 = ~n1206 & n1238;
  assign n1240 = ~n1203 & n1239;
  assign n1241 = n1200 & ~n1240;
  assign n1242 = ~n148 & n385;
  assign n1243 = n1192 & n1242;
  assign n1244 = ~n148 & ~n385;
  assign n1245 = ~n1192 & n1244;
  assign n1246 = n93 & n278;
  assign n1247 = n121 & n276;
  assign n1248 = n126 & n887;
  assign n1249 = n130 & n813;
  assign n1250 = n135 & n733;
  assign n1251 = n120 & ~n833;
  assign n1252 = ~n100 & n1251;
  assign n1253 = ~n214 & ~n1241;
  assign n1254 = ~n282 & ~n1253;
  assign n1255 = ~n1252 & n1254;
  assign n1256 = ~n1250 & n1255;
  assign n1257 = ~n1249 & n1256;
  assign n1258 = ~n1248 & n1257;
  assign n1259 = ~n1247 & n1258;
  assign n1260 = ~n1246 & n1259;
  assign n1261 = ~n1245 & n1260;
  assign O7 = n1243 | ~n1261;
  assign n1263 = inC8 & n184;
  assign n1264 = n107 & n1263;
  assign n1265 = inA8 & n104;
  assign n1266 = ~n184 & n215;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = ~n1264 & n1267;
  assign n1269 = inC8 & n110;
  assign n1270 = n1268 & ~n1269;
  assign n1271 = ~inA8 & ~musel2;
  assign n1272 = ~n225 & n1271;
  assign n1273 = ~n224 & n1272;
  assign n1274 = ~inC8 & musel2;
  assign n1275 = ~n225 & n1274;
  assign n1276 = ~n224 & n1275;
  assign n1277 = ~inA8 & ~inB8;
  assign n1278 = ~musel2 & n1277;
  assign n1279 = ~n224 & n1278;
  assign n1280 = ~inB8 & ~inC8;
  assign n1281 = musel2 & n1280;
  assign n1282 = ~n224 & n1281;
  assign n1283 = ~inA8 & ~inD8;
  assign n1284 = ~musel2 & n1283;
  assign n1285 = ~n225 & n1284;
  assign n1286 = ~inC8 & ~inD8;
  assign n1287 = musel2 & n1286;
  assign n1288 = ~n225 & n1287;
  assign n1289 = ~inD8 & n1277;
  assign n1290 = ~musel2 & n1289;
  assign n1291 = ~inD8 & n1280;
  assign n1292 = musel2 & n1291;
  assign n1293 = ~inB8 & ~n226;
  assign n1294 = ~n224 & n1293;
  assign n1295 = ~inD8 & ~n226;
  assign n1296 = ~n225 & n1295;
  assign n1297 = ~inB8 & ~inD8;
  assign n1298 = ~n226 & n1297;
  assign n1299 = ~musel4 & ~n1298;
  assign n1300 = ~n1296 & n1299;
  assign n1301 = ~n1294 & n1300;
  assign n1302 = ~n250 & n1301;
  assign n1303 = ~n1292 & n1302;
  assign n1304 = ~n1290 & n1303;
  assign n1305 = ~n1288 & n1304;
  assign n1306 = ~n1285 & n1305;
  assign n1307 = ~n1282 & n1306;
  assign n1308 = ~n1279 & n1307;
  assign n1309 = ~n1276 & n1308;
  assign n1310 = ~n1273 & n1309;
  assign n1311 = n1270 & ~n1310;
  assign n1312 = n93 & n1028;
  assign n1313 = ~n129 & ~n358;
  assign n1314 = n121 & n1313;
  assign n1315 = ~n138 & ~n358;
  assign n1316 = n126 & n1315;
  assign n1317 = ~n187 & ~n209;
  assign n1318 = ~n148 & n1317;
  assign n1319 = n359 & ~n755;
  assign n1320 = n360 & ~n661;
  assign n1321 = ~n141 & n361;
  assign n1322 = n144 & ~n358;
  assign n1323 = ~n214 & ~n1311;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1321 & n1324;
  assign n1326 = ~n1320 & n1325;
  assign n1327 = ~n1319 & n1326;
  assign n1328 = ~n1318 & n1327;
  assign n1329 = ~n1316 & n1328;
  assign n1330 = ~n1314 & n1329;
  assign O8 = n1312 | ~n1330;
  assign n1332 = inC9 & n190;
  assign n1333 = n107 & n1332;
  assign n1334 = inA9 & n104;
  assign n1335 = ~n190 & n215;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~n1333 & n1336;
  assign n1338 = inC9 & n110;
  assign n1339 = n1337 & ~n1338;
  assign n1340 = ~inA9 & ~musel2;
  assign n1341 = ~n225 & n1340;
  assign n1342 = ~n224 & n1341;
  assign n1343 = ~inC9 & musel2;
  assign n1344 = ~n225 & n1343;
  assign n1345 = ~n224 & n1344;
  assign n1346 = ~inA9 & ~inB9;
  assign n1347 = ~musel2 & n1346;
  assign n1348 = ~n224 & n1347;
  assign n1349 = ~inB9 & ~inC9;
  assign n1350 = musel2 & n1349;
  assign n1351 = ~n224 & n1350;
  assign n1352 = ~inA9 & ~inD9;
  assign n1353 = ~musel2 & n1352;
  assign n1354 = ~n225 & n1353;
  assign n1355 = ~inC9 & ~inD9;
  assign n1356 = musel2 & n1355;
  assign n1357 = ~n225 & n1356;
  assign n1358 = ~inD9 & n1346;
  assign n1359 = ~musel2 & n1358;
  assign n1360 = ~inD9 & n1349;
  assign n1361 = musel2 & n1360;
  assign n1362 = ~inB9 & ~n226;
  assign n1363 = ~n224 & n1362;
  assign n1364 = ~inD9 & ~n226;
  assign n1365 = ~n225 & n1364;
  assign n1366 = ~inB9 & ~inD9;
  assign n1367 = ~n226 & n1366;
  assign n1368 = ~musel4 & ~n1367;
  assign n1369 = ~n1365 & n1368;
  assign n1370 = ~n1363 & n1369;
  assign n1371 = ~n250 & n1370;
  assign n1372 = ~n1361 & n1371;
  assign n1373 = ~n1359 & n1372;
  assign n1374 = ~n1357 & n1373;
  assign n1375 = ~n1354 & n1374;
  assign n1376 = ~n1351 & n1375;
  assign n1377 = ~n1348 & n1376;
  assign n1378 = ~n1345 & n1377;
  assign n1379 = ~n1342 & n1378;
  assign n1380 = n1339 & ~n1379;
  assign n1381 = ~n148 & ~n193;
  assign n1382 = ~n209 & n1381;
  assign n1383 = n93 & n274;
  assign n1384 = n121 & n270;
  assign n1385 = n126 & n276;
  assign n1386 = n130 & n278;
  assign n1387 = ~n141 & n465;
  assign n1388 = n466 & ~n755;
  assign n1389 = ~n214 & ~n1380;
  assign n1390 = ~n282 & ~n1389;
  assign n1391 = ~n1388 & n1390;
  assign n1392 = ~n1387 & n1391;
  assign n1393 = ~n1386 & n1392;
  assign n1394 = ~n1385 & n1393;
  assign n1395 = ~n1384 & n1394;
  assign n1396 = ~n1383 & n1395;
  assign O9 = n1382 | ~n1396;
endmodule


