// Benchmark "i9" written by ABC on Tue May 16 16:07:51 2017

module i9 ( 
    \V88(21) , \V88(20) , \V88(27) , \V9(0) , \V88(0) , \V88(26) , \V9(1) ,
    \V88(1) , \V88(29) , \V9(2) , \V88(2) , \V88(28) , \V9(3) , \V88(3) ,
    \V88(4) , \V9(5) , \V88(5) , \V9(6) , \V88(6) , \V56(13) , \V9(7) ,
    \V88(7) , \V56(12) , \V9(8) , \V9(10) , \V88(8) , \V56(15) , \V88(9) ,
    \V88(31) , \V56(14) , \V88(30) , \V56(11) , \V56(10) , \V56(17) ,
    \V56(0) , \V56(16) , \V56(1) , \V56(19) , \V56(2) , \V56(18) ,
    \V56(3) , \V56(23) , \V56(4) , \V56(22) , \V56(5) , \V56(25) ,
    \V56(6) , \V56(24) , \V56(7) , \V56(8) , \V56(9) , \V56(21) ,
    \V56(20) , \V56(27) , \V56(26) , \V56(29) , \V56(28) , \V24(0) ,
    \V88(13) , \V24(1) , \V88(12) , \V24(2) , \V88(15) , \V24(3) ,
    \V24(13) , \V88(14) , \V24(4) , \V24(12) , \V24(5) , \V56(31) ,
    \V24(6) , \V24(14) , \V88(11) , \V56(30) , \V24(7) , \V88(10) ,
    \V24(8) , \V24(9) , \V24(11) , \V24(10) , \V88(17) , \V88(16) ,
    \V88(19) , \V88(18) , \V88(23) , \V88(22) , \V88(25) , \V88(24) ,
    \V119(21) , \V151(16) , \V119(20) , \V151(19) , \V119(23) , \V151(18) ,
    \V119(22) , \V119(25) , \V119(24) , \V119(17) , \V119(16) , \V119(3) ,
    \V119(19) , \V119(2) , \V119(18) , \V151(11) , \V119(5) , \V151(10) ,
    \V119(4) , \V151(13) , \V151(12) , \V151(15) , \V119(1) , \V151(14) ,
    \V119(0) , \V119(11) , \V119(10) , \V119(13) , \V119(12) , \V119(7) ,
    \V119(15) , \V119(6) , \V119(14) , \V119(9) , \V119(8) , \V151(3) ,
    \V151(2) , \V151(5) , \V151(4) , \V151(1) , \V151(0) , \V151(7) ,
    \V151(6) , \V151(9) , \V151(8) , \V151(31) , \V151(30) , \V119(30) ,
    \V151(27) , \V151(26) , \V151(29) , \V151(28) , \V119(27) , \V119(26) ,
    \V119(29) , \V119(28) , \V151(21) , \V151(20) , \V151(23) , \V151(22) ,
    \V151(25) , \V151(24) , \V151(17)   );
  input  \V88(21) , \V88(20) , \V88(27) , \V9(0) , \V88(0) , \V88(26) ,
    \V9(1) , \V88(1) , \V88(29) , \V9(2) , \V88(2) , \V88(28) , \V9(3) ,
    \V88(3) , \V88(4) , \V9(5) , \V88(5) , \V9(6) , \V88(6) , \V56(13) ,
    \V9(7) , \V88(7) , \V56(12) , \V9(8) , \V9(10) , \V88(8) , \V56(15) ,
    \V88(9) , \V88(31) , \V56(14) , \V88(30) , \V56(11) , \V56(10) ,
    \V56(17) , \V56(0) , \V56(16) , \V56(1) , \V56(19) , \V56(2) ,
    \V56(18) , \V56(3) , \V56(23) , \V56(4) , \V56(22) , \V56(5) ,
    \V56(25) , \V56(6) , \V56(24) , \V56(7) , \V56(8) , \V56(9) ,
    \V56(21) , \V56(20) , \V56(27) , \V56(26) , \V56(29) , \V56(28) ,
    \V24(0) , \V88(13) , \V24(1) , \V88(12) , \V24(2) , \V88(15) ,
    \V24(3) , \V24(13) , \V88(14) , \V24(4) , \V24(12) , \V24(5) ,
    \V56(31) , \V24(6) , \V24(14) , \V88(11) , \V56(30) , \V24(7) ,
    \V88(10) , \V24(8) , \V24(9) , \V24(11) , \V24(10) , \V88(17) ,
    \V88(16) , \V88(19) , \V88(18) , \V88(23) , \V88(22) , \V88(25) ,
    \V88(24) ;
  output \V119(21) , \V151(16) , \V119(20) , \V151(19) , \V119(23) ,
    \V151(18) , \V119(22) , \V119(25) , \V119(24) , \V119(17) , \V119(16) ,
    \V119(3) , \V119(19) , \V119(2) , \V119(18) , \V151(11) , \V119(5) ,
    \V151(10) , \V119(4) , \V151(13) , \V151(12) , \V151(15) , \V119(1) ,
    \V151(14) , \V119(0) , \V119(11) , \V119(10) , \V119(13) , \V119(12) ,
    \V119(7) , \V119(15) , \V119(6) , \V119(14) , \V119(9) , \V119(8) ,
    \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) , \V151(0) ,
    \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V151(31) , \V151(30) ,
    \V119(30) , \V151(27) , \V151(26) , \V151(29) , \V151(28) , \V119(27) ,
    \V119(26) , \V119(29) , \V119(28) , \V151(21) , \V151(20) , \V151(23) ,
    \V151(22) , \V151(25) , \V151(24) , \V151(17) ;
  wire n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n208, n209, n210, n211, n212,
    n213, n214, n216, n217, n218, n219, n220, n221, n222, n224, n225, n226,
    n227, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238, n240,
    n241, n242, n243, n244, n245, n246, n248, n249, n250, n251, n252, n253,
    n254, n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267,
    n268, n269, n270, n272, n273, n274, n275, n276, n277, n278, n280, n281,
    n282, n283, n284, n285, n287, n288, n289, n290, n291, n292, n293, n295,
    n296, n297, n298, n299, n301, n302, n303, n304, n305, n306, n307, n309,
    n310, n311, n312, n313, n314, n315, n317, n318, n319, n320, n321, n323,
    n324, n325, n326, n327, n328, n329, n331, n332, n333, n334, n336, n337,
    n338, n339, n340, n341, n342, n344, n345, n346, n347, n348, n349, n350,
    n352, n353, n354, n355, n356, n357, n359, n360, n361, n362, n364, n365,
    n366, n367, n368, n369, n371, n372, n373, n374, n376, n377, n378, n379,
    n380, n381, n382, n384, n385, n386, n387, n388, n389, n390, n392, n393,
    n394, n395, n396, n397, n398, n400, n401, n402, n403, n404, n405, n406,
    n408, n409, n410, n411, n412, n414, n415, n416, n417, n418, n419, n420,
    n422, n423, n424, n425, n427, n428, n429, n430, n431, n432, n433, n435,
    n436, n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n448,
    n449, n451, n452, n453, n454, n455, n456, n457, n459, n460, n461, n462,
    n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n475, n476,
    n477, n478, n479, n480, n481, n483, n484, n485, n486, n487, n488, n489,
    n491, n492, n493, n494, n495, n496, n497, n499, n500, n501, n502, n503,
    n504, n505, n507, n508, n509, n510, n511, n512, n513, n515, n516, n517,
    n518, n519, n520, n521, n523, n524, n525, n526, n527, n528, n529, n531,
    n532, n533, n534, n535, n536, n537, n539, n540, n541, n542, n543, n544,
    n545, n547, n548, n549, n550, n551, n552, n553, n555, n556, n557, n558,
    n559, n560, n561, n563, n564, n565, n566, n567, n568, n569, n571, n572,
    n573, n574, n575, n576, n577, n579, n580, n581, n582, n583, n584, n585,
    n587, n588, n589, n590, n591, n592, n593, n595, n596, n597, n598, n599,
    n600, n601, n603, n604, n605, n606, n607, n608, n609, n611, n612, n613,
    n614, n615, n616, n617, n619, n620, n621, n622, n623, n625, n626, n627,
    n628, n629, n631, n632, n633, n634, n635, n636, n637, n639, n640, n641,
    n642, n643, n645, n646, n647, n648, n649, n650, n651, n653, n654, n655,
    n656, n657, n658, n659, n661, n662, n663, n664, n665, n666;
  assign n152 = ~\V9(7)  & ~\V9(10) ;
  assign n153 = ~\V9(2)  & ~\V9(10) ;
  assign n154 = ~\V9(5)  & n153;
  assign n155 = ~\V9(6)  & n154;
  assign n156 = ~\V9(1)  & ~\V9(2) ;
  assign n157 = ~n152 & n156;
  assign n158 = \V9(1)  & ~\V9(10) ;
  assign n159 = \V9(8)  & n158;
  assign n160 = ~\V9(0)  & ~\V9(10) ;
  assign n161 = \V9(7)  & n160;
  assign n162 = ~\V9(5)  & n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = ~n159 & n163;
  assign n165 = ~n157 & n164;
  assign n166 = ~n155 & n165;
  assign n167 = ~\V9(1)  & ~\V9(10) ;
  assign n168 = \V9(0)  & n167;
  assign n169 = ~\V9(5)  & n168;
  assign n170 = ~\V9(6)  & n169;
  assign n171 = ~\V9(1)  & \V9(2) ;
  assign n172 = ~\V9(10)  & n171;
  assign n173 = \V9(8)  & n172;
  assign n174 = ~\V9(5)  & n156;
  assign n175 = ~\V9(6)  & n174;
  assign n176 = \V9(1)  & ~\V9(3) ;
  assign n177 = \V9(2)  & n176;
  assign n178 = ~\V9(10)  & n177;
  assign n179 = ~n157 & ~n178;
  assign n180 = ~n175 & n179;
  assign n181 = ~n173 & n180;
  assign n182 = ~n170 & n181;
  assign n183 = ~n166 & ~n182;
  assign n184 = n166 & n182;
  assign n185 = n166 & ~n182;
  assign n186 = ~n166 & n182;
  assign n187 = \V9(1)  & \V9(2) ;
  assign n188 = ~\V9(10)  & n184;
  assign n189 = ~n187 & n188;
  assign n190 = \V56(7)  & n183;
  assign n191 = \V56(22)  & n184;
  assign n192 = \V56(11)  & n185;
  assign n193 = \V56(14)  & n186;
  assign n194 = ~n189 & ~n193;
  assign n195 = ~n192 & n194;
  assign n196 = ~n191 & n195;
  assign \V119(21)  = n190 | ~n196;
  assign n198 = ~n166 & ~n186;
  assign n199 = n182 & ~n186;
  assign n200 = \V88(1)  & n198;
  assign n201 = \V88(16)  & n199;
  assign n202 = \V88(5)  & n185;
  assign n203 = \V88(8)  & n186;
  assign n204 = ~n189 & ~n203;
  assign n205 = ~n202 & n204;
  assign n206 = ~n201 & n205;
  assign \V151(16)  = n200 | ~n206;
  assign n208 = \V56(6)  & n183;
  assign n209 = \V56(21)  & n184;
  assign n210 = \V56(10)  & n185;
  assign n211 = \V56(13)  & n186;
  assign n212 = ~n189 & ~n211;
  assign n213 = ~n210 & n212;
  assign n214 = ~n209 & n213;
  assign \V119(20)  = n208 | ~n214;
  assign n216 = \V88(8)  & n185;
  assign n217 = ~n189 & ~n216;
  assign n218 = \V88(4)  & n198;
  assign n219 = \V88(19)  & n199;
  assign n220 = \V88(11)  & n186;
  assign n221 = n217 & ~n220;
  assign n222 = ~n219 & n221;
  assign \V151(19)  = n218 | ~n222;
  assign n224 = \V56(9)  & n183;
  assign n225 = \V56(24)  & n184;
  assign n226 = \V56(13)  & n185;
  assign n227 = \V56(16)  & n186;
  assign n228 = ~n189 & ~n227;
  assign n229 = ~n226 & n228;
  assign n230 = ~n225 & n229;
  assign \V119(23)  = n224 | ~n230;
  assign n232 = \V88(3)  & n198;
  assign n233 = \V88(18)  & n199;
  assign n234 = \V88(7)  & n185;
  assign n235 = \V88(10)  & n186;
  assign n236 = ~n189 & ~n235;
  assign n237 = ~n234 & n236;
  assign n238 = ~n233 & n237;
  assign \V151(18)  = n232 | ~n238;
  assign n240 = \V56(8)  & n183;
  assign n241 = \V56(23)  & n184;
  assign n242 = \V56(12)  & n185;
  assign n243 = \V56(15)  & n186;
  assign n244 = ~n189 & ~n243;
  assign n245 = ~n242 & n244;
  assign n246 = ~n241 & n245;
  assign \V119(22)  = n240 | ~n246;
  assign n248 = \V56(11)  & n183;
  assign n249 = \V56(26)  & n184;
  assign n250 = \V56(15)  & n185;
  assign n251 = \V56(18)  & n186;
  assign n252 = ~n189 & ~n251;
  assign n253 = ~n250 & n252;
  assign n254 = ~n249 & n253;
  assign \V119(25)  = n248 | ~n254;
  assign n256 = \V56(10)  & n183;
  assign n257 = \V56(25)  & n184;
  assign n258 = \V56(14)  & n185;
  assign n259 = \V56(17)  & n186;
  assign n260 = ~n189 & ~n259;
  assign n261 = ~n258 & n260;
  assign n262 = ~n257 & n261;
  assign \V119(24)  = n256 | ~n262;
  assign n264 = \V56(3)  & n183;
  assign n265 = \V56(18)  & n184;
  assign n266 = \V56(7)  & n185;
  assign n267 = \V56(10)  & n186;
  assign n268 = ~n189 & ~n267;
  assign n269 = ~n266 & n268;
  assign n270 = ~n265 & n269;
  assign \V119(17)  = n264 | ~n270;
  assign n272 = \V56(2)  & n183;
  assign n273 = \V56(17)  & n184;
  assign n274 = \V56(6)  & n185;
  assign n275 = \V56(9)  & n186;
  assign n276 = ~n189 & ~n275;
  assign n277 = ~n274 & n276;
  assign n278 = ~n273 & n277;
  assign \V119(16)  = n272 | ~n278;
  assign n280 = ~n186 & ~n189;
  assign n281 = \V88(4)  & n185;
  assign n282 = \V24(3)  & ~n166;
  assign n283 = \V56(4)  & n182;
  assign n284 = n280 & ~n283;
  assign n285 = ~n282 & n284;
  assign \V119(3)  = n281 | ~n285;
  assign n287 = \V56(5)  & n183;
  assign n288 = \V56(20)  & n184;
  assign n289 = \V56(9)  & n185;
  assign n290 = \V56(12)  & n186;
  assign n291 = ~n189 & ~n290;
  assign n292 = ~n289 & n291;
  assign n293 = ~n288 & n292;
  assign \V119(19)  = n287 | ~n293;
  assign n295 = \V88(3)  & n185;
  assign n296 = \V24(2)  & ~n166;
  assign n297 = \V56(3)  & n182;
  assign n298 = n280 & ~n297;
  assign n299 = ~n296 & n298;
  assign \V119(2)  = n295 | ~n299;
  assign n301 = \V56(4)  & n183;
  assign n302 = \V56(19)  & n184;
  assign n303 = \V56(8)  & n185;
  assign n304 = \V56(11)  & n186;
  assign n305 = ~n189 & ~n304;
  assign n306 = ~n303 & n305;
  assign n307 = ~n302 & n306;
  assign \V119(18)  = n301 | ~n307;
  assign n309 = \V56(28)  & n198;
  assign n310 = \V88(11)  & n199;
  assign n311 = \V88(0)  & n185;
  assign n312 = \V88(3)  & n186;
  assign n313 = ~n189 & ~n312;
  assign n314 = ~n311 & n313;
  assign n315 = ~n310 & n314;
  assign \V151(11)  = n309 | ~n315;
  assign n317 = \V88(6)  & n185;
  assign n318 = \V24(5)  & ~n166;
  assign n319 = \V56(6)  & n182;
  assign n320 = n280 & ~n319;
  assign n321 = ~n318 & n320;
  assign \V119(5)  = n317 | ~n321;
  assign n323 = \V56(27)  & n198;
  assign n324 = \V88(10)  & n199;
  assign n325 = \V56(31)  & n185;
  assign n326 = \V88(2)  & n186;
  assign n327 = ~n189 & ~n326;
  assign n328 = ~n325 & n327;
  assign n329 = ~n324 & n328;
  assign \V151(10)  = n323 | ~n329;
  assign n331 = \V24(4)  & ~n166;
  assign n332 = \V56(5)  & n182;
  assign n333 = n280 & ~n332;
  assign n334 = ~n331 & n333;
  assign \V119(4)  = n202 | ~n334;
  assign n336 = \V56(30)  & n198;
  assign n337 = \V88(13)  & n199;
  assign n338 = \V88(2)  & n185;
  assign n339 = \V88(5)  & n186;
  assign n340 = ~n189 & ~n339;
  assign n341 = ~n338 & n340;
  assign n342 = ~n337 & n341;
  assign \V151(13)  = n336 | ~n342;
  assign n344 = \V56(29)  & n198;
  assign n345 = \V88(12)  & n199;
  assign n346 = \V88(1)  & n185;
  assign n347 = \V88(4)  & n186;
  assign n348 = ~n189 & ~n347;
  assign n349 = ~n346 & n348;
  assign n350 = ~n345 & n349;
  assign \V151(12)  = n344 | ~n350;
  assign n352 = \V88(0)  & n198;
  assign n353 = \V88(15)  & n199;
  assign n354 = \V88(7)  & n186;
  assign n355 = ~n189 & ~n354;
  assign n356 = ~n281 & n355;
  assign n357 = ~n353 & n356;
  assign \V151(15)  = n352 | ~n357;
  assign n359 = \V24(1)  & ~n166;
  assign n360 = \V56(2)  & n182;
  assign n361 = n280 & ~n360;
  assign n362 = ~n359 & n361;
  assign \V119(1)  = n338 | ~n362;
  assign n364 = \V56(31)  & n198;
  assign n365 = \V88(14)  & n199;
  assign n366 = \V88(6)  & n186;
  assign n367 = ~n189 & ~n366;
  assign n368 = ~n295 & n367;
  assign n369 = ~n365 & n368;
  assign \V151(14)  = n364 | ~n369;
  assign n371 = \V24(0)  & ~n166;
  assign n372 = \V56(1)  & n182;
  assign n373 = n280 & ~n372;
  assign n374 = ~n371 & n373;
  assign \V119(0)  = n346 | ~n374;
  assign n376 = \V24(11)  & n183;
  assign n377 = \V56(12)  & n184;
  assign n378 = \V56(1)  & n185;
  assign n379 = \V56(4)  & n186;
  assign n380 = ~n189 & ~n379;
  assign n381 = ~n378 & n380;
  assign n382 = ~n377 & n381;
  assign \V119(11)  = n376 | ~n382;
  assign n384 = \V88(11)  & n185;
  assign n385 = ~n189 & ~n384;
  assign n386 = \V24(10)  & n183;
  assign n387 = \V56(3)  & n186;
  assign n388 = n385 & ~n387;
  assign n389 = \V56(11)  & n184;
  assign n390 = n388 & ~n389;
  assign \V119(10)  = n386 | ~n390;
  assign n392 = \V24(13)  & n183;
  assign n393 = \V56(14)  & n184;
  assign n394 = \V56(3)  & n185;
  assign n395 = \V56(6)  & n186;
  assign n396 = ~n189 & ~n395;
  assign n397 = ~n394 & n396;
  assign n398 = ~n393 & n397;
  assign \V119(13)  = n392 | ~n398;
  assign n400 = \V24(12)  & n183;
  assign n401 = \V56(13)  & n184;
  assign n402 = \V56(2)  & n185;
  assign n403 = \V56(5)  & n186;
  assign n404 = ~n189 & ~n403;
  assign n405 = ~n402 & n404;
  assign n406 = ~n401 & n405;
  assign \V119(12)  = n400 | ~n406;
  assign n408 = \V24(7)  & n183;
  assign n409 = \V56(0)  & n186;
  assign n410 = n217 & ~n409;
  assign n411 = \V56(8)  & n184;
  assign n412 = n410 & ~n411;
  assign \V119(7)  = n408 | ~n412;
  assign n414 = \V56(1)  & n183;
  assign n415 = \V56(16)  & n184;
  assign n416 = \V56(5)  & n185;
  assign n417 = \V56(8)  & n186;
  assign n418 = ~n189 & ~n417;
  assign n419 = ~n416 & n418;
  assign n420 = ~n415 & n419;
  assign \V119(15)  = n414 | ~n420;
  assign n422 = \V24(6)  & ~n166;
  assign n423 = \V56(7)  & n182;
  assign n424 = n280 & ~n423;
  assign n425 = ~n422 & n424;
  assign \V119(6)  = n234 | ~n425;
  assign n427 = \V24(14)  & n183;
  assign n428 = \V56(15)  & n184;
  assign n429 = \V56(4)  & n185;
  assign n430 = \V56(7)  & n186;
  assign n431 = ~n189 & ~n430;
  assign n432 = ~n429 & n431;
  assign n433 = ~n428 & n432;
  assign \V119(14)  = n427 | ~n433;
  assign n435 = \V88(10)  & n185;
  assign n436 = ~n189 & ~n435;
  assign n437 = \V24(9)  & n183;
  assign n438 = \V56(2)  & n186;
  assign n439 = n436 & ~n438;
  assign n440 = \V56(10)  & n184;
  assign n441 = n439 & ~n440;
  assign \V119(9)  = n437 | ~n441;
  assign n443 = \V88(9)  & n185;
  assign n444 = ~n189 & ~n443;
  assign n445 = \V24(8)  & n183;
  assign n446 = \V56(1)  & n186;
  assign n447 = n444 & ~n446;
  assign n448 = \V56(9)  & n184;
  assign n449 = n447 & ~n448;
  assign \V119(8)  = n445 | ~n449;
  assign n451 = \V56(20)  & n198;
  assign n452 = \V88(3)  & n199;
  assign n453 = \V56(24)  & n185;
  assign n454 = \V56(27)  & n186;
  assign n455 = ~n189 & ~n454;
  assign n456 = ~n453 & n455;
  assign n457 = ~n452 & n456;
  assign \V151(3)  = n451 | ~n457;
  assign n459 = \V56(19)  & n198;
  assign n460 = \V88(2)  & n199;
  assign n461 = \V56(23)  & n185;
  assign n462 = \V56(26)  & n186;
  assign n463 = ~n189 & ~n462;
  assign n464 = ~n461 & n463;
  assign n465 = ~n460 & n464;
  assign \V151(2)  = n459 | ~n465;
  assign n467 = \V56(22)  & n198;
  assign n468 = \V88(5)  & n199;
  assign n469 = \V56(26)  & n185;
  assign n470 = \V56(29)  & n186;
  assign n471 = ~n189 & ~n470;
  assign n472 = ~n469 & n471;
  assign n473 = ~n468 & n472;
  assign \V151(5)  = n467 | ~n473;
  assign n475 = \V56(21)  & n198;
  assign n476 = \V88(4)  & n199;
  assign n477 = \V56(25)  & n185;
  assign n478 = \V56(28)  & n186;
  assign n479 = ~n189 & ~n478;
  assign n480 = ~n477 & n479;
  assign n481 = ~n476 & n480;
  assign \V151(4)  = n475 | ~n481;
  assign n483 = \V56(18)  & n198;
  assign n484 = \V88(1)  & n199;
  assign n485 = \V56(22)  & n185;
  assign n486 = \V56(25)  & n186;
  assign n487 = ~n189 & ~n486;
  assign n488 = ~n485 & n487;
  assign n489 = ~n484 & n488;
  assign \V151(1)  = n483 | ~n489;
  assign n491 = \V56(17)  & n198;
  assign n492 = \V88(0)  & n199;
  assign n493 = \V56(21)  & n185;
  assign n494 = \V56(24)  & n186;
  assign n495 = ~n189 & ~n494;
  assign n496 = ~n493 & n495;
  assign n497 = ~n492 & n496;
  assign \V151(0)  = n491 | ~n497;
  assign n499 = \V56(24)  & n198;
  assign n500 = \V88(7)  & n199;
  assign n501 = \V56(28)  & n185;
  assign n502 = \V56(31)  & n186;
  assign n503 = ~n189 & ~n502;
  assign n504 = ~n501 & n503;
  assign n505 = ~n500 & n504;
  assign \V151(7)  = n499 | ~n505;
  assign n507 = \V56(23)  & n198;
  assign n508 = \V88(6)  & n199;
  assign n509 = \V56(27)  & n185;
  assign n510 = \V56(30)  & n186;
  assign n511 = ~n189 & ~n510;
  assign n512 = ~n509 & n511;
  assign n513 = ~n508 & n512;
  assign \V151(6)  = n507 | ~n513;
  assign n515 = \V56(26)  & n198;
  assign n516 = \V88(9)  & n199;
  assign n517 = \V56(30)  & n185;
  assign n518 = \V88(1)  & n186;
  assign n519 = ~n189 & ~n518;
  assign n520 = ~n517 & n519;
  assign n521 = ~n516 & n520;
  assign \V151(9)  = n515 | ~n521;
  assign n523 = \V56(25)  & n198;
  assign n524 = \V88(8)  & n199;
  assign n525 = \V56(29)  & n185;
  assign n526 = \V88(0)  & n186;
  assign n527 = ~n189 & ~n526;
  assign n528 = ~n525 & n527;
  assign n529 = ~n524 & n528;
  assign \V151(8)  = n523 | ~n529;
  assign n531 = \V88(16)  & n198;
  assign n532 = \V88(31)  & n199;
  assign n533 = \V88(20)  & n185;
  assign n534 = \V88(23)  & n186;
  assign n535 = ~n189 & ~n534;
  assign n536 = ~n533 & n535;
  assign n537 = ~n532 & n536;
  assign \V151(31)  = n531 | ~n537;
  assign n539 = \V88(15)  & n198;
  assign n540 = \V88(30)  & n199;
  assign n541 = \V88(19)  & n185;
  assign n542 = \V88(22)  & n186;
  assign n543 = ~n189 & ~n542;
  assign n544 = ~n541 & n543;
  assign n545 = ~n540 & n544;
  assign \V151(30)  = n539 | ~n545;
  assign n547 = \V56(16)  & n183;
  assign n548 = \V56(31)  & n184;
  assign n549 = \V56(20)  & n185;
  assign n550 = \V56(23)  & n186;
  assign n551 = ~n189 & ~n550;
  assign n552 = ~n549 & n551;
  assign n553 = ~n548 & n552;
  assign \V119(30)  = n547 | ~n553;
  assign n555 = \V88(12)  & n198;
  assign n556 = \V88(27)  & n199;
  assign n557 = \V88(16)  & n185;
  assign n558 = \V88(19)  & n186;
  assign n559 = ~n189 & ~n558;
  assign n560 = ~n557 & n559;
  assign n561 = ~n556 & n560;
  assign \V151(27)  = n555 | ~n561;
  assign n563 = \V88(11)  & n198;
  assign n564 = \V88(26)  & n199;
  assign n565 = \V88(15)  & n185;
  assign n566 = \V88(18)  & n186;
  assign n567 = ~n189 & ~n566;
  assign n568 = ~n565 & n567;
  assign n569 = ~n564 & n568;
  assign \V151(26)  = n563 | ~n569;
  assign n571 = \V88(14)  & n198;
  assign n572 = \V88(29)  & n199;
  assign n573 = \V88(18)  & n185;
  assign n574 = \V88(21)  & n186;
  assign n575 = ~n189 & ~n574;
  assign n576 = ~n573 & n575;
  assign n577 = ~n572 & n576;
  assign \V151(29)  = n571 | ~n577;
  assign n579 = \V88(13)  & n198;
  assign n580 = \V88(28)  & n199;
  assign n581 = \V88(17)  & n185;
  assign n582 = \V88(20)  & n186;
  assign n583 = ~n189 & ~n582;
  assign n584 = ~n581 & n583;
  assign n585 = ~n580 & n584;
  assign \V151(28)  = n579 | ~n585;
  assign n587 = \V56(13)  & n183;
  assign n588 = \V56(28)  & n184;
  assign n589 = \V56(17)  & n185;
  assign n590 = \V56(20)  & n186;
  assign n591 = ~n189 & ~n590;
  assign n592 = ~n589 & n591;
  assign n593 = ~n588 & n592;
  assign \V119(27)  = n587 | ~n593;
  assign n595 = \V56(12)  & n183;
  assign n596 = \V56(27)  & n184;
  assign n597 = \V56(16)  & n185;
  assign n598 = \V56(19)  & n186;
  assign n599 = ~n189 & ~n598;
  assign n600 = ~n597 & n599;
  assign n601 = ~n596 & n600;
  assign \V119(26)  = n595 | ~n601;
  assign n603 = \V56(15)  & n183;
  assign n604 = \V56(30)  & n184;
  assign n605 = \V56(19)  & n185;
  assign n606 = \V56(22)  & n186;
  assign n607 = ~n189 & ~n606;
  assign n608 = ~n605 & n607;
  assign n609 = ~n604 & n608;
  assign \V119(29)  = n603 | ~n609;
  assign n611 = \V56(14)  & n183;
  assign n612 = \V56(29)  & n184;
  assign n613 = \V56(18)  & n185;
  assign n614 = \V56(21)  & n186;
  assign n615 = ~n189 & ~n614;
  assign n616 = ~n613 & n615;
  assign n617 = ~n612 & n616;
  assign \V119(28)  = n611 | ~n617;
  assign n619 = \V88(6)  & n198;
  assign n620 = \V88(21)  & n199;
  assign n621 = \V88(13)  & n186;
  assign n622 = n436 & ~n621;
  assign n623 = ~n620 & n622;
  assign \V151(21)  = n619 | ~n623;
  assign n625 = \V88(5)  & n198;
  assign n626 = \V88(20)  & n199;
  assign n627 = \V88(12)  & n186;
  assign n628 = n444 & ~n627;
  assign n629 = ~n626 & n628;
  assign \V151(20)  = n625 | ~n629;
  assign n631 = \V88(8)  & n198;
  assign n632 = \V88(23)  & n199;
  assign n633 = \V88(12)  & n185;
  assign n634 = \V88(15)  & n186;
  assign n635 = ~n189 & ~n634;
  assign n636 = ~n633 & n635;
  assign n637 = ~n632 & n636;
  assign \V151(23)  = n631 | ~n637;
  assign n639 = \V88(7)  & n198;
  assign n640 = \V88(22)  & n199;
  assign n641 = \V88(14)  & n186;
  assign n642 = n385 & ~n641;
  assign n643 = ~n640 & n642;
  assign \V151(22)  = n639 | ~n643;
  assign n645 = \V88(10)  & n198;
  assign n646 = \V88(25)  & n199;
  assign n647 = \V88(14)  & n185;
  assign n648 = \V88(17)  & n186;
  assign n649 = ~n189 & ~n648;
  assign n650 = ~n647 & n649;
  assign n651 = ~n646 & n650;
  assign \V151(25)  = n645 | ~n651;
  assign n653 = \V88(9)  & n198;
  assign n654 = \V88(24)  & n199;
  assign n655 = \V88(13)  & n185;
  assign n656 = \V88(16)  & n186;
  assign n657 = ~n189 & ~n656;
  assign n658 = ~n655 & n657;
  assign n659 = ~n654 & n658;
  assign \V151(24)  = n653 | ~n659;
  assign n661 = \V88(2)  & n198;
  assign n662 = \V88(17)  & n199;
  assign n663 = \V88(9)  & n186;
  assign n664 = ~n189 & ~n663;
  assign n665 = ~n317 & n664;
  assign n666 = ~n662 & n665;
  assign \V151(17)  = n661 | ~n666;
endmodule


