// Benchmark "i7" written by ABC on Tue May 16 16:07:50 2017

module i7 ( 
    \V32(30) , \V199(1) , \V199(0) , \V128(21) , \V128(20) , \V192(31) ,
    \V128(23) , \V192(30) , \V128(22) , \V160(3) , \V128(25) , \V160(2) ,
    \V128(24) , \V160(5) , \V128(17) , \V160(4) , \V128(16) , \V128(19) ,
    \V128(18) , \V160(1) , \V160(0) , \V160(7) , \V128(11) , \V160(6) ,
    \V128(10) , \V160(9) , \V128(13) , \V160(8) , \V160(31) , \V128(12) ,
    \V160(30) , \V128(15) , \V128(3) , \V128(14) , \V128(2) , \V128(5) ,
    \V128(4) , \V128(1) , \V128(0) , \V32(0) , \V32(1) , \V32(2) ,
    \V32(3) , \V128(7) , \V32(4) , \V128(6) , \V32(5) , \V128(9) ,
    \V32(6) , \V128(8) , \V32(7) , \V32(8) , \V32(9) , \V96(0) , \V96(1) ,
    \V96(2) , \V96(3) , \V96(4) , \V96(13) , \V96(5) , \V128(31) ,
    \V96(12) , \V96(6) , \V128(30) , \V96(15) , \V96(7) , \V96(14) ,
    \V96(8) , \V96(9) , \V96(11) , \V96(10) , \V96(17) , \V96(16) ,
    \V96(19) , \V96(18) , \V96(23) , \V96(22) , \V64(13) , \V96(25) ,
    \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V192(27) , \V96(21) ,
    \V192(26) , \V96(20) , \V192(29) , \V64(11) , \V192(28) , \V64(10) ,
    \V192(3) , \V192(2) , \V192(5) , \V96(27) , \V192(4) , \V96(26) ,
    \V64(17) , \V96(29) , \V64(16) , \V96(28) , \V192(21) , \V64(19) ,
    \V192(1) , \V192(20) , \V64(18) , \V192(0) , \V192(23) , \V64(23) ,
    \V192(22) , \V64(22) , \V32(13) , \V192(25) , \V64(25) , \V32(12) ,
    \V192(24) , \V64(24) , \V32(15) , \V192(17) , \V192(7) , \V32(14) ,
    \V96(31) , \V192(16) , \V160(27) , \V192(6) , \V96(30) , \V192(19) ,
    \V64(21) , \V160(26) , \V192(9) , \V192(18) , \V64(20) , \V160(29) ,
    \V192(8) , \V32(11) , \V160(28) , \V32(10) , \V194(1) , \V194(0) ,
    \V64(27) , \V64(26) , \V32(17) , \V192(11) , \V64(29) , \V32(16) ,
    \V192(10) , \V64(28) , \V160(21) , \V32(19) , \V192(13) , \V160(20) ,
    \V32(18) , \V192(12) , \V160(23) , \V32(23) , \V64(0) , \V192(15) ,
    \V160(22) , \V195(0) , \V32(22) , \V64(1) , \V192(14) , \V160(25) ,
    \V32(25) , \V64(2) , \V160(24) , \V32(24) , \V64(3) , \V160(17) ,
    \V64(4) , \V64(31) , \V160(16) , \V64(5) , \V64(30) , \V160(19) ,
    \V32(21) , \V64(6) , \V160(18) , \V32(20) , \V64(7) , \V64(8) ,
    \V64(9) , \V32(27) , \V32(26) , \V160(11) , \V32(29) , \V160(10) ,
    \V32(28) , \V160(13) , \V160(12) , \V128(27) , \V160(15) , \V128(26) ,
    \V160(14) , \V128(29) , \V199(3) , \V128(28) , \V32(31) , \V199(4) ,
    \V259(27) , \V259(26) , \V259(29) , \V227(3) , \V259(28) , \V227(2) ,
    \V227(5) , \V227(4) , \V227(1) , \V227(0) , \V259(21) , \V259(20) ,
    \V259(23) , \V259(22) , \V259(25) , \V227(7) , \V259(24) , \V227(6) ,
    \V259(17) , \V227(9) , \V259(16) , \V227(8) , \V227(27) , \V259(19) ,
    \V227(26) , \V259(18) , \V259(11) , \V259(10) , \V227(21) , \V259(13) ,
    \V227(20) , \V259(12) , \V227(23) , \V266(3) , \V259(15) , \V227(22) ,
    \V266(2) , \V259(14) , \V227(25) , \V266(5) , \V227(24) , \V266(4) ,
    \V227(17) , \V227(16) , \V227(19) , \V266(1) , \V227(18) , \V266(0) ,
    \V266(6) , \V227(11) , \V227(10) , \V227(13) , \V227(12) , \V227(15) ,
    \V227(14) , \V259(31) , \V259(30) , \V259(3) , \V259(2) , \V259(5) ,
    \V259(4) , \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) ,
    \V259(8)   );
  input  \V32(30) , \V199(1) , \V199(0) , \V128(21) , \V128(20) ,
    \V192(31) , \V128(23) , \V192(30) , \V128(22) , \V160(3) , \V128(25) ,
    \V160(2) , \V128(24) , \V160(5) , \V128(17) , \V160(4) , \V128(16) ,
    \V128(19) , \V128(18) , \V160(1) , \V160(0) , \V160(7) , \V128(11) ,
    \V160(6) , \V128(10) , \V160(9) , \V128(13) , \V160(8) , \V160(31) ,
    \V128(12) , \V160(30) , \V128(15) , \V128(3) , \V128(14) , \V128(2) ,
    \V128(5) , \V128(4) , \V128(1) , \V128(0) , \V32(0) , \V32(1) ,
    \V32(2) , \V32(3) , \V128(7) , \V32(4) , \V128(6) , \V32(5) ,
    \V128(9) , \V32(6) , \V128(8) , \V32(7) , \V32(8) , \V32(9) , \V96(0) ,
    \V96(1) , \V96(2) , \V96(3) , \V96(4) , \V96(13) , \V96(5) ,
    \V128(31) , \V96(12) , \V96(6) , \V128(30) , \V96(15) , \V96(7) ,
    \V96(14) , \V96(8) , \V96(9) , \V96(11) , \V96(10) , \V96(17) ,
    \V96(16) , \V96(19) , \V96(18) , \V96(23) , \V96(22) , \V64(13) ,
    \V96(25) , \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V192(27) ,
    \V96(21) , \V192(26) , \V96(20) , \V192(29) , \V64(11) , \V192(28) ,
    \V64(10) , \V192(3) , \V192(2) , \V192(5) , \V96(27) , \V192(4) ,
    \V96(26) , \V64(17) , \V96(29) , \V64(16) , \V96(28) , \V192(21) ,
    \V64(19) , \V192(1) , \V192(20) , \V64(18) , \V192(0) , \V192(23) ,
    \V64(23) , \V192(22) , \V64(22) , \V32(13) , \V192(25) , \V64(25) ,
    \V32(12) , \V192(24) , \V64(24) , \V32(15) , \V192(17) , \V192(7) ,
    \V32(14) , \V96(31) , \V192(16) , \V160(27) , \V192(6) , \V96(30) ,
    \V192(19) , \V64(21) , \V160(26) , \V192(9) , \V192(18) , \V64(20) ,
    \V160(29) , \V192(8) , \V32(11) , \V160(28) , \V32(10) , \V194(1) ,
    \V194(0) , \V64(27) , \V64(26) , \V32(17) , \V192(11) , \V64(29) ,
    \V32(16) , \V192(10) , \V64(28) , \V160(21) , \V32(19) , \V192(13) ,
    \V160(20) , \V32(18) , \V192(12) , \V160(23) , \V32(23) , \V64(0) ,
    \V192(15) , \V160(22) , \V195(0) , \V32(22) , \V64(1) , \V192(14) ,
    \V160(25) , \V32(25) , \V64(2) , \V160(24) , \V32(24) , \V64(3) ,
    \V160(17) , \V64(4) , \V64(31) , \V160(16) , \V64(5) , \V64(30) ,
    \V160(19) , \V32(21) , \V64(6) , \V160(18) , \V32(20) , \V64(7) ,
    \V64(8) , \V64(9) , \V32(27) , \V32(26) , \V160(11) , \V32(29) ,
    \V160(10) , \V32(28) , \V160(13) , \V160(12) , \V128(27) , \V160(15) ,
    \V128(26) , \V160(14) , \V128(29) , \V199(3) , \V128(28) , \V32(31) ,
    \V199(4) ;
  output \V259(27) , \V259(26) , \V259(29) , \V227(3) , \V259(28) , \V227(2) ,
    \V227(5) , \V227(4) , \V227(1) , \V227(0) , \V259(21) , \V259(20) ,
    \V259(23) , \V259(22) , \V259(25) , \V227(7) , \V259(24) , \V227(6) ,
    \V259(17) , \V227(9) , \V259(16) , \V227(8) , \V227(27) , \V259(19) ,
    \V227(26) , \V259(18) , \V259(11) , \V259(10) , \V227(21) , \V259(13) ,
    \V227(20) , \V259(12) , \V227(23) , \V266(3) , \V259(15) , \V227(22) ,
    \V266(2) , \V259(14) , \V227(25) , \V266(5) , \V227(24) , \V266(4) ,
    \V227(17) , \V227(16) , \V227(19) , \V266(1) , \V227(18) , \V266(0) ,
    \V266(6) , \V227(11) , \V227(10) , \V227(13) , \V227(12) , \V227(15) ,
    \V227(14) , \V259(31) , \V259(30) , \V259(3) , \V259(2) , \V259(5) ,
    \V259(4) , \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) ,
    \V259(8) ;
  wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n282, n283, n284, n285, n286, n287, n288, n290, n291,
    n292, n293, n294, n295, n296, n298, n299, n300, n301, n302, n303, n305,
    n306, n307, n308, n309, n310, n311, n313, n314, n315, n316, n317, n318,
    n320, n321, n322, n323, n324, n325, n327, n328, n329, n330, n331, n332,
    n334, n335, n336, n337, n338, n339, n341, n342, n343, n344, n345, n346,
    n348, n349, n350, n351, n352, n353, n354, n356, n357, n358, n359, n360,
    n361, n362, n364, n365, n366, n367, n368, n369, n370, n372, n373, n374,
    n375, n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n388,
    n389, n390, n391, n392, n393, n395, n396, n397, n398, n399, n400, n401,
    n403, n404, n405, n406, n407, n408, n410, n411, n412, n413, n414, n415,
    n416, n418, n419, n420, n421, n422, n423, n425, n426, n427, n428, n429,
    n430, n431, n433, n434, n435, n436, n437, n438, n440, n441, n442, n443,
    n444, n445, n447, n448, n449, n450, n451, n452, n453, n455, n456, n457,
    n458, n459, n460, n462, n463, n464, n465, n466, n467, n468, n470, n471,
    n472, n473, n474, n475, n476, n478, n479, n480, n481, n482, n483, n484,
    n486, n487, n488, n489, n490, n491, n493, n494, n495, n496, n497, n498,
    n499, n501, n502, n503, n504, n505, n506, n508, n509, n510, n511, n512,
    n513, n514, n516, n517, n518, n519, n520, n521, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n534, n535, n536, n537, n538, n539,
    n540, n542, n543, n544, n545, n546, n547, n549, n550, n551, n552, n553,
    n554, n555, n557, n558, n559, n560, n561, n562, n563, n565, n566, n567,
    n568, n569, n570, n572, n573, n574, n575, n577, n578, n579, n580, n581,
    n582, n584, n585, n586, n588, n589, n590, n591, n592, n593, n595, n596,
    n597, n598, n599, n600, n602, n603, n604, n605, n606, n607, n609, n610,
    n611, n612, n613, n614, n615, n617, n618, n619, n620, n621, n622, n624,
    n625, n626, n627, n628, n629, n630, n632, n634, n635, n636, n637, n638,
    n639, n641, n642, n643, n644, n645, n646, n648, n649, n650, n651, n652,
    n653, n655, n656, n657, n658, n659, n660, n662, n663, n664, n665, n666,
    n667, n669, n670, n671, n672, n673, n674, n676, n677, n678, n679, n680,
    n681, n682, n684, n685, n686, n687, n688, n689, n690, n692, n693, n694,
    n695, n696, n697, n698, n700, n701, n702, n703, n704, n705, n706, n708,
    n709, n710, n711, n712, n713, n714, n716, n717, n718, n719, n720, n721,
    n722, n724, n725, n726, n727, n728, n729, n730, n732, n733, n734, n735,
    n736, n737, n738, n740, n741, n742, n743, n744, n745, n746, n748, n749,
    n750, n751, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762,
    n764, n765, n766, n767, n768, n769, n770;
  assign n267 = ~\V199(1)  & ~\V199(0) ;
  assign n268 = \V199(4)  & n267;
  assign n269 = ~\V199(1)  & \V199(0) ;
  assign n270 = \V199(4)  & n269;
  assign n271 = \V199(1)  & \V199(0) ;
  assign n272 = \V199(1)  & ~\V199(0) ;
  assign n273 = \V199(1)  & ~\V199(4) ;
  assign n274 = \V192(23)  & n268;
  assign n275 = \V128(23)  & n270;
  assign n276 = \V160(23)  & n271;
  assign n277 = ~\V192(23)  & n272;
  assign n278 = ~n273 & ~n277;
  assign n279 = ~n276 & n278;
  assign n280 = ~n275 & n279;
  assign \V259(27)  = n274 | ~n280;
  assign n282 = \V192(22)  & n268;
  assign n283 = \V128(22)  & n270;
  assign n284 = \V160(22)  & n271;
  assign n285 = ~\V192(22)  & n272;
  assign n286 = ~n273 & ~n285;
  assign n287 = ~n284 & n286;
  assign n288 = ~n283 & n287;
  assign \V259(26)  = n282 | ~n288;
  assign n290 = \V192(25)  & n268;
  assign n291 = \V128(25)  & n270;
  assign n292 = \V160(25)  & n271;
  assign n293 = ~\V192(25)  & n272;
  assign n294 = ~n273 & ~n293;
  assign n295 = ~n292 & n294;
  assign n296 = ~n291 & n295;
  assign \V259(29)  = n290 | ~n296;
  assign n298 = \V64(3)  & n271;
  assign n299 = \V32(3)  & n269;
  assign n300 = \V96(3)  & n267;
  assign n301 = ~\V96(3)  & n272;
  assign n302 = ~n300 & ~n301;
  assign n303 = ~n299 & n302;
  assign \V227(3)  = n298 | ~n303;
  assign n305 = \V192(24)  & n268;
  assign n306 = \V128(24)  & n270;
  assign n307 = \V160(24)  & n271;
  assign n308 = ~\V192(24)  & n272;
  assign n309 = ~n273 & ~n308;
  assign n310 = ~n307 & n309;
  assign n311 = ~n306 & n310;
  assign \V259(28)  = n305 | ~n311;
  assign n313 = \V64(2)  & n271;
  assign n314 = \V32(2)  & n269;
  assign n315 = \V96(2)  & n267;
  assign n316 = ~\V96(2)  & n272;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~n314 & n317;
  assign \V227(2)  = n313 | ~n318;
  assign n320 = \V64(5)  & n271;
  assign n321 = \V32(5)  & n269;
  assign n322 = \V96(5)  & n267;
  assign n323 = ~\V96(5)  & n272;
  assign n324 = ~n322 & ~n323;
  assign n325 = ~n321 & n324;
  assign \V227(5)  = n320 | ~n325;
  assign n327 = \V64(4)  & n271;
  assign n328 = \V32(4)  & n269;
  assign n329 = \V96(4)  & n267;
  assign n330 = ~\V96(4)  & n272;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n328 & n331;
  assign \V227(4)  = n327 | ~n332;
  assign n334 = \V64(1)  & n271;
  assign n335 = \V32(1)  & n269;
  assign n336 = \V96(1)  & n267;
  assign n337 = ~\V96(1)  & n272;
  assign n338 = ~n336 & ~n337;
  assign n339 = ~n335 & n338;
  assign \V227(1)  = n334 | ~n339;
  assign n341 = \V64(0)  & n271;
  assign n342 = \V32(0)  & n269;
  assign n343 = \V96(0)  & n267;
  assign n344 = ~\V96(0)  & n272;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~n342 & n345;
  assign \V227(0)  = n341 | ~n346;
  assign n348 = \V192(17)  & n268;
  assign n349 = \V128(17)  & n270;
  assign n350 = \V160(17)  & n271;
  assign n351 = ~\V192(17)  & n272;
  assign n352 = ~n273 & ~n351;
  assign n353 = ~n350 & n352;
  assign n354 = ~n349 & n353;
  assign \V259(21)  = n348 | ~n354;
  assign n356 = \V192(16)  & n268;
  assign n357 = \V128(16)  & n270;
  assign n358 = \V160(16)  & n271;
  assign n359 = ~\V192(16)  & n272;
  assign n360 = ~n273 & ~n359;
  assign n361 = ~n358 & n360;
  assign n362 = ~n357 & n361;
  assign \V259(20)  = n356 | ~n362;
  assign n364 = \V192(19)  & n268;
  assign n365 = \V128(19)  & n270;
  assign n366 = \V160(19)  & n271;
  assign n367 = ~\V192(19)  & n272;
  assign n368 = ~n273 & ~n367;
  assign n369 = ~n366 & n368;
  assign n370 = ~n365 & n369;
  assign \V259(23)  = n364 | ~n370;
  assign n372 = \V192(18)  & n268;
  assign n373 = \V128(18)  & n270;
  assign n374 = \V160(18)  & n271;
  assign n375 = ~\V192(18)  & n272;
  assign n376 = ~n273 & ~n375;
  assign n377 = ~n374 & n376;
  assign n378 = ~n373 & n377;
  assign \V259(22)  = n372 | ~n378;
  assign n380 = \V192(21)  & n268;
  assign n381 = \V128(21)  & n270;
  assign n382 = \V160(21)  & n271;
  assign n383 = ~\V192(21)  & n272;
  assign n384 = ~n273 & ~n383;
  assign n385 = ~n382 & n384;
  assign n386 = ~n381 & n385;
  assign \V259(25)  = n380 | ~n386;
  assign n388 = \V64(7)  & n271;
  assign n389 = \V32(7)  & n269;
  assign n390 = \V96(7)  & n267;
  assign n391 = ~\V96(7)  & n272;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n389 & n392;
  assign \V227(7)  = n388 | ~n393;
  assign n395 = \V192(20)  & n268;
  assign n396 = \V128(20)  & n270;
  assign n397 = \V160(20)  & n271;
  assign n398 = ~\V192(20)  & n272;
  assign n399 = ~n273 & ~n398;
  assign n400 = ~n397 & n399;
  assign n401 = ~n396 & n400;
  assign \V259(24)  = n395 | ~n401;
  assign n403 = \V64(6)  & n271;
  assign n404 = \V32(6)  & n269;
  assign n405 = \V96(6)  & n267;
  assign n406 = ~\V96(6)  & n272;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n404 & n407;
  assign \V227(6)  = n403 | ~n408;
  assign n410 = \V192(13)  & n268;
  assign n411 = \V128(13)  & n270;
  assign n412 = \V160(13)  & n271;
  assign n413 = ~\V192(13)  & n272;
  assign n414 = ~n273 & ~n413;
  assign n415 = ~n412 & n414;
  assign n416 = ~n411 & n415;
  assign \V259(17)  = n410 | ~n416;
  assign n418 = \V64(9)  & n271;
  assign n419 = \V32(9)  & n269;
  assign n420 = \V96(9)  & n267;
  assign n421 = ~\V96(9)  & n272;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~n419 & n422;
  assign \V227(9)  = n418 | ~n423;
  assign n425 = \V192(12)  & n268;
  assign n426 = \V128(12)  & n270;
  assign n427 = \V160(12)  & n271;
  assign n428 = ~\V192(12)  & n272;
  assign n429 = ~n273 & ~n428;
  assign n430 = ~n427 & n429;
  assign n431 = ~n426 & n430;
  assign \V259(16)  = n425 | ~n431;
  assign n433 = \V64(8)  & n271;
  assign n434 = \V32(8)  & n269;
  assign n435 = \V96(8)  & n267;
  assign n436 = ~\V96(8)  & n272;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n434 & n437;
  assign \V227(8)  = n433 | ~n438;
  assign n440 = \V64(27)  & n271;
  assign n441 = \V32(27)  & n269;
  assign n442 = \V96(27)  & n267;
  assign n443 = ~\V96(27)  & n272;
  assign n444 = ~n442 & ~n443;
  assign n445 = ~n441 & n444;
  assign \V227(27)  = n440 | ~n445;
  assign n447 = \V192(15)  & n268;
  assign n448 = \V128(15)  & n270;
  assign n449 = \V160(15)  & n271;
  assign n450 = ~\V192(15)  & n272;
  assign n451 = ~n273 & ~n450;
  assign n452 = ~n449 & n451;
  assign n453 = ~n448 & n452;
  assign \V259(19)  = n447 | ~n453;
  assign n455 = \V64(26)  & n271;
  assign n456 = \V32(26)  & n269;
  assign n457 = \V96(26)  & n267;
  assign n458 = ~\V96(26)  & n272;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~n456 & n459;
  assign \V227(26)  = n455 | ~n460;
  assign n462 = \V192(14)  & n268;
  assign n463 = \V128(14)  & n270;
  assign n464 = \V160(14)  & n271;
  assign n465 = ~\V192(14)  & n272;
  assign n466 = ~n273 & ~n465;
  assign n467 = ~n464 & n466;
  assign n468 = ~n463 & n467;
  assign \V259(18)  = n462 | ~n468;
  assign n470 = \V192(7)  & n268;
  assign n471 = \V128(7)  & n270;
  assign n472 = \V160(7)  & n271;
  assign n473 = ~\V192(7)  & n272;
  assign n474 = ~n273 & ~n473;
  assign n475 = ~n472 & n474;
  assign n476 = ~n471 & n475;
  assign \V259(11)  = n470 | ~n476;
  assign n478 = \V192(6)  & n268;
  assign n479 = \V128(6)  & n270;
  assign n480 = \V160(6)  & n271;
  assign n481 = ~\V192(6)  & n272;
  assign n482 = ~n273 & ~n481;
  assign n483 = ~n480 & n482;
  assign n484 = ~n479 & n483;
  assign \V259(10)  = n478 | ~n484;
  assign n486 = \V64(21)  & n271;
  assign n487 = \V32(21)  & n269;
  assign n488 = \V96(21)  & n267;
  assign n489 = ~\V96(21)  & n272;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n487 & n490;
  assign \V227(21)  = n486 | ~n491;
  assign n493 = \V192(9)  & n268;
  assign n494 = \V128(9)  & n270;
  assign n495 = \V160(9)  & n271;
  assign n496 = ~\V192(9)  & n272;
  assign n497 = ~n273 & ~n496;
  assign n498 = ~n495 & n497;
  assign n499 = ~n494 & n498;
  assign \V259(13)  = n493 | ~n499;
  assign n501 = \V64(20)  & n271;
  assign n502 = \V32(20)  & n269;
  assign n503 = \V96(20)  & n267;
  assign n504 = ~\V96(20)  & n272;
  assign n505 = ~n503 & ~n504;
  assign n506 = ~n502 & n505;
  assign \V227(20)  = n501 | ~n506;
  assign n508 = \V192(8)  & n268;
  assign n509 = \V128(8)  & n270;
  assign n510 = \V160(8)  & n271;
  assign n511 = ~\V192(8)  & n272;
  assign n512 = ~n273 & ~n511;
  assign n513 = ~n510 & n512;
  assign n514 = ~n509 & n513;
  assign \V259(12)  = n508 | ~n514;
  assign n516 = \V64(23)  & n271;
  assign n517 = \V32(23)  & n269;
  assign n518 = \V96(23)  & n267;
  assign n519 = ~\V96(23)  & n272;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n517 & n520;
  assign \V227(23)  = n516 | ~n521;
  assign n523 = \V199(3)  & n269;
  assign n524 = \V199(3)  & n267;
  assign n525 = \V199(1)  & ~\V199(3) ;
  assign n526 = \V128(31)  & n523;
  assign n527 = \V192(31)  & n524;
  assign n528 = ~\V192(31)  & n272;
  assign n529 = \V160(31)  & n271;
  assign n530 = ~n525 & ~n529;
  assign n531 = ~n528 & n530;
  assign n532 = ~n527 & n531;
  assign \V266(3)  = n526 | ~n532;
  assign n534 = \V192(11)  & n268;
  assign n535 = \V128(11)  & n270;
  assign n536 = \V160(11)  & n271;
  assign n537 = ~\V192(11)  & n272;
  assign n538 = ~n273 & ~n537;
  assign n539 = ~n536 & n538;
  assign n540 = ~n535 & n539;
  assign \V259(15)  = n534 | ~n540;
  assign n542 = \V64(22)  & n271;
  assign n543 = \V32(22)  & n269;
  assign n544 = \V96(22)  & n267;
  assign n545 = ~\V96(22)  & n272;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n543 & n546;
  assign \V227(22)  = n542 | ~n547;
  assign n549 = \V128(30)  & n523;
  assign n550 = \V192(30)  & n524;
  assign n551 = ~\V192(30)  & n272;
  assign n552 = \V160(30)  & n271;
  assign n553 = ~n525 & ~n552;
  assign n554 = ~n551 & n553;
  assign n555 = ~n550 & n554;
  assign \V266(2)  = n549 | ~n555;
  assign n557 = \V192(10)  & n268;
  assign n558 = \V128(10)  & n270;
  assign n559 = \V160(10)  & n271;
  assign n560 = ~\V192(10)  & n272;
  assign n561 = ~n273 & ~n560;
  assign n562 = ~n559 & n561;
  assign n563 = ~n558 & n562;
  assign \V259(14)  = n557 | ~n563;
  assign n565 = \V64(25)  & n271;
  assign n566 = \V32(25)  & n269;
  assign n567 = \V96(25)  & n267;
  assign n568 = ~\V96(25)  & n272;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n566 & n569;
  assign \V227(25)  = n565 | ~n570;
  assign n572 = \V194(1)  & n524;
  assign n573 = \V199(1)  & ~\V194(1) ;
  assign n574 = ~n271 & ~n525;
  assign n575 = ~n573 & n574;
  assign \V266(5)  = n572 | ~n575;
  assign n577 = \V64(24)  & n271;
  assign n578 = \V32(24)  & n269;
  assign n579 = \V96(24)  & n267;
  assign n580 = ~\V96(24)  & n272;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n578 & n581;
  assign \V227(24)  = n577 | ~n582;
  assign n584 = \V194(0)  & n524;
  assign n585 = \V199(1)  & ~\V194(0) ;
  assign n586 = n574 & ~n585;
  assign \V266(4)  = n584 | ~n586;
  assign n588 = \V64(17)  & n271;
  assign n589 = \V32(17)  & n269;
  assign n590 = \V96(17)  & n267;
  assign n591 = ~\V96(17)  & n272;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n589 & n592;
  assign \V227(17)  = n588 | ~n593;
  assign n595 = \V64(16)  & n271;
  assign n596 = \V32(16)  & n269;
  assign n597 = \V96(16)  & n267;
  assign n598 = ~\V96(16)  & n272;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n596 & n599;
  assign \V227(16)  = n595 | ~n600;
  assign n602 = \V64(19)  & n271;
  assign n603 = \V32(19)  & n269;
  assign n604 = \V96(19)  & n267;
  assign n605 = ~\V96(19)  & n272;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n603 & n606;
  assign \V227(19)  = n602 | ~n607;
  assign n609 = \V128(29)  & n523;
  assign n610 = \V192(29)  & n524;
  assign n611 = ~\V192(29)  & n272;
  assign n612 = \V160(29)  & n271;
  assign n613 = ~n525 & ~n612;
  assign n614 = ~n611 & n613;
  assign n615 = ~n610 & n614;
  assign \V266(1)  = n609 | ~n615;
  assign n617 = \V64(18)  & n271;
  assign n618 = \V32(18)  & n269;
  assign n619 = \V96(18)  & n267;
  assign n620 = ~\V96(18)  & n272;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n618 & n621;
  assign \V227(18)  = n617 | ~n622;
  assign n624 = \V128(28)  & n523;
  assign n625 = \V192(28)  & n524;
  assign n626 = ~\V192(28)  & n272;
  assign n627 = \V160(28)  & n271;
  assign n628 = ~n525 & ~n627;
  assign n629 = ~n626 & n628;
  assign n630 = ~n625 & n629;
  assign \V266(0)  = n624 | ~n630;
  assign n632 = ~\V199(0)  & \V199(3) ;
  assign \V266(6)  = \V195(0)  & n632;
  assign n634 = \V64(11)  & n271;
  assign n635 = \V32(11)  & n269;
  assign n636 = \V96(11)  & n267;
  assign n637 = ~\V96(11)  & n272;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~n635 & n638;
  assign \V227(11)  = n634 | ~n639;
  assign n641 = \V64(10)  & n271;
  assign n642 = \V32(10)  & n269;
  assign n643 = \V96(10)  & n267;
  assign n644 = ~\V96(10)  & n272;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~n642 & n645;
  assign \V227(10)  = n641 | ~n646;
  assign n648 = \V64(13)  & n271;
  assign n649 = \V32(13)  & n269;
  assign n650 = \V96(13)  & n267;
  assign n651 = ~\V96(13)  & n272;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n649 & n652;
  assign \V227(13)  = n648 | ~n653;
  assign n655 = \V64(12)  & n271;
  assign n656 = \V32(12)  & n269;
  assign n657 = \V96(12)  & n267;
  assign n658 = ~\V96(12)  & n272;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n656 & n659;
  assign \V227(12)  = n655 | ~n660;
  assign n662 = \V64(15)  & n271;
  assign n663 = \V32(15)  & n269;
  assign n664 = \V96(15)  & n267;
  assign n665 = ~\V96(15)  & n272;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~n663 & n666;
  assign \V227(15)  = n662 | ~n667;
  assign n669 = \V64(14)  & n271;
  assign n670 = \V32(14)  & n269;
  assign n671 = \V96(14)  & n267;
  assign n672 = ~\V96(14)  & n272;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n670 & n673;
  assign \V227(14)  = n669 | ~n674;
  assign n676 = \V192(27)  & n268;
  assign n677 = \V128(27)  & n270;
  assign n678 = \V160(27)  & n271;
  assign n679 = ~\V192(27)  & n272;
  assign n680 = ~n273 & ~n679;
  assign n681 = ~n678 & n680;
  assign n682 = ~n677 & n681;
  assign \V259(31)  = n676 | ~n682;
  assign n684 = \V192(26)  & n268;
  assign n685 = \V128(26)  & n270;
  assign n686 = \V160(26)  & n271;
  assign n687 = ~\V192(26)  & n272;
  assign n688 = ~n273 & ~n687;
  assign n689 = ~n686 & n688;
  assign n690 = ~n685 & n689;
  assign \V259(30)  = n684 | ~n690;
  assign n692 = \V96(31)  & n268;
  assign n693 = \V32(31)  & n270;
  assign n694 = \V64(31)  & n271;
  assign n695 = ~\V96(31)  & n272;
  assign n696 = ~n273 & ~n695;
  assign n697 = ~n694 & n696;
  assign n698 = ~n693 & n697;
  assign \V259(3)  = n692 | ~n698;
  assign n700 = \V96(30)  & n268;
  assign n701 = \V32(30)  & n270;
  assign n702 = \V64(30)  & n271;
  assign n703 = ~\V96(30)  & n272;
  assign n704 = ~n273 & ~n703;
  assign n705 = ~n702 & n704;
  assign n706 = ~n701 & n705;
  assign \V259(2)  = n700 | ~n706;
  assign n708 = \V192(1)  & n268;
  assign n709 = \V128(1)  & n270;
  assign n710 = \V160(1)  & n271;
  assign n711 = ~\V192(1)  & n272;
  assign n712 = ~n273 & ~n711;
  assign n713 = ~n710 & n712;
  assign n714 = ~n709 & n713;
  assign \V259(5)  = n708 | ~n714;
  assign n716 = \V192(0)  & n268;
  assign n717 = \V128(0)  & n270;
  assign n718 = \V160(0)  & n271;
  assign n719 = ~\V192(0)  & n272;
  assign n720 = ~n273 & ~n719;
  assign n721 = ~n718 & n720;
  assign n722 = ~n717 & n721;
  assign \V259(4)  = n716 | ~n722;
  assign n724 = \V96(29)  & n268;
  assign n725 = \V32(29)  & n270;
  assign n726 = \V64(29)  & n271;
  assign n727 = ~\V96(29)  & n272;
  assign n728 = ~n273 & ~n727;
  assign n729 = ~n726 & n728;
  assign n730 = ~n725 & n729;
  assign \V259(1)  = n724 | ~n730;
  assign n732 = \V96(28)  & n268;
  assign n733 = \V32(28)  & n270;
  assign n734 = \V64(28)  & n271;
  assign n735 = ~\V96(28)  & n272;
  assign n736 = ~n273 & ~n735;
  assign n737 = ~n734 & n736;
  assign n738 = ~n733 & n737;
  assign \V259(0)  = n732 | ~n738;
  assign n740 = \V192(3)  & n268;
  assign n741 = \V128(3)  & n270;
  assign n742 = \V160(3)  & n271;
  assign n743 = ~\V192(3)  & n272;
  assign n744 = ~n273 & ~n743;
  assign n745 = ~n742 & n744;
  assign n746 = ~n741 & n745;
  assign \V259(7)  = n740 | ~n746;
  assign n748 = \V192(2)  & n268;
  assign n749 = \V128(2)  & n270;
  assign n750 = \V160(2)  & n271;
  assign n751 = ~\V192(2)  & n272;
  assign n752 = ~n273 & ~n751;
  assign n753 = ~n750 & n752;
  assign n754 = ~n749 & n753;
  assign \V259(6)  = n748 | ~n754;
  assign n756 = \V192(5)  & n268;
  assign n757 = \V128(5)  & n270;
  assign n758 = \V160(5)  & n271;
  assign n759 = ~\V192(5)  & n272;
  assign n760 = ~n273 & ~n759;
  assign n761 = ~n758 & n760;
  assign n762 = ~n757 & n761;
  assign \V259(9)  = n756 | ~n762;
  assign n764 = \V192(4)  & n268;
  assign n765 = \V128(4)  & n270;
  assign n766 = \V160(4)  & n271;
  assign n767 = ~\V192(4)  & n272;
  assign n768 = ~n273 & ~n767;
  assign n769 = ~n766 & n768;
  assign n770 = ~n765 & n769;
  assign \V259(8)  = n764 | ~n770;
endmodule


