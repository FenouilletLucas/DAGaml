// Benchmark "i7" written by ABC on Tue May 16 16:07:50 2017

module i7 ( 
    \V160(21) , \V160(20) , \V160(23) , \V160(22) , \V128(27) , \V160(25) ,
    \V128(26) , \V160(24) , \V128(29) , \V160(17) , \V128(28) , \V160(16) ,
    \V160(19) , \V160(18) , \V96(0) , \V96(1) , \V64(13) , \V96(2) ,
    \V64(12) , \V96(3) , \V64(15) , \V128(21) , \V96(4) , \V64(14) ,
    \V128(20) , \V96(5) , \V128(23) , \V160(11) , \V96(6) , \V128(22) ,
    \V160(10) , \V96(7) , \V64(11) , \V128(25) , \V160(13) , \V96(8) ,
    \V64(10) , \V128(24) , \V192(3) , \V160(12) , \V96(9) , \V128(17) ,
    \V192(2) , \V160(15) , \V128(16) , \V192(5) , \V160(14) , \V128(19) ,
    \V192(4) , \V128(18) , \V64(17) , \V64(16) , \V192(1) , \V64(19) ,
    \V192(0) , \V64(18) , \V64(23) , \V64(22) , \V64(25) , \V128(11) ,
    \V64(24) , \V128(10) , \V192(7) , \V128(13) , \V192(6) , \V128(12) ,
    \V192(9) , \V64(21) , \V128(15) , \V192(8) , \V64(20) , \V128(14) ,
    \V64(27) , \V64(26) , \V64(29) , \V64(28) , \V194(1) , \V160(31) ,
    \V194(0) , \V160(30) , \V64(31) , \V64(30) , \V128(3) , \V128(2) ,
    \V128(5) , \V195(0) , \V128(4) , \V128(31) , \V128(30) , \V128(1) ,
    \V128(0) , \V128(7) , \V128(6) , \V128(9) , \V128(8) , \V199(3) ,
    \V199(4) , \V199(1) , \V199(0) , \V32(0) , \V32(1) , \V32(2) ,
    \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) , \V32(15) ,
    \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) , \V32(11) ,
    \V32(10) , \V192(27) , \V192(26) , \V192(29) , \V192(28) , \V32(17) ,
    \V32(16) , \V32(19) , \V32(18) , \V32(23) , \V32(22) , \V192(21) ,
    \V32(25) , \V192(20) , \V32(24) , \V192(23) , \V192(22) , \V192(25) ,
    \V32(21) , \V192(24) , \V32(20) , \V192(17) , \V192(16) , \V192(19) ,
    \V192(18) , \V32(27) , \V96(13) , \V32(26) , \V96(12) , \V32(29) ,
    \V96(15) , \V32(28) , \V96(14) , \V192(11) , \V192(10) , \V96(11) ,
    \V192(13) , \V96(10) , \V192(12) , \V192(15) , \V32(31) , \V192(14) ,
    \V32(30) , \V96(17) , \V96(16) , \V96(19) , \V96(18) , \V96(23) ,
    \V96(22) , \V96(25) , \V96(24) , \V96(21) , \V96(20) , \V96(27) ,
    \V96(26) , \V96(29) , \V96(28) , \V192(31) , \V64(0) , \V192(30) ,
    \V96(31) , \V64(1) , \V96(30) , \V64(2) , \V64(3) , \V64(4) , \V64(5) ,
    \V64(6) , \V64(7) , \V64(8) , \V160(3) , \V64(9) , \V160(2) ,
    \V160(5) , \V160(4) , \V160(1) , \V160(0) , \V160(7) , \V160(6) ,
    \V160(9) , \V160(8) , \V160(27) , \V160(26) , \V160(29) , \V160(28) ,
    \V259(27) , \V259(26) , \V259(29) , \V259(28) , \V259(21) , \V259(20) ,
    \V259(23) , \V259(22) , \V259(25) , \V259(24) , \V259(17) , \V259(16) ,
    \V259(19) , \V259(18) , \V259(11) , \V259(10) , \V259(13) , \V259(12) ,
    \V259(15) , \V259(14) , \V259(3) , \V259(2) , \V259(5) , \V259(4) ,
    \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) , \V259(8) ,
    \V259(31) , \V259(30) , \V227(27) , \V227(26) , \V227(21) , \V227(20) ,
    \V227(23) , \V227(22) , \V227(25) , \V227(24) , \V227(17) , \V227(16) ,
    \V227(19) , \V227(18) , \V227(11) , \V227(10) , \V227(13) , \V227(12) ,
    \V227(15) , \V227(14) , \V266(3) , \V266(2) , \V266(5) , \V266(4) ,
    \V266(1) , \V266(0) , \V266(6) , \V227(3) , \V227(2) , \V227(5) ,
    \V227(4) , \V227(1) , \V227(0) , \V227(7) , \V227(6) , \V227(9) ,
    \V227(8)   );
  input  \V160(21) , \V160(20) , \V160(23) , \V160(22) , \V128(27) ,
    \V160(25) , \V128(26) , \V160(24) , \V128(29) , \V160(17) , \V128(28) ,
    \V160(16) , \V160(19) , \V160(18) , \V96(0) , \V96(1) , \V64(13) ,
    \V96(2) , \V64(12) , \V96(3) , \V64(15) , \V128(21) , \V96(4) ,
    \V64(14) , \V128(20) , \V96(5) , \V128(23) , \V160(11) , \V96(6) ,
    \V128(22) , \V160(10) , \V96(7) , \V64(11) , \V128(25) , \V160(13) ,
    \V96(8) , \V64(10) , \V128(24) , \V192(3) , \V160(12) , \V96(9) ,
    \V128(17) , \V192(2) , \V160(15) , \V128(16) , \V192(5) , \V160(14) ,
    \V128(19) , \V192(4) , \V128(18) , \V64(17) , \V64(16) , \V192(1) ,
    \V64(19) , \V192(0) , \V64(18) , \V64(23) , \V64(22) , \V64(25) ,
    \V128(11) , \V64(24) , \V128(10) , \V192(7) , \V128(13) , \V192(6) ,
    \V128(12) , \V192(9) , \V64(21) , \V128(15) , \V192(8) , \V64(20) ,
    \V128(14) , \V64(27) , \V64(26) , \V64(29) , \V64(28) , \V194(1) ,
    \V160(31) , \V194(0) , \V160(30) , \V64(31) , \V64(30) , \V128(3) ,
    \V128(2) , \V128(5) , \V195(0) , \V128(4) , \V128(31) , \V128(30) ,
    \V128(1) , \V128(0) , \V128(7) , \V128(6) , \V128(9) , \V128(8) ,
    \V199(3) , \V199(4) , \V199(1) , \V199(0) , \V32(0) , \V32(1) ,
    \V32(2) , \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) ,
    \V32(15) , \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) ,
    \V32(11) , \V32(10) , \V192(27) , \V192(26) , \V192(29) , \V192(28) ,
    \V32(17) , \V32(16) , \V32(19) , \V32(18) , \V32(23) , \V32(22) ,
    \V192(21) , \V32(25) , \V192(20) , \V32(24) , \V192(23) , \V192(22) ,
    \V192(25) , \V32(21) , \V192(24) , \V32(20) , \V192(17) , \V192(16) ,
    \V192(19) , \V192(18) , \V32(27) , \V96(13) , \V32(26) , \V96(12) ,
    \V32(29) , \V96(15) , \V32(28) , \V96(14) , \V192(11) , \V192(10) ,
    \V96(11) , \V192(13) , \V96(10) , \V192(12) , \V192(15) , \V32(31) ,
    \V192(14) , \V32(30) , \V96(17) , \V96(16) , \V96(19) , \V96(18) ,
    \V96(23) , \V96(22) , \V96(25) , \V96(24) , \V96(21) , \V96(20) ,
    \V96(27) , \V96(26) , \V96(29) , \V96(28) , \V192(31) , \V64(0) ,
    \V192(30) , \V96(31) , \V64(1) , \V96(30) , \V64(2) , \V64(3) ,
    \V64(4) , \V64(5) , \V64(6) , \V64(7) , \V64(8) , \V160(3) , \V64(9) ,
    \V160(2) , \V160(5) , \V160(4) , \V160(1) , \V160(0) , \V160(7) ,
    \V160(6) , \V160(9) , \V160(8) , \V160(27) , \V160(26) , \V160(29) ,
    \V160(28) ;
  output \V259(27) , \V259(26) , \V259(29) , \V259(28) , \V259(21) ,
    \V259(20) , \V259(23) , \V259(22) , \V259(25) , \V259(24) , \V259(17) ,
    \V259(16) , \V259(19) , \V259(18) , \V259(11) , \V259(10) , \V259(13) ,
    \V259(12) , \V259(15) , \V259(14) , \V259(3) , \V259(2) , \V259(5) ,
    \V259(4) , \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) ,
    \V259(8) , \V259(31) , \V259(30) , \V227(27) , \V227(26) , \V227(21) ,
    \V227(20) , \V227(23) , \V227(22) , \V227(25) , \V227(24) , \V227(17) ,
    \V227(16) , \V227(19) , \V227(18) , \V227(11) , \V227(10) , \V227(13) ,
    \V227(12) , \V227(15) , \V227(14) , \V266(3) , \V266(2) , \V266(5) ,
    \V266(4) , \V266(1) , \V266(0) , \V266(6) , \V227(3) , \V227(2) ,
    \V227(5) , \V227(4) , \V227(1) , \V227(0) , \V227(7) , \V227(6) ,
    \V227(9) , \V227(8) ;
  wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1055, n1056, n1057, n1058, n1059, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169;
  assign n267 = ~\V199(4)  & \V199(1) ;
  assign n268 = ~\V199(0)  & ~\V192(23) ;
  assign n269 = \V199(1)  & n268;
  assign n270 = \V199(4)  & n269;
  assign n271 = \V160(23)  & \V199(0) ;
  assign n272 = \V199(1)  & n271;
  assign n273 = \V199(4)  & n272;
  assign n274 = ~\V199(0)  & \V192(23) ;
  assign n275 = ~\V199(1)  & n274;
  assign n276 = \V199(4)  & n275;
  assign n277 = \V128(23)  & \V199(0) ;
  assign n278 = ~\V199(1)  & n277;
  assign n279 = \V199(4)  & n278;
  assign n280 = ~n276 & ~n279;
  assign n281 = ~n273 & n280;
  assign n282 = ~n270 & n281;
  assign \V259(27)  = n267 | ~n282;
  assign n284 = ~\V199(0)  & ~\V192(22) ;
  assign n285 = \V199(1)  & n284;
  assign n286 = \V199(4)  & n285;
  assign n287 = \V160(22)  & \V199(0) ;
  assign n288 = \V199(1)  & n287;
  assign n289 = \V199(4)  & n288;
  assign n290 = ~\V199(0)  & \V192(22) ;
  assign n291 = ~\V199(1)  & n290;
  assign n292 = \V199(4)  & n291;
  assign n293 = \V128(22)  & \V199(0) ;
  assign n294 = ~\V199(1)  & n293;
  assign n295 = \V199(4)  & n294;
  assign n296 = ~n292 & ~n295;
  assign n297 = ~n289 & n296;
  assign n298 = ~n286 & n297;
  assign \V259(26)  = n267 | ~n298;
  assign n300 = ~\V199(0)  & ~\V192(25) ;
  assign n301 = \V199(1)  & n300;
  assign n302 = \V199(4)  & n301;
  assign n303 = \V160(25)  & \V199(0) ;
  assign n304 = \V199(1)  & n303;
  assign n305 = \V199(4)  & n304;
  assign n306 = ~\V199(0)  & \V192(25) ;
  assign n307 = ~\V199(1)  & n306;
  assign n308 = \V199(4)  & n307;
  assign n309 = \V128(25)  & \V199(0) ;
  assign n310 = ~\V199(1)  & n309;
  assign n311 = \V199(4)  & n310;
  assign n312 = ~n308 & ~n311;
  assign n313 = ~n305 & n312;
  assign n314 = ~n302 & n313;
  assign \V259(29)  = n267 | ~n314;
  assign n316 = ~\V199(0)  & ~\V192(24) ;
  assign n317 = \V199(1)  & n316;
  assign n318 = \V199(4)  & n317;
  assign n319 = \V160(24)  & \V199(0) ;
  assign n320 = \V199(1)  & n319;
  assign n321 = \V199(4)  & n320;
  assign n322 = ~\V199(0)  & \V192(24) ;
  assign n323 = ~\V199(1)  & n322;
  assign n324 = \V199(4)  & n323;
  assign n325 = \V128(24)  & \V199(0) ;
  assign n326 = ~\V199(1)  & n325;
  assign n327 = \V199(4)  & n326;
  assign n328 = ~n324 & ~n327;
  assign n329 = ~n321 & n328;
  assign n330 = ~n318 & n329;
  assign \V259(28)  = n267 | ~n330;
  assign n332 = ~\V199(0)  & ~\V192(17) ;
  assign n333 = \V199(1)  & n332;
  assign n334 = \V199(4)  & n333;
  assign n335 = \V160(17)  & \V199(0) ;
  assign n336 = \V199(1)  & n335;
  assign n337 = \V199(4)  & n336;
  assign n338 = ~\V199(0)  & \V192(17) ;
  assign n339 = ~\V199(1)  & n338;
  assign n340 = \V199(4)  & n339;
  assign n341 = \V128(17)  & \V199(0) ;
  assign n342 = ~\V199(1)  & n341;
  assign n343 = \V199(4)  & n342;
  assign n344 = ~n340 & ~n343;
  assign n345 = ~n337 & n344;
  assign n346 = ~n334 & n345;
  assign \V259(21)  = n267 | ~n346;
  assign n348 = ~\V199(0)  & ~\V192(16) ;
  assign n349 = \V199(1)  & n348;
  assign n350 = \V199(4)  & n349;
  assign n351 = \V160(16)  & \V199(0) ;
  assign n352 = \V199(1)  & n351;
  assign n353 = \V199(4)  & n352;
  assign n354 = ~\V199(0)  & \V192(16) ;
  assign n355 = ~\V199(1)  & n354;
  assign n356 = \V199(4)  & n355;
  assign n357 = \V128(16)  & \V199(0) ;
  assign n358 = ~\V199(1)  & n357;
  assign n359 = \V199(4)  & n358;
  assign n360 = ~n356 & ~n359;
  assign n361 = ~n353 & n360;
  assign n362 = ~n350 & n361;
  assign \V259(20)  = n267 | ~n362;
  assign n364 = ~\V199(0)  & ~\V192(19) ;
  assign n365 = \V199(1)  & n364;
  assign n366 = \V199(4)  & n365;
  assign n367 = \V160(19)  & \V199(0) ;
  assign n368 = \V199(1)  & n367;
  assign n369 = \V199(4)  & n368;
  assign n370 = ~\V199(0)  & \V192(19) ;
  assign n371 = ~\V199(1)  & n370;
  assign n372 = \V199(4)  & n371;
  assign n373 = \V128(19)  & \V199(0) ;
  assign n374 = ~\V199(1)  & n373;
  assign n375 = \V199(4)  & n374;
  assign n376 = ~n372 & ~n375;
  assign n377 = ~n369 & n376;
  assign n378 = ~n366 & n377;
  assign \V259(23)  = n267 | ~n378;
  assign n380 = ~\V199(0)  & ~\V192(18) ;
  assign n381 = \V199(1)  & n380;
  assign n382 = \V199(4)  & n381;
  assign n383 = \V160(18)  & \V199(0) ;
  assign n384 = \V199(1)  & n383;
  assign n385 = \V199(4)  & n384;
  assign n386 = ~\V199(0)  & \V192(18) ;
  assign n387 = ~\V199(1)  & n386;
  assign n388 = \V199(4)  & n387;
  assign n389 = \V128(18)  & \V199(0) ;
  assign n390 = ~\V199(1)  & n389;
  assign n391 = \V199(4)  & n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = ~n385 & n392;
  assign n394 = ~n382 & n393;
  assign \V259(22)  = n267 | ~n394;
  assign n396 = ~\V199(0)  & ~\V192(21) ;
  assign n397 = \V199(1)  & n396;
  assign n398 = \V199(4)  & n397;
  assign n399 = \V160(21)  & \V199(0) ;
  assign n400 = \V199(1)  & n399;
  assign n401 = \V199(4)  & n400;
  assign n402 = ~\V199(0)  & \V192(21) ;
  assign n403 = ~\V199(1)  & n402;
  assign n404 = \V199(4)  & n403;
  assign n405 = \V128(21)  & \V199(0) ;
  assign n406 = ~\V199(1)  & n405;
  assign n407 = \V199(4)  & n406;
  assign n408 = ~n404 & ~n407;
  assign n409 = ~n401 & n408;
  assign n410 = ~n398 & n409;
  assign \V259(25)  = n267 | ~n410;
  assign n412 = ~\V199(0)  & ~\V192(20) ;
  assign n413 = \V199(1)  & n412;
  assign n414 = \V199(4)  & n413;
  assign n415 = \V160(20)  & \V199(0) ;
  assign n416 = \V199(1)  & n415;
  assign n417 = \V199(4)  & n416;
  assign n418 = ~\V199(0)  & \V192(20) ;
  assign n419 = ~\V199(1)  & n418;
  assign n420 = \V199(4)  & n419;
  assign n421 = \V128(20)  & \V199(0) ;
  assign n422 = ~\V199(1)  & n421;
  assign n423 = \V199(4)  & n422;
  assign n424 = ~n420 & ~n423;
  assign n425 = ~n417 & n424;
  assign n426 = ~n414 & n425;
  assign \V259(24)  = n267 | ~n426;
  assign n428 = ~\V199(0)  & ~\V192(13) ;
  assign n429 = \V199(1)  & n428;
  assign n430 = \V199(4)  & n429;
  assign n431 = \V160(13)  & \V199(0) ;
  assign n432 = \V199(1)  & n431;
  assign n433 = \V199(4)  & n432;
  assign n434 = ~\V199(0)  & \V192(13) ;
  assign n435 = ~\V199(1)  & n434;
  assign n436 = \V199(4)  & n435;
  assign n437 = \V128(13)  & \V199(0) ;
  assign n438 = ~\V199(1)  & n437;
  assign n439 = \V199(4)  & n438;
  assign n440 = ~n436 & ~n439;
  assign n441 = ~n433 & n440;
  assign n442 = ~n430 & n441;
  assign \V259(17)  = n267 | ~n442;
  assign n444 = ~\V199(0)  & ~\V192(12) ;
  assign n445 = \V199(1)  & n444;
  assign n446 = \V199(4)  & n445;
  assign n447 = \V160(12)  & \V199(0) ;
  assign n448 = \V199(1)  & n447;
  assign n449 = \V199(4)  & n448;
  assign n450 = ~\V199(0)  & \V192(12) ;
  assign n451 = ~\V199(1)  & n450;
  assign n452 = \V199(4)  & n451;
  assign n453 = \V128(12)  & \V199(0) ;
  assign n454 = ~\V199(1)  & n453;
  assign n455 = \V199(4)  & n454;
  assign n456 = ~n452 & ~n455;
  assign n457 = ~n449 & n456;
  assign n458 = ~n446 & n457;
  assign \V259(16)  = n267 | ~n458;
  assign n460 = ~\V199(0)  & ~\V192(15) ;
  assign n461 = \V199(1)  & n460;
  assign n462 = \V199(4)  & n461;
  assign n463 = \V160(15)  & \V199(0) ;
  assign n464 = \V199(1)  & n463;
  assign n465 = \V199(4)  & n464;
  assign n466 = ~\V199(0)  & \V192(15) ;
  assign n467 = ~\V199(1)  & n466;
  assign n468 = \V199(4)  & n467;
  assign n469 = \V128(15)  & \V199(0) ;
  assign n470 = ~\V199(1)  & n469;
  assign n471 = \V199(4)  & n470;
  assign n472 = ~n468 & ~n471;
  assign n473 = ~n465 & n472;
  assign n474 = ~n462 & n473;
  assign \V259(19)  = n267 | ~n474;
  assign n476 = ~\V199(0)  & ~\V192(14) ;
  assign n477 = \V199(1)  & n476;
  assign n478 = \V199(4)  & n477;
  assign n479 = \V160(14)  & \V199(0) ;
  assign n480 = \V199(1)  & n479;
  assign n481 = \V199(4)  & n480;
  assign n482 = ~\V199(0)  & \V192(14) ;
  assign n483 = ~\V199(1)  & n482;
  assign n484 = \V199(4)  & n483;
  assign n485 = \V128(14)  & \V199(0) ;
  assign n486 = ~\V199(1)  & n485;
  assign n487 = \V199(4)  & n486;
  assign n488 = ~n484 & ~n487;
  assign n489 = ~n481 & n488;
  assign n490 = ~n478 & n489;
  assign \V259(18)  = n267 | ~n490;
  assign n492 = ~\V192(7)  & ~\V199(0) ;
  assign n493 = \V199(1)  & n492;
  assign n494 = \V199(4)  & n493;
  assign n495 = \V199(0)  & \V160(7) ;
  assign n496 = \V199(1)  & n495;
  assign n497 = \V199(4)  & n496;
  assign n498 = \V192(7)  & ~\V199(0) ;
  assign n499 = ~\V199(1)  & n498;
  assign n500 = \V199(4)  & n499;
  assign n501 = \V128(7)  & \V199(0) ;
  assign n502 = ~\V199(1)  & n501;
  assign n503 = \V199(4)  & n502;
  assign n504 = ~n500 & ~n503;
  assign n505 = ~n497 & n504;
  assign n506 = ~n494 & n505;
  assign \V259(11)  = n267 | ~n506;
  assign n508 = ~\V192(6)  & ~\V199(0) ;
  assign n509 = \V199(1)  & n508;
  assign n510 = \V199(4)  & n509;
  assign n511 = \V199(0)  & \V160(6) ;
  assign n512 = \V199(1)  & n511;
  assign n513 = \V199(4)  & n512;
  assign n514 = \V192(6)  & ~\V199(0) ;
  assign n515 = ~\V199(1)  & n514;
  assign n516 = \V199(4)  & n515;
  assign n517 = \V128(6)  & \V199(0) ;
  assign n518 = ~\V199(1)  & n517;
  assign n519 = \V199(4)  & n518;
  assign n520 = ~n516 & ~n519;
  assign n521 = ~n513 & n520;
  assign n522 = ~n510 & n521;
  assign \V259(10)  = n267 | ~n522;
  assign n524 = ~\V192(9)  & ~\V199(0) ;
  assign n525 = \V199(1)  & n524;
  assign n526 = \V199(4)  & n525;
  assign n527 = \V199(0)  & \V160(9) ;
  assign n528 = \V199(1)  & n527;
  assign n529 = \V199(4)  & n528;
  assign n530 = \V192(9)  & ~\V199(0) ;
  assign n531 = ~\V199(1)  & n530;
  assign n532 = \V199(4)  & n531;
  assign n533 = \V128(9)  & \V199(0) ;
  assign n534 = ~\V199(1)  & n533;
  assign n535 = \V199(4)  & n534;
  assign n536 = ~n532 & ~n535;
  assign n537 = ~n529 & n536;
  assign n538 = ~n526 & n537;
  assign \V259(13)  = n267 | ~n538;
  assign n540 = ~\V192(8)  & ~\V199(0) ;
  assign n541 = \V199(1)  & n540;
  assign n542 = \V199(4)  & n541;
  assign n543 = \V199(0)  & \V160(8) ;
  assign n544 = \V199(1)  & n543;
  assign n545 = \V199(4)  & n544;
  assign n546 = \V192(8)  & ~\V199(0) ;
  assign n547 = ~\V199(1)  & n546;
  assign n548 = \V199(4)  & n547;
  assign n549 = \V128(8)  & \V199(0) ;
  assign n550 = ~\V199(1)  & n549;
  assign n551 = \V199(4)  & n550;
  assign n552 = ~n548 & ~n551;
  assign n553 = ~n545 & n552;
  assign n554 = ~n542 & n553;
  assign \V259(12)  = n267 | ~n554;
  assign n556 = ~\V199(0)  & ~\V192(11) ;
  assign n557 = \V199(1)  & n556;
  assign n558 = \V199(4)  & n557;
  assign n559 = \V160(11)  & \V199(0) ;
  assign n560 = \V199(1)  & n559;
  assign n561 = \V199(4)  & n560;
  assign n562 = ~\V199(0)  & \V192(11) ;
  assign n563 = ~\V199(1)  & n562;
  assign n564 = \V199(4)  & n563;
  assign n565 = \V128(11)  & \V199(0) ;
  assign n566 = ~\V199(1)  & n565;
  assign n567 = \V199(4)  & n566;
  assign n568 = ~n564 & ~n567;
  assign n569 = ~n561 & n568;
  assign n570 = ~n558 & n569;
  assign \V259(15)  = n267 | ~n570;
  assign n572 = ~\V199(0)  & ~\V192(10) ;
  assign n573 = \V199(1)  & n572;
  assign n574 = \V199(4)  & n573;
  assign n575 = \V160(10)  & \V199(0) ;
  assign n576 = \V199(1)  & n575;
  assign n577 = \V199(4)  & n576;
  assign n578 = ~\V199(0)  & \V192(10) ;
  assign n579 = ~\V199(1)  & n578;
  assign n580 = \V199(4)  & n579;
  assign n581 = \V128(10)  & \V199(0) ;
  assign n582 = ~\V199(1)  & n581;
  assign n583 = \V199(4)  & n582;
  assign n584 = ~n580 & ~n583;
  assign n585 = ~n577 & n584;
  assign n586 = ~n574 & n585;
  assign \V259(14)  = n267 | ~n586;
  assign n588 = ~\V199(0)  & ~\V96(31) ;
  assign n589 = \V199(1)  & n588;
  assign n590 = \V199(4)  & n589;
  assign n591 = \V64(31)  & \V199(0) ;
  assign n592 = \V199(1)  & n591;
  assign n593 = \V199(4)  & n592;
  assign n594 = ~\V199(0)  & \V96(31) ;
  assign n595 = ~\V199(1)  & n594;
  assign n596 = \V199(4)  & n595;
  assign n597 = \V199(0)  & \V32(31) ;
  assign n598 = ~\V199(1)  & n597;
  assign n599 = \V199(4)  & n598;
  assign n600 = ~n596 & ~n599;
  assign n601 = ~n593 & n600;
  assign n602 = ~n590 & n601;
  assign \V259(3)  = n267 | ~n602;
  assign n604 = ~\V199(0)  & ~\V96(30) ;
  assign n605 = \V199(1)  & n604;
  assign n606 = \V199(4)  & n605;
  assign n607 = \V64(30)  & \V199(0) ;
  assign n608 = \V199(1)  & n607;
  assign n609 = \V199(4)  & n608;
  assign n610 = ~\V199(0)  & \V96(30) ;
  assign n611 = ~\V199(1)  & n610;
  assign n612 = \V199(4)  & n611;
  assign n613 = \V199(0)  & \V32(30) ;
  assign n614 = ~\V199(1)  & n613;
  assign n615 = \V199(4)  & n614;
  assign n616 = ~n612 & ~n615;
  assign n617 = ~n609 & n616;
  assign n618 = ~n606 & n617;
  assign \V259(2)  = n267 | ~n618;
  assign n620 = ~\V192(1)  & ~\V199(0) ;
  assign n621 = \V199(1)  & n620;
  assign n622 = \V199(4)  & n621;
  assign n623 = \V199(0)  & \V160(1) ;
  assign n624 = \V199(1)  & n623;
  assign n625 = \V199(4)  & n624;
  assign n626 = \V192(1)  & ~\V199(0) ;
  assign n627 = ~\V199(1)  & n626;
  assign n628 = \V199(4)  & n627;
  assign n629 = \V128(1)  & \V199(0) ;
  assign n630 = ~\V199(1)  & n629;
  assign n631 = \V199(4)  & n630;
  assign n632 = ~n628 & ~n631;
  assign n633 = ~n625 & n632;
  assign n634 = ~n622 & n633;
  assign \V259(5)  = n267 | ~n634;
  assign n636 = ~\V192(0)  & ~\V199(0) ;
  assign n637 = \V199(1)  & n636;
  assign n638 = \V199(4)  & n637;
  assign n639 = \V199(0)  & \V160(0) ;
  assign n640 = \V199(1)  & n639;
  assign n641 = \V199(4)  & n640;
  assign n642 = \V192(0)  & ~\V199(0) ;
  assign n643 = ~\V199(1)  & n642;
  assign n644 = \V199(4)  & n643;
  assign n645 = \V128(0)  & \V199(0) ;
  assign n646 = ~\V199(1)  & n645;
  assign n647 = \V199(4)  & n646;
  assign n648 = ~n644 & ~n647;
  assign n649 = ~n641 & n648;
  assign n650 = ~n638 & n649;
  assign \V259(4)  = n267 | ~n650;
  assign n652 = ~\V199(0)  & ~\V96(29) ;
  assign n653 = \V199(1)  & n652;
  assign n654 = \V199(4)  & n653;
  assign n655 = \V64(29)  & \V199(0) ;
  assign n656 = \V199(1)  & n655;
  assign n657 = \V199(4)  & n656;
  assign n658 = ~\V199(0)  & \V96(29) ;
  assign n659 = ~\V199(1)  & n658;
  assign n660 = \V199(4)  & n659;
  assign n661 = \V199(0)  & \V32(29) ;
  assign n662 = ~\V199(1)  & n661;
  assign n663 = \V199(4)  & n662;
  assign n664 = ~n660 & ~n663;
  assign n665 = ~n657 & n664;
  assign n666 = ~n654 & n665;
  assign \V259(1)  = n267 | ~n666;
  assign n668 = ~\V199(0)  & ~\V96(28) ;
  assign n669 = \V199(1)  & n668;
  assign n670 = \V199(4)  & n669;
  assign n671 = \V64(28)  & \V199(0) ;
  assign n672 = \V199(1)  & n671;
  assign n673 = \V199(4)  & n672;
  assign n674 = ~\V199(0)  & \V96(28) ;
  assign n675 = ~\V199(1)  & n674;
  assign n676 = \V199(4)  & n675;
  assign n677 = \V199(0)  & \V32(28) ;
  assign n678 = ~\V199(1)  & n677;
  assign n679 = \V199(4)  & n678;
  assign n680 = ~n676 & ~n679;
  assign n681 = ~n673 & n680;
  assign n682 = ~n670 & n681;
  assign \V259(0)  = n267 | ~n682;
  assign n684 = ~\V192(3)  & ~\V199(0) ;
  assign n685 = \V199(1)  & n684;
  assign n686 = \V199(4)  & n685;
  assign n687 = \V199(0)  & \V160(3) ;
  assign n688 = \V199(1)  & n687;
  assign n689 = \V199(4)  & n688;
  assign n690 = \V192(3)  & ~\V199(0) ;
  assign n691 = ~\V199(1)  & n690;
  assign n692 = \V199(4)  & n691;
  assign n693 = \V128(3)  & \V199(0) ;
  assign n694 = ~\V199(1)  & n693;
  assign n695 = \V199(4)  & n694;
  assign n696 = ~n692 & ~n695;
  assign n697 = ~n689 & n696;
  assign n698 = ~n686 & n697;
  assign \V259(7)  = n267 | ~n698;
  assign n700 = ~\V192(2)  & ~\V199(0) ;
  assign n701 = \V199(1)  & n700;
  assign n702 = \V199(4)  & n701;
  assign n703 = \V199(0)  & \V160(2) ;
  assign n704 = \V199(1)  & n703;
  assign n705 = \V199(4)  & n704;
  assign n706 = \V192(2)  & ~\V199(0) ;
  assign n707 = ~\V199(1)  & n706;
  assign n708 = \V199(4)  & n707;
  assign n709 = \V128(2)  & \V199(0) ;
  assign n710 = ~\V199(1)  & n709;
  assign n711 = \V199(4)  & n710;
  assign n712 = ~n708 & ~n711;
  assign n713 = ~n705 & n712;
  assign n714 = ~n702 & n713;
  assign \V259(6)  = n267 | ~n714;
  assign n716 = ~\V192(5)  & ~\V199(0) ;
  assign n717 = \V199(1)  & n716;
  assign n718 = \V199(4)  & n717;
  assign n719 = \V199(0)  & \V160(5) ;
  assign n720 = \V199(1)  & n719;
  assign n721 = \V199(4)  & n720;
  assign n722 = \V192(5)  & ~\V199(0) ;
  assign n723 = ~\V199(1)  & n722;
  assign n724 = \V199(4)  & n723;
  assign n725 = \V128(5)  & \V199(0) ;
  assign n726 = ~\V199(1)  & n725;
  assign n727 = \V199(4)  & n726;
  assign n728 = ~n724 & ~n727;
  assign n729 = ~n721 & n728;
  assign n730 = ~n718 & n729;
  assign \V259(9)  = n267 | ~n730;
  assign n732 = ~\V192(4)  & ~\V199(0) ;
  assign n733 = \V199(1)  & n732;
  assign n734 = \V199(4)  & n733;
  assign n735 = \V199(0)  & \V160(4) ;
  assign n736 = \V199(1)  & n735;
  assign n737 = \V199(4)  & n736;
  assign n738 = \V192(4)  & ~\V199(0) ;
  assign n739 = ~\V199(1)  & n738;
  assign n740 = \V199(4)  & n739;
  assign n741 = \V128(4)  & \V199(0) ;
  assign n742 = ~\V199(1)  & n741;
  assign n743 = \V199(4)  & n742;
  assign n744 = ~n740 & ~n743;
  assign n745 = ~n737 & n744;
  assign n746 = ~n734 & n745;
  assign \V259(8)  = n267 | ~n746;
  assign n748 = ~\V199(0)  & ~\V192(27) ;
  assign n749 = \V199(1)  & n748;
  assign n750 = \V199(4)  & n749;
  assign n751 = \V199(0)  & \V160(27) ;
  assign n752 = \V199(1)  & n751;
  assign n753 = \V199(4)  & n752;
  assign n754 = ~\V199(0)  & \V192(27) ;
  assign n755 = ~\V199(1)  & n754;
  assign n756 = \V199(4)  & n755;
  assign n757 = \V128(27)  & \V199(0) ;
  assign n758 = ~\V199(1)  & n757;
  assign n759 = \V199(4)  & n758;
  assign n760 = ~n756 & ~n759;
  assign n761 = ~n753 & n760;
  assign n762 = ~n750 & n761;
  assign \V259(31)  = n267 | ~n762;
  assign n764 = ~\V199(0)  & ~\V192(26) ;
  assign n765 = \V199(1)  & n764;
  assign n766 = \V199(4)  & n765;
  assign n767 = \V199(0)  & \V160(26) ;
  assign n768 = \V199(1)  & n767;
  assign n769 = \V199(4)  & n768;
  assign n770 = ~\V199(0)  & \V192(26) ;
  assign n771 = ~\V199(1)  & n770;
  assign n772 = \V199(4)  & n771;
  assign n773 = \V128(26)  & \V199(0) ;
  assign n774 = ~\V199(1)  & n773;
  assign n775 = \V199(4)  & n774;
  assign n776 = ~n772 & ~n775;
  assign n777 = ~n769 & n776;
  assign n778 = ~n766 & n777;
  assign \V259(30)  = n267 | ~n778;
  assign n780 = \V199(1)  & ~\V96(27) ;
  assign n781 = ~\V199(0)  & n780;
  assign n782 = \V64(27)  & \V199(1) ;
  assign n783 = \V199(0)  & n782;
  assign n784 = ~\V199(1)  & \V96(27) ;
  assign n785 = ~\V199(0)  & n784;
  assign n786 = ~\V199(1)  & \V32(27) ;
  assign n787 = \V199(0)  & n786;
  assign n788 = ~n785 & ~n787;
  assign n789 = ~n783 & n788;
  assign \V227(27)  = n781 | ~n789;
  assign n791 = \V199(1)  & ~\V96(26) ;
  assign n792 = ~\V199(0)  & n791;
  assign n793 = \V64(26)  & \V199(1) ;
  assign n794 = \V199(0)  & n793;
  assign n795 = ~\V199(1)  & \V96(26) ;
  assign n796 = ~\V199(0)  & n795;
  assign n797 = ~\V199(1)  & \V32(26) ;
  assign n798 = \V199(0)  & n797;
  assign n799 = ~n796 & ~n798;
  assign n800 = ~n794 & n799;
  assign \V227(26)  = n792 | ~n800;
  assign n802 = \V199(1)  & ~\V96(21) ;
  assign n803 = ~\V199(0)  & n802;
  assign n804 = \V64(21)  & \V199(1) ;
  assign n805 = \V199(0)  & n804;
  assign n806 = ~\V199(1)  & \V96(21) ;
  assign n807 = ~\V199(0)  & n806;
  assign n808 = ~\V199(1)  & \V32(21) ;
  assign n809 = \V199(0)  & n808;
  assign n810 = ~n807 & ~n809;
  assign n811 = ~n805 & n810;
  assign \V227(21)  = n803 | ~n811;
  assign n813 = \V199(1)  & ~\V96(20) ;
  assign n814 = ~\V199(0)  & n813;
  assign n815 = \V64(20)  & \V199(1) ;
  assign n816 = \V199(0)  & n815;
  assign n817 = ~\V199(1)  & \V96(20) ;
  assign n818 = ~\V199(0)  & n817;
  assign n819 = ~\V199(1)  & \V32(20) ;
  assign n820 = \V199(0)  & n819;
  assign n821 = ~n818 & ~n820;
  assign n822 = ~n816 & n821;
  assign \V227(20)  = n814 | ~n822;
  assign n824 = \V199(1)  & ~\V96(23) ;
  assign n825 = ~\V199(0)  & n824;
  assign n826 = \V64(23)  & \V199(1) ;
  assign n827 = \V199(0)  & n826;
  assign n828 = ~\V199(1)  & \V96(23) ;
  assign n829 = ~\V199(0)  & n828;
  assign n830 = ~\V199(1)  & \V32(23) ;
  assign n831 = \V199(0)  & n830;
  assign n832 = ~n829 & ~n831;
  assign n833 = ~n827 & n832;
  assign \V227(23)  = n825 | ~n833;
  assign n835 = \V199(1)  & ~\V96(22) ;
  assign n836 = ~\V199(0)  & n835;
  assign n837 = \V64(22)  & \V199(1) ;
  assign n838 = \V199(0)  & n837;
  assign n839 = ~\V199(1)  & \V96(22) ;
  assign n840 = ~\V199(0)  & n839;
  assign n841 = ~\V199(1)  & \V32(22) ;
  assign n842 = \V199(0)  & n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = ~n838 & n843;
  assign \V227(22)  = n836 | ~n844;
  assign n846 = \V199(1)  & ~\V96(25) ;
  assign n847 = ~\V199(0)  & n846;
  assign n848 = \V64(25)  & \V199(1) ;
  assign n849 = \V199(0)  & n848;
  assign n850 = ~\V199(1)  & \V96(25) ;
  assign n851 = ~\V199(0)  & n850;
  assign n852 = ~\V199(1)  & \V32(25) ;
  assign n853 = \V199(0)  & n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = ~n849 & n854;
  assign \V227(25)  = n847 | ~n855;
  assign n857 = \V199(1)  & ~\V96(24) ;
  assign n858 = ~\V199(0)  & n857;
  assign n859 = \V64(24)  & \V199(1) ;
  assign n860 = \V199(0)  & n859;
  assign n861 = ~\V199(1)  & \V96(24) ;
  assign n862 = ~\V199(0)  & n861;
  assign n863 = ~\V199(1)  & \V32(24) ;
  assign n864 = \V199(0)  & n863;
  assign n865 = ~n862 & ~n864;
  assign n866 = ~n860 & n865;
  assign \V227(24)  = n858 | ~n866;
  assign n868 = \V199(1)  & ~\V96(17) ;
  assign n869 = ~\V199(0)  & n868;
  assign n870 = \V64(17)  & \V199(1) ;
  assign n871 = \V199(0)  & n870;
  assign n872 = ~\V199(1)  & \V96(17) ;
  assign n873 = ~\V199(0)  & n872;
  assign n874 = ~\V199(1)  & \V32(17) ;
  assign n875 = \V199(0)  & n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = ~n871 & n876;
  assign \V227(17)  = n869 | ~n877;
  assign n879 = \V199(1)  & ~\V96(16) ;
  assign n880 = ~\V199(0)  & n879;
  assign n881 = \V64(16)  & \V199(1) ;
  assign n882 = \V199(0)  & n881;
  assign n883 = ~\V199(1)  & \V96(16) ;
  assign n884 = ~\V199(0)  & n883;
  assign n885 = ~\V199(1)  & \V32(16) ;
  assign n886 = \V199(0)  & n885;
  assign n887 = ~n884 & ~n886;
  assign n888 = ~n882 & n887;
  assign \V227(16)  = n880 | ~n888;
  assign n890 = \V199(1)  & ~\V96(19) ;
  assign n891 = ~\V199(0)  & n890;
  assign n892 = \V64(19)  & \V199(1) ;
  assign n893 = \V199(0)  & n892;
  assign n894 = ~\V199(1)  & \V96(19) ;
  assign n895 = ~\V199(0)  & n894;
  assign n896 = ~\V199(1)  & \V32(19) ;
  assign n897 = \V199(0)  & n896;
  assign n898 = ~n895 & ~n897;
  assign n899 = ~n893 & n898;
  assign \V227(19)  = n891 | ~n899;
  assign n901 = \V199(1)  & ~\V96(18) ;
  assign n902 = ~\V199(0)  & n901;
  assign n903 = \V64(18)  & \V199(1) ;
  assign n904 = \V199(0)  & n903;
  assign n905 = ~\V199(1)  & \V96(18) ;
  assign n906 = ~\V199(0)  & n905;
  assign n907 = ~\V199(1)  & \V32(18) ;
  assign n908 = \V199(0)  & n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = ~n904 & n909;
  assign \V227(18)  = n902 | ~n910;
  assign n912 = \V199(1)  & ~\V96(11) ;
  assign n913 = ~\V199(0)  & n912;
  assign n914 = \V64(11)  & \V199(1) ;
  assign n915 = \V199(0)  & n914;
  assign n916 = ~\V199(1)  & \V96(11) ;
  assign n917 = ~\V199(0)  & n916;
  assign n918 = ~\V199(1)  & \V32(11) ;
  assign n919 = \V199(0)  & n918;
  assign n920 = ~n917 & ~n919;
  assign n921 = ~n915 & n920;
  assign \V227(11)  = n913 | ~n921;
  assign n923 = \V199(1)  & ~\V96(10) ;
  assign n924 = ~\V199(0)  & n923;
  assign n925 = \V64(10)  & \V199(1) ;
  assign n926 = \V199(0)  & n925;
  assign n927 = ~\V199(1)  & \V96(10) ;
  assign n928 = ~\V199(0)  & n927;
  assign n929 = ~\V199(1)  & \V32(10) ;
  assign n930 = \V199(0)  & n929;
  assign n931 = ~n928 & ~n930;
  assign n932 = ~n926 & n931;
  assign \V227(10)  = n924 | ~n932;
  assign n934 = \V199(1)  & ~\V96(13) ;
  assign n935 = ~\V199(0)  & n934;
  assign n936 = \V64(13)  & \V199(1) ;
  assign n937 = \V199(0)  & n936;
  assign n938 = ~\V199(1)  & \V96(13) ;
  assign n939 = ~\V199(0)  & n938;
  assign n940 = ~\V199(1)  & \V32(13) ;
  assign n941 = \V199(0)  & n940;
  assign n942 = ~n939 & ~n941;
  assign n943 = ~n937 & n942;
  assign \V227(13)  = n935 | ~n943;
  assign n945 = \V199(1)  & ~\V96(12) ;
  assign n946 = ~\V199(0)  & n945;
  assign n947 = \V64(12)  & \V199(1) ;
  assign n948 = \V199(0)  & n947;
  assign n949 = ~\V199(1)  & \V96(12) ;
  assign n950 = ~\V199(0)  & n949;
  assign n951 = ~\V199(1)  & \V32(12) ;
  assign n952 = \V199(0)  & n951;
  assign n953 = ~n950 & ~n952;
  assign n954 = ~n948 & n953;
  assign \V227(12)  = n946 | ~n954;
  assign n956 = \V199(1)  & ~\V96(15) ;
  assign n957 = ~\V199(0)  & n956;
  assign n958 = \V64(15)  & \V199(1) ;
  assign n959 = \V199(0)  & n958;
  assign n960 = ~\V199(1)  & \V96(15) ;
  assign n961 = ~\V199(0)  & n960;
  assign n962 = ~\V199(1)  & \V32(15) ;
  assign n963 = \V199(0)  & n962;
  assign n964 = ~n961 & ~n963;
  assign n965 = ~n959 & n964;
  assign \V227(15)  = n957 | ~n965;
  assign n967 = \V199(1)  & ~\V96(14) ;
  assign n968 = ~\V199(0)  & n967;
  assign n969 = \V64(14)  & \V199(1) ;
  assign n970 = \V199(0)  & n969;
  assign n971 = ~\V199(1)  & \V96(14) ;
  assign n972 = ~\V199(0)  & n971;
  assign n973 = ~\V199(1)  & \V32(14) ;
  assign n974 = \V199(0)  & n973;
  assign n975 = ~n972 & ~n974;
  assign n976 = ~n970 & n975;
  assign \V227(14)  = n968 | ~n976;
  assign n978 = ~\V199(3)  & \V199(1) ;
  assign n979 = ~\V199(0)  & ~\V192(31) ;
  assign n980 = \V199(1)  & n979;
  assign n981 = \V199(3)  & n980;
  assign n982 = \V199(3)  & \V199(1) ;
  assign n983 = \V199(0)  & n982;
  assign n984 = \V160(31)  & n983;
  assign n985 = ~\V199(0)  & \V192(31) ;
  assign n986 = ~\V199(1)  & n985;
  assign n987 = \V199(3)  & n986;
  assign n988 = \V128(31)  & \V199(0) ;
  assign n989 = ~\V199(1)  & n988;
  assign n990 = \V199(3)  & n989;
  assign n991 = ~n987 & ~n990;
  assign n992 = ~n984 & n991;
  assign n993 = ~n981 & n992;
  assign \V266(3)  = n978 | ~n993;
  assign n995 = ~\V199(0)  & ~\V192(30) ;
  assign n996 = \V199(1)  & n995;
  assign n997 = \V199(3)  & n996;
  assign n998 = \V160(30)  & n983;
  assign n999 = ~\V199(0)  & \V192(30) ;
  assign n1000 = ~\V199(1)  & n999;
  assign n1001 = \V199(3)  & n1000;
  assign n1002 = \V128(30)  & \V199(0) ;
  assign n1003 = ~\V199(1)  & n1002;
  assign n1004 = \V199(3)  & n1003;
  assign n1005 = ~n1001 & ~n1004;
  assign n1006 = ~n998 & n1005;
  assign n1007 = ~n997 & n1006;
  assign \V266(2)  = n978 | ~n1007;
  assign n1009 = ~\V194(1)  & ~\V199(0) ;
  assign n1010 = \V199(1)  & n1009;
  assign n1011 = \V199(3)  & n1010;
  assign n1012 = \V194(1)  & ~\V199(0) ;
  assign n1013 = ~\V199(1)  & n1012;
  assign n1014 = \V199(3)  & n1013;
  assign n1015 = ~n978 & ~n1014;
  assign n1016 = ~n983 & n1015;
  assign \V266(5)  = n1011 | ~n1016;
  assign n1018 = ~\V194(0)  & ~\V199(0) ;
  assign n1019 = \V199(1)  & n1018;
  assign n1020 = \V199(3)  & n1019;
  assign n1021 = \V194(0)  & ~\V199(0) ;
  assign n1022 = ~\V199(1)  & n1021;
  assign n1023 = \V199(3)  & n1022;
  assign n1024 = ~n978 & ~n1023;
  assign n1025 = ~n983 & n1024;
  assign \V266(4)  = n1020 | ~n1025;
  assign n1027 = ~\V199(0)  & ~\V192(29) ;
  assign n1028 = \V199(1)  & n1027;
  assign n1029 = \V199(3)  & n1028;
  assign n1030 = \V160(29)  & n983;
  assign n1031 = ~\V199(0)  & \V192(29) ;
  assign n1032 = ~\V199(1)  & n1031;
  assign n1033 = \V199(3)  & n1032;
  assign n1034 = \V128(29)  & \V199(0) ;
  assign n1035 = ~\V199(1)  & n1034;
  assign n1036 = \V199(3)  & n1035;
  assign n1037 = ~n1033 & ~n1036;
  assign n1038 = ~n1030 & n1037;
  assign n1039 = ~n1029 & n1038;
  assign \V266(1)  = n978 | ~n1039;
  assign n1041 = ~\V199(0)  & ~\V192(28) ;
  assign n1042 = \V199(1)  & n1041;
  assign n1043 = \V199(3)  & n1042;
  assign n1044 = \V160(28)  & n983;
  assign n1045 = ~\V199(0)  & \V192(28) ;
  assign n1046 = ~\V199(1)  & n1045;
  assign n1047 = \V199(3)  & n1046;
  assign n1048 = \V128(28)  & \V199(0) ;
  assign n1049 = ~\V199(1)  & n1048;
  assign n1050 = \V199(3)  & n1049;
  assign n1051 = ~n1047 & ~n1050;
  assign n1052 = ~n1044 & n1051;
  assign n1053 = ~n1043 & n1052;
  assign \V266(0)  = n978 | ~n1053;
  assign n1055 = \V195(0)  & ~\V199(0) ;
  assign n1056 = ~\V199(1)  & n1055;
  assign n1057 = \V199(3)  & n1056;
  assign n1058 = \V199(1)  & n1055;
  assign n1059 = \V199(3)  & n1058;
  assign \V266(6)  = n1057 | n1059;
  assign n1061 = ~\V96(3)  & \V199(1) ;
  assign n1062 = ~\V199(0)  & n1061;
  assign n1063 = \V199(1)  & \V64(3) ;
  assign n1064 = \V199(0)  & n1063;
  assign n1065 = \V96(3)  & ~\V199(1) ;
  assign n1066 = ~\V199(0)  & n1065;
  assign n1067 = ~\V199(1)  & \V32(3) ;
  assign n1068 = \V199(0)  & n1067;
  assign n1069 = ~n1066 & ~n1068;
  assign n1070 = ~n1064 & n1069;
  assign \V227(3)  = n1062 | ~n1070;
  assign n1072 = ~\V96(2)  & \V199(1) ;
  assign n1073 = ~\V199(0)  & n1072;
  assign n1074 = \V199(1)  & \V64(2) ;
  assign n1075 = \V199(0)  & n1074;
  assign n1076 = \V96(2)  & ~\V199(1) ;
  assign n1077 = ~\V199(0)  & n1076;
  assign n1078 = ~\V199(1)  & \V32(2) ;
  assign n1079 = \V199(0)  & n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = ~n1075 & n1080;
  assign \V227(2)  = n1073 | ~n1081;
  assign n1083 = ~\V96(5)  & \V199(1) ;
  assign n1084 = ~\V199(0)  & n1083;
  assign n1085 = \V199(1)  & \V64(5) ;
  assign n1086 = \V199(0)  & n1085;
  assign n1087 = \V96(5)  & ~\V199(1) ;
  assign n1088 = ~\V199(0)  & n1087;
  assign n1089 = ~\V199(1)  & \V32(5) ;
  assign n1090 = \V199(0)  & n1089;
  assign n1091 = ~n1088 & ~n1090;
  assign n1092 = ~n1086 & n1091;
  assign \V227(5)  = n1084 | ~n1092;
  assign n1094 = ~\V96(4)  & \V199(1) ;
  assign n1095 = ~\V199(0)  & n1094;
  assign n1096 = \V199(1)  & \V64(4) ;
  assign n1097 = \V199(0)  & n1096;
  assign n1098 = \V96(4)  & ~\V199(1) ;
  assign n1099 = ~\V199(0)  & n1098;
  assign n1100 = ~\V199(1)  & \V32(4) ;
  assign n1101 = \V199(0)  & n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~n1097 & n1102;
  assign \V227(4)  = n1095 | ~n1103;
  assign n1105 = ~\V96(1)  & \V199(1) ;
  assign n1106 = ~\V199(0)  & n1105;
  assign n1107 = \V199(1)  & \V64(1) ;
  assign n1108 = \V199(0)  & n1107;
  assign n1109 = \V96(1)  & ~\V199(1) ;
  assign n1110 = ~\V199(0)  & n1109;
  assign n1111 = ~\V199(1)  & \V32(1) ;
  assign n1112 = \V199(0)  & n1111;
  assign n1113 = ~n1110 & ~n1112;
  assign n1114 = ~n1108 & n1113;
  assign \V227(1)  = n1106 | ~n1114;
  assign n1116 = ~\V96(0)  & \V199(1) ;
  assign n1117 = ~\V199(0)  & n1116;
  assign n1118 = \V199(1)  & \V64(0) ;
  assign n1119 = \V199(0)  & n1118;
  assign n1120 = \V96(0)  & ~\V199(1) ;
  assign n1121 = ~\V199(0)  & n1120;
  assign n1122 = ~\V199(1)  & \V32(0) ;
  assign n1123 = \V199(0)  & n1122;
  assign n1124 = ~n1121 & ~n1123;
  assign n1125 = ~n1119 & n1124;
  assign \V227(0)  = n1117 | ~n1125;
  assign n1127 = ~\V96(7)  & \V199(1) ;
  assign n1128 = ~\V199(0)  & n1127;
  assign n1129 = \V199(1)  & \V64(7) ;
  assign n1130 = \V199(0)  & n1129;
  assign n1131 = \V96(7)  & ~\V199(1) ;
  assign n1132 = ~\V199(0)  & n1131;
  assign n1133 = ~\V199(1)  & \V32(7) ;
  assign n1134 = \V199(0)  & n1133;
  assign n1135 = ~n1132 & ~n1134;
  assign n1136 = ~n1130 & n1135;
  assign \V227(7)  = n1128 | ~n1136;
  assign n1138 = ~\V96(6)  & \V199(1) ;
  assign n1139 = ~\V199(0)  & n1138;
  assign n1140 = \V199(1)  & \V64(6) ;
  assign n1141 = \V199(0)  & n1140;
  assign n1142 = \V96(6)  & ~\V199(1) ;
  assign n1143 = ~\V199(0)  & n1142;
  assign n1144 = ~\V199(1)  & \V32(6) ;
  assign n1145 = \V199(0)  & n1144;
  assign n1146 = ~n1143 & ~n1145;
  assign n1147 = ~n1141 & n1146;
  assign \V227(6)  = n1139 | ~n1147;
  assign n1149 = ~\V96(9)  & \V199(1) ;
  assign n1150 = ~\V199(0)  & n1149;
  assign n1151 = \V199(1)  & \V64(9) ;
  assign n1152 = \V199(0)  & n1151;
  assign n1153 = \V96(9)  & ~\V199(1) ;
  assign n1154 = ~\V199(0)  & n1153;
  assign n1155 = ~\V199(1)  & \V32(9) ;
  assign n1156 = \V199(0)  & n1155;
  assign n1157 = ~n1154 & ~n1156;
  assign n1158 = ~n1152 & n1157;
  assign \V227(9)  = n1150 | ~n1158;
  assign n1160 = ~\V96(8)  & \V199(1) ;
  assign n1161 = ~\V199(0)  & n1160;
  assign n1162 = \V199(1)  & \V64(8) ;
  assign n1163 = \V199(0)  & n1162;
  assign n1164 = \V96(8)  & ~\V199(1) ;
  assign n1165 = ~\V199(0)  & n1164;
  assign n1166 = ~\V199(1)  & \V32(8) ;
  assign n1167 = \V199(0)  & n1166;
  assign n1168 = ~n1165 & ~n1167;
  assign n1169 = ~n1163 & n1168;
  assign \V227(8)  = n1161 | ~n1169;
endmodule


