// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:01 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_,
    i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_,
    i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_,
    o_0_, o_1_, o_2_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_,
    i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_,
    i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_;
  output o_0_, o_1_, o_2_;
  wire n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306;
  assign n43 = i_13_ & i_14_;
  assign n44 = ~i_16_ & ~i_23_;
  assign n45 = ~n43 & n44;
  assign n46 = ~i_4_ & ~i_5_;
  assign n47 = ~i_2_ & n46;
  assign n48 = ~i_6_ & ~i_12_;
  assign n49 = n47 & n48;
  assign n50 = n45 & n49;
  assign n51 = ~i_8_ & ~i_31_;
  assign n52 = n50 & n51;
  assign n53 = ~i_31_ & ~i_32_;
  assign n54 = ~i_6_ & n46;
  assign n55 = ~i_1_ & n54;
  assign n56 = ~i_2_ & n55;
  assign n57 = ~i_23_ & n56;
  assign n58 = ~i_16_ & ~i_17_;
  assign n59 = ~i_13_ & n58;
  assign n60 = n57 & n59;
  assign n61 = ~i_14_ & ~i_16_;
  assign n62 = ~i_17_ & n61;
  assign n63 = n57 & n62;
  assign n64 = ~n60 & ~n63;
  assign n65 = n53 & ~n64;
  assign n66 = ~i_11_ & ~i_19_;
  assign n67 = i_3_ & ~i_18_;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~i_9_ & ~n68;
  assign n70 = n54 & n69;
  assign n71 = ~i_23_ & n59;
  assign n72 = ~i_2_ & ~i_8_;
  assign n73 = n71 & n72;
  assign n74 = n70 & n73;
  assign n75 = ~n65 & ~n74;
  assign n76 = ~n52 & n75;
  assign n77 = ~i_24_ & ~i_28_;
  assign n78 = ~i_29_ & n77;
  assign n79 = ~i_27_ & n78;
  assign n80 = ~n76 & n79;
  assign n81 = ~i_6_ & ~i_9_;
  assign n82 = ~i_10_ & n81;
  assign n83 = n59 & n82;
  assign n84 = n47 & n83;
  assign n85 = n47 & n81;
  assign n86 = i_13_ & n85;
  assign n87 = n62 & n86;
  assign n88 = ~n84 & ~n87;
  assign n89 = ~i_28_ & ~i_29_;
  assign n90 = ~i_27_ & n89;
  assign n91 = ~i_23_ & ~i_24_;
  assign n92 = n90 & n91;
  assign n93 = ~i_32_ & n92;
  assign n94 = ~n88 & n93;
  assign n95 = i_10_ & ~i_13_;
  assign n96 = ~i_13_ & ~i_16_;
  assign n97 = ~n61 & ~n96;
  assign n98 = ~n95 & ~n97;
  assign n99 = ~i_23_ & ~i_27_;
  assign n100 = ~i_17_ & n99;
  assign n101 = n78 & n100;
  assign n102 = ~i_8_ & n81;
  assign n103 = n47 & n102;
  assign n104 = n101 & n103;
  assign n105 = n98 & n104;
  assign n106 = ~i_31_ & n56;
  assign n107 = ~i_17_ & ~n97;
  assign n108 = ~i_8_ & n107;
  assign n109 = n106 & n108;
  assign n110 = n92 & n109;
  assign n111 = ~n105 & ~n110;
  assign n112 = ~n94 & n111;
  assign n113 = ~n80 & n112;
  assign n114 = ~i_35_ & ~n113;
  assign n115 = ~i_7_ & n56;
  assign n116 = ~n97 & n115;
  assign n117 = ~i_8_ & n116;
  assign n118 = ~i_7_ & n85;
  assign n119 = ~i_32_ & n118;
  assign n120 = n98 & n119;
  assign n121 = ~n117 & ~n120;
  assign n122 = n101 & ~n121;
  assign n123 = ~i_7_ & ~i_32_;
  assign n124 = n107 & n123;
  assign n125 = n56 & n124;
  assign n126 = n92 & n125;
  assign n127 = ~n122 & ~n126;
  assign n128 = ~n114 & n127;
  assign n129 = i_34_ & ~n128;
  assign n130 = ~i_24_ & ~i_26_;
  assign n131 = n99 & n130;
  assign n132 = ~i_17_ & ~i_21_;
  assign n133 = n131 & n132;
  assign n134 = ~i_7_ & ~i_8_;
  assign n135 = n54 & n134;
  assign n136 = ~i_9_ & n135;
  assign n137 = ~i_28_ & i_29_;
  assign n138 = n98 & n137;
  assign n139 = n136 & n138;
  assign n140 = ~i_8_ & ~i_28_;
  assign n141 = n116 & n140;
  assign n142 = ~n139 & ~n141;
  assign n143 = n133 & ~n142;
  assign n144 = ~i_28_ & ~i_30_;
  assign n145 = n53 & n144;
  assign n146 = ~i_34_ & i_35_;
  assign n147 = ~i_29_ & n146;
  assign n148 = n145 & n147;
  assign n149 = ~i_14_ & n44;
  assign n150 = ~i_24_ & i_34_;
  assign n151 = ~n146 & ~n150;
  assign n152 = n90 & ~n151;
  assign n153 = ~i_32_ & n152;
  assign n154 = n149 & n153;
  assign n155 = n49 & n154;
  assign n156 = ~n148 & ~n155;
  assign n157 = ~i_27_ & ~i_28_;
  assign n158 = ~i_26_ & n157;
  assign n159 = ~i_21_ & n91;
  assign n160 = n158 & n159;
  assign n161 = n107 & n160;
  assign n162 = ~i_2_ & ~i_30_;
  assign n163 = n161 & n162;
  assign n164 = ~i_30_ & ~i_31_;
  assign n165 = ~i_28_ & n164;
  assign n166 = ~i_29_ & n91;
  assign n167 = i_34_ & n166;
  assign n168 = n165 & n167;
  assign n169 = ~n163 & ~n168;
  assign n170 = ~i_32_ & ~n169;
  assign n171 = n156 & ~n170;
  assign n172 = ~i_7_ & ~n171;
  assign n173 = ~n143 & ~n172;
  assign n174 = ~i_28_ & n147;
  assign n175 = n100 & n174;
  assign n176 = ~n121 & n175;
  assign n177 = ~i_27_ & n130;
  assign n178 = n89 & n123;
  assign n179 = n50 & n178;
  assign n180 = ~i_32_ & n144;
  assign n181 = ~i_32_ & n137;
  assign n182 = n54 & n181;
  assign n183 = ~n180 & ~n182;
  assign n184 = ~i_12_ & ~n43;
  assign n185 = ~i_7_ & n184;
  assign n186 = ~i_21_ & n44;
  assign n187 = n185 & n186;
  assign n188 = ~n183 & n187;
  assign n189 = ~n179 & ~n188;
  assign n190 = n177 & ~n189;
  assign n191 = n147 & n157;
  assign n192 = ~i_23_ & n191;
  assign n193 = ~i_28_ & n130;
  assign n194 = n99 & n193;
  assign n195 = i_21_ & i_29_;
  assign n196 = n194 & ~n195;
  assign n197 = ~n192 & ~n196;
  assign n198 = n125 & ~n197;
  assign n199 = ~n190 & ~n198;
  assign n200 = n96 & n134;
  assign n201 = n132 & n200;
  assign n202 = i_29_ & n54;
  assign n203 = n69 & n194;
  assign n204 = n202 & n203;
  assign n205 = n201 & n204;
  assign n206 = ~i_30_ & ~i_32_;
  assign n207 = n185 & n206;
  assign n208 = n44 & n191;
  assign n209 = n207 & n208;
  assign n210 = n49 & n134;
  assign n211 = ~i_26_ & n91;
  assign n212 = n90 & n211;
  assign n213 = ~n97 & n212;
  assign n214 = n210 & n213;
  assign n215 = ~n209 & ~n214;
  assign n216 = ~n205 & n215;
  assign n217 = n199 & n216;
  assign n218 = ~n176 & n217;
  assign n219 = n173 & n218;
  assign n220 = ~i_8_ & n118;
  assign n221 = ~i_10_ & n220;
  assign n222 = n71 & n221;
  assign n223 = ~i_2_ & n70;
  assign n224 = ~i_17_ & n223;
  assign n225 = ~n49 & ~n224;
  assign n226 = n200 & ~n225;
  assign n227 = n61 & n210;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~i_23_ & ~n228;
  assign n230 = ~i_13_ & n44;
  assign n231 = ~i_7_ & ~n225;
  assign n232 = n230 & n231;
  assign n233 = ~i_32_ & n232;
  assign n234 = ~i_23_ & n134;
  assign n235 = n87 & n234;
  assign n236 = ~n233 & ~n235;
  assign n237 = ~n229 & n236;
  assign n238 = ~n222 & n237;
  assign n239 = n152 & ~n238;
  assign n240 = n219 & ~n239;
  assign n241 = ~n129 & n240;
  assign n242 = i_36_ & ~n241;
  assign n243 = i_31_ & n157;
  assign n244 = i_21_ & ~i_23_;
  assign n245 = ~n151 & n244;
  assign n246 = n243 & n245;
  assign n247 = i_7_ & ~i_9_;
  assign n248 = ~i_12_ & n247;
  assign n249 = n246 & n248;
  assign n250 = ~i_32_ & i_34_;
  assign n251 = n101 & n250;
  assign n252 = ~i_32_ & n175;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~i_30_ & ~n253;
  assign n255 = ~i_29_ & n206;
  assign n256 = n193 & n255;
  assign n257 = n100 & n256;
  assign n258 = ~n254 & ~n257;
  assign n259 = ~i_7_ & ~n258;
  assign n260 = i_30_ & ~n202;
  assign n261 = ~i_8_ & ~i_12_;
  assign n262 = ~i_7_ & n261;
  assign n263 = ~n260 & n262;
  assign n264 = n160 & n263;
  assign n265 = ~n259 & ~n264;
  assign n266 = i_36_ & ~n265;
  assign n267 = i_0_ & n137;
  assign n268 = ~i_35_ & i_36_;
  assign n269 = ~i_32_ & n268;
  assign n270 = ~i_2_ & n269;
  assign n271 = n165 & n270;
  assign n272 = ~n267 & ~n271;
  assign n273 = n133 & ~n272;
  assign n274 = ~n266 & ~n273;
  assign n275 = ~n249 & n274;
  assign n276 = ~n97 & ~n275;
  assign n277 = n131 & n137;
  assign n278 = ~i_8_ & ~i_35_;
  assign n279 = ~n123 & ~n278;
  assign n280 = i_36_ & n54;
  assign n281 = ~n279 & n280;
  assign n282 = ~i_2_ & ~n281;
  assign n283 = n59 & n69;
  assign n284 = ~n282 & n283;
  assign n285 = n277 & n284;
  assign n286 = n164 & n181;
  assign n287 = ~i_23_ & n150;
  assign n288 = ~i_34_ & n130;
  assign n289 = ~n146 & ~n288;
  assign n290 = ~n287 & n289;
  assign n291 = n286 & ~n290;
  assign n292 = i_20_ & n291;
  assign n293 = ~n285 & ~n292;
  assign n294 = ~i_21_ & ~n293;
  assign n295 = i_7_ & i_10_;
  assign n296 = i_12_ & i_17_;
  assign n297 = n96 & ~n296;
  assign n298 = i_31_ & n297;
  assign n299 = ~n68 & n298;
  assign n300 = n295 & n299;
  assign n301 = n61 & ~n296;
  assign n302 = i_25_ & i_33_;
  assign n303 = n301 & n302;
  assign n304 = n245 & n303;
  assign n305 = ~n300 & ~n304;
  assign n306 = ~n167 & ~n211;
  assign n307 = ~n245 & n306;
  assign n308 = n157 & ~n307;
  assign n309 = ~n305 & n308;
  assign n310 = ~n43 & ~n296;
  assign n311 = ~i_16_ & n310;
  assign n312 = n277 & n311;
  assign n313 = ~i_21_ & ~i_22_;
  assign n314 = i_20_ & n313;
  assign n315 = n312 & n314;
  assign n316 = n45 & ~n296;
  assign n317 = ~i_27_ & n316;
  assign n318 = n137 & n146;
  assign n319 = i_22_ & n318;
  assign n320 = n317 & n319;
  assign n321 = ~n315 & ~n320;
  assign n322 = i_14_ & i_33_;
  assign n323 = ~n302 & ~n322;
  assign n324 = ~i_21_ & i_29_;
  assign n325 = n145 & ~n289;
  assign n326 = ~n324 & n325;
  assign n327 = ~n323 & n326;
  assign n328 = n321 & ~n327;
  assign n329 = ~n309 & n328;
  assign n330 = ~n294 & n329;
  assign n331 = n243 & n301;
  assign n332 = i_13_ & n331;
  assign n333 = n295 & n332;
  assign n334 = n244 & n333;
  assign n335 = i_20_ & ~i_23_;
  assign n336 = n157 & n335;
  assign n337 = n324 & n336;
  assign n338 = n311 & n337;
  assign n339 = ~n334 & ~n338;
  assign n340 = ~i_31_ & n206;
  assign n341 = ~i_28_ & n244;
  assign n342 = n340 & n341;
  assign n343 = ~n323 & n342;
  assign n344 = n339 & ~n343;
  assign n345 = n150 & ~n344;
  assign n346 = n297 & n322;
  assign n347 = ~n300 & ~n346;
  assign n348 = ~n303 & n347;
  assign n349 = n192 & ~n348;
  assign n350 = ~n130 & ~n147;
  assign n351 = ~i_23_ & ~n350;
  assign n352 = ~n167 & ~n351;
  assign n353 = n333 & ~n352;
  assign n354 = ~n349 & ~n353;
  assign n355 = ~n345 & n354;
  assign n356 = i_22_ & n286;
  assign n357 = n339 & ~n356;
  assign n358 = n146 & ~n357;
  assign n359 = ~n307 & n346;
  assign n360 = n303 & ~n306;
  assign n361 = ~i_12_ & ~n97;
  assign n362 = ~i_30_ & n123;
  assign n363 = ~i_29_ & i_36_;
  assign n364 = n91 & n363;
  assign n365 = n362 & n364;
  assign n366 = n361 & n365;
  assign n367 = i_34_ & n366;
  assign n368 = ~n360 & ~n367;
  assign n369 = ~n359 & n368;
  assign n370 = n157 & ~n369;
  assign n371 = n184 & n186;
  assign n372 = n267 & n371;
  assign n373 = n177 & n372;
  assign n374 = ~n370 & ~n373;
  assign n375 = ~n358 & n374;
  assign n376 = n355 & n375;
  assign n377 = n145 & n166;
  assign n378 = n322 & n377;
  assign n379 = n302 & n377;
  assign n380 = ~n62 & ~n361;
  assign n381 = i_22_ & n91;
  assign n382 = ~i_27_ & n137;
  assign n383 = n381 & n382;
  assign n384 = ~n380 & n383;
  assign n385 = ~n379 & ~n384;
  assign n386 = ~i_8_ & ~i_24_;
  assign n387 = ~n296 & n386;
  assign n388 = n164 & n387;
  assign n389 = n45 & n388;
  assign n390 = n268 & n389;
  assign n391 = n90 & n390;
  assign n392 = n385 & ~n391;
  assign n393 = ~n378 & n392;
  assign n394 = i_34_ & ~n393;
  assign n395 = n90 & n150;
  assign n396 = n157 & ~n350;
  assign n397 = ~n395 & ~n396;
  assign n398 = i_31_ & ~n397;
  assign n399 = ~i_23_ & n398;
  assign n400 = ~n246 & ~n399;
  assign n401 = n107 & n247;
  assign n402 = ~n400 & n401;
  assign n403 = ~n394 & ~n402;
  assign n404 = n248 & n398;
  assign n405 = ~i_30_ & n157;
  assign n406 = ~n130 & n151;
  assign n407 = n363 & ~n406;
  assign n408 = n405 & n407;
  assign n409 = n262 & n408;
  assign n410 = ~n404 & ~n409;
  assign n411 = n45 & ~n410;
  assign n412 = n59 & n382;
  assign n413 = ~n286 & ~n412;
  assign n414 = i_34_ & ~n413;
  assign n415 = ~n62 & ~n297;
  assign n416 = n158 & ~n415;
  assign n417 = i_29_ & n416;
  assign n418 = ~n414 & ~n417;
  assign n419 = n381 & ~n418;
  assign n420 = n288 & n356;
  assign n421 = ~i_12_ & i_29_;
  assign n422 = ~i_20_ & ~i_21_;
  assign n423 = n421 & n422;
  assign n424 = i_2_ & ~n97;
  assign n425 = n423 & n424;
  assign n426 = n194 & n425;
  assign n427 = ~n420 & ~n426;
  assign n428 = ~n419 & n427;
  assign n429 = n107 & n234;
  assign n430 = n408 & n429;
  assign n431 = n428 & ~n430;
  assign n432 = ~n411 & n431;
  assign n433 = n403 & n432;
  assign n434 = n376 & n433;
  assign n435 = n330 & n434;
  assign n436 = ~i_17_ & n91;
  assign n437 = ~i_32_ & n96;
  assign n438 = n223 & n437;
  assign n439 = ~i_35_ & n438;
  assign n440 = ~n117 & ~n439;
  assign n441 = n436 & ~n440;
  assign n442 = n50 & n53;
  assign n443 = ~i_24_ & n442;
  assign n444 = n103 & n436;
  assign n445 = n98 & n444;
  assign n446 = ~n389 & ~n445;
  assign n447 = ~n443 & n446;
  assign n448 = ~i_35_ & ~n447;
  assign n449 = ~n441 & ~n448;
  assign n450 = n363 & ~n449;
  assign n451 = ~i_31_ & ~n260;
  assign n452 = n361 & n451;
  assign n453 = n202 & n283;
  assign n454 = ~n452 & ~n453;
  assign n455 = n159 & ~n454;
  assign n456 = n269 & n455;
  assign n457 = ~i_30_ & n134;
  assign n458 = ~i_2_ & n457;
  assign n459 = i_36_ & n458;
  assign n460 = i_29_ & ~n95;
  assign n461 = ~i_9_ & n460;
  assign n462 = ~n282 & n461;
  assign n463 = ~n459 & ~n462;
  assign n464 = n107 & n159;
  assign n465 = ~n463 & n464;
  assign n466 = n61 & n381;
  assign n467 = n421 & n466;
  assign n468 = ~n366 & ~n467;
  assign n469 = ~n465 & n468;
  assign n470 = ~n456 & n469;
  assign n471 = ~n450 & n470;
  assign n472 = n158 & ~n471;
  assign n473 = n435 & ~n472;
  assign n474 = ~n276 & n473;
  assign n475 = ~i_29_ & n288;
  assign n476 = n165 & n475;
  assign n477 = n54 & n461;
  assign n478 = ~n106 & ~n477;
  assign n479 = n161 & ~n478;
  assign n480 = ~n88 & n212;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n476 & n481;
  assign n483 = ~i_32_ & ~n482;
  assign n484 = n109 & n196;
  assign n485 = n395 & n442;
  assign n486 = ~n484 & ~n485;
  assign n487 = n96 & n223;
  assign n488 = n251 & n487;
  assign n489 = n145 & n167;
  assign n490 = n51 & n163;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~n488 & n491;
  assign n493 = n486 & n492;
  assign n494 = ~n76 & n89;
  assign n495 = n140 & n371;
  assign n496 = n451 & n495;
  assign n497 = ~n494 & ~n496;
  assign n498 = n177 & ~n497;
  assign n499 = n493 & ~n498;
  assign n500 = ~n483 & n499;
  assign n501 = n268 & ~n500;
  assign n502 = n474 & ~n501;
  assign o_0_ = n242 | ~n502;
  assign n504 = ~i_31_ & n89;
  assign n505 = n362 & n504;
  assign n506 = i_37_ & n146;
  assign n507 = n505 & n506;
  assign n508 = ~i_35_ & i_37_;
  assign n509 = n489 & n508;
  assign n510 = i_37_ & n123;
  assign n511 = n168 & n510;
  assign n512 = ~n509 & ~n511;
  assign n513 = ~i_23_ & n152;
  assign n514 = n134 & n223;
  assign n515 = ~n221 & ~n514;
  assign n516 = ~n457 & n515;
  assign n517 = n513 & ~n516;
  assign n518 = n81 & ~n95;
  assign n519 = ~i_20_ & n211;
  assign n520 = n382 & n519;
  assign n521 = ~i_0_ & ~i_4_;
  assign n522 = ~i_5_ & n521;
  assign n523 = n134 & n522;
  assign n524 = n520 & n523;
  assign n525 = n518 & n524;
  assign n526 = ~n517 & ~n525;
  assign n527 = i_37_ & n58;
  assign n528 = ~n526 & n527;
  assign n529 = n512 & ~n528;
  assign n530 = ~n507 & n529;
  assign n531 = ~i_14_ & ~n530;
  assign n532 = n148 & n302;
  assign n533 = ~i_10_ & n96;
  assign n534 = ~i_33_ & n533;
  assign n535 = ~i_29_ & n158;
  assign n536 = n508 & n535;
  assign n537 = n444 & n536;
  assign n538 = n534 & n537;
  assign n539 = ~i_8_ & n211;
  assign n540 = ~i_0_ & ~i_20_;
  assign n541 = ~n322 & n508;
  assign n542 = n540 & n541;
  assign n543 = n311 & n405;
  assign n544 = n542 & n543;
  assign n545 = n539 & n544;
  assign n546 = ~n538 & ~n545;
  assign n547 = n428 & n546;
  assign n548 = ~n532 & n547;
  assign n549 = ~n531 & n548;
  assign n550 = ~i_33_ & n230;
  assign n551 = ~i_8_ & ~n225;
  assign n552 = n550 & n551;
  assign n553 = ~i_8_ & n63;
  assign n554 = ~n552 & ~n553;
  assign n555 = n395 & n508;
  assign n556 = ~n554 & n555;
  assign n557 = n108 & n541;
  assign n558 = ~i_1_ & n521;
  assign n559 = ~i_32_ & ~i_33_;
  assign n560 = i_37_ & n559;
  assign n561 = n59 & n560;
  assign n562 = n558 & n561;
  assign n563 = ~i_7_ & n562;
  assign n564 = ~n557 & ~n563;
  assign n565 = ~i_0_ & n55;
  assign n566 = ~i_5_ & ~i_6_;
  assign n567 = n67 & n521;
  assign n568 = ~i_9_ & n567;
  assign n569 = n566 & n568;
  assign n570 = ~n565 & ~n569;
  assign n571 = ~n564 & ~n570;
  assign n572 = ~i_6_ & ~n322;
  assign n573 = i_37_ & n523;
  assign n574 = n69 & n107;
  assign n575 = ~n361 & ~n574;
  assign n576 = n573 & ~n575;
  assign n577 = n572 & n576;
  assign n578 = ~n571 & ~n577;
  assign n579 = n520 & ~n578;
  assign n580 = ~i_33_ & n89;
  assign n581 = ~i_23_ & n506;
  assign n582 = ~i_27_ & n581;
  assign n583 = n580 & n582;
  assign n584 = n226 & n583;
  assign n585 = ~n579 & ~n584;
  assign n586 = n56 & n557;
  assign n587 = ~i_35_ & n84;
  assign n588 = ~i_30_ & n298;
  assign n589 = ~n587 & ~n588;
  assign n590 = n560 & ~n589;
  assign n591 = ~n586 & ~n590;
  assign n592 = n212 & ~n591;
  assign n593 = n508 & n522;
  assign n594 = ~n97 & ~n322;
  assign n595 = ~i_20_ & n48;
  assign n596 = ~i_8_ & n595;
  assign n597 = n277 & n596;
  assign n598 = ~i_17_ & n520;
  assign n599 = n66 & n102;
  assign n600 = n598 & n599;
  assign n601 = ~n597 & ~n600;
  assign n602 = n594 & ~n601;
  assign n603 = n593 & n602;
  assign n604 = ~n592 & ~n603;
  assign n605 = n585 & n604;
  assign n606 = ~n556 & n605;
  assign n607 = n117 & ~n322;
  assign n608 = n61 & ~n95;
  assign n609 = n119 & n608;
  assign n610 = ~n607 & ~n609;
  assign n611 = n175 & ~n610;
  assign n612 = i_37_ & n611;
  assign n613 = i_37_ & n152;
  assign n614 = n235 & n613;
  assign n615 = n150 & n244;
  assign n616 = n286 & n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = n192 & n561;
  assign n619 = n115 & n618;
  assign n620 = ~i_20_ & ~n475;
  assign n621 = n325 & ~n620;
  assign n622 = n302 & n621;
  assign n623 = ~n619 & ~n622;
  assign n624 = ~i_33_ & n506;
  assign n625 = n505 & n624;
  assign n626 = n623 & ~n625;
  assign n627 = n617 & n626;
  assign n628 = i_34_ & ~n385;
  assign n629 = n627 & ~n628;
  assign n630 = ~n612 & n629;
  assign n631 = ~n313 & n318;
  assign n632 = n99 & n631;
  assign n633 = i_7_ & i_31_;
  assign n634 = ~n302 & ~n633;
  assign n635 = ~i_20_ & ~n147;
  assign n636 = ~i_23_ & ~n635;
  assign n637 = ~n151 & n636;
  assign n638 = n306 & ~n637;
  assign n639 = n157 & ~n638;
  assign n640 = ~n634 & n639;
  assign n641 = n382 & n615;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n632 & n642;
  assign n644 = n311 & ~n643;
  assign n645 = n630 & ~n644;
  assign n646 = n606 & n645;
  assign n647 = i_34_ & n508;
  assign n648 = n104 & n534;
  assign n649 = n149 & n551;
  assign n650 = ~i_32_ & n63;
  assign n651 = ~n649 & ~n650;
  assign n652 = n79 & ~n651;
  assign n653 = n85 & ~n95;
  assign n654 = n62 & n653;
  assign n655 = ~i_33_ & n84;
  assign n656 = ~n654 & ~n655;
  assign n657 = n93 & ~n656;
  assign n658 = ~n652 & ~n657;
  assign n659 = ~n648 & n658;
  assign n660 = n647 & ~n659;
  assign n661 = n646 & ~n660;
  assign n662 = n549 & n661;
  assign n663 = ~i_17_ & ~i_23_;
  assign n664 = ~i_20_ & n663;
  assign n665 = ~i_7_ & n566;
  assign n666 = i_37_ & n558;
  assign n667 = n665 & n666;
  assign n668 = ~i_8_ & n594;
  assign n669 = n667 & n668;
  assign n670 = ~n534 & ~n608;
  assign n671 = n102 & ~n670;
  assign n672 = n593 & n671;
  assign n673 = ~n424 & ~n672;
  assign n674 = ~n669 & n673;
  assign n675 = n664 & ~n674;
  assign n676 = n137 & n675;
  assign n677 = ~i_23_ & n54;
  assign n678 = n542 & n677;
  assign n679 = n574 & n678;
  assign n680 = ~i_7_ & n81;
  assign n681 = i_37_ & n680;
  assign n682 = n664 & n681;
  assign n683 = ~n670 & n682;
  assign n684 = n541 & n595;
  assign n685 = n45 & n684;
  assign n686 = ~n683 & ~n685;
  assign n687 = n522 & ~n686;
  assign n688 = ~n679 & ~n687;
  assign n689 = n181 & ~n688;
  assign n690 = ~i_22_ & i_29_;
  assign n691 = n341 & n690;
  assign n692 = n311 & n691;
  assign n693 = n316 & n542;
  assign n694 = n180 & n693;
  assign n695 = ~n692 & ~n694;
  assign n696 = ~n689 & n695;
  assign n697 = n60 & n559;
  assign n698 = n651 & ~n697;
  assign n699 = ~n552 & n698;
  assign n700 = n89 & n508;
  assign n701 = ~n699 & n700;
  assign n702 = n696 & ~n701;
  assign n703 = ~n676 & n702;
  assign n704 = n177 & ~n703;
  assign n705 = n662 & ~n704;
  assign n706 = n66 & n680;
  assign n707 = n522 & n706;
  assign n708 = n568 & n665;
  assign n709 = ~n707 & ~n708;
  assign n710 = n598 & ~n709;
  assign n711 = ~i_0_ & ~i_7_;
  assign n712 = n46 & n711;
  assign n713 = n48 & n712;
  assign n714 = n382 & n713;
  assign n715 = n405 & n711;
  assign n716 = ~n296 & n715;
  assign n717 = ~n714 & ~n716;
  assign n718 = n519 & ~n717;
  assign n719 = ~n710 & ~n718;
  assign n720 = n61 & ~n719;
  assign n721 = n61 & n565;
  assign n722 = n598 & n721;
  assign n723 = n212 & n654;
  assign n724 = ~i_14_ & n476;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n722 & n725;
  assign n727 = ~i_35_ & ~n726;
  assign n728 = ~n720 & ~n727;
  assign n729 = n62 & n115;
  assign n730 = n192 & n729;
  assign n731 = ~i_29_ & ~i_30_;
  assign n732 = n211 & n731;
  assign n733 = n331 & n732;
  assign n734 = ~n730 & ~n733;
  assign n735 = ~i_35_ & n60;
  assign n736 = ~n232 & ~n735;
  assign n737 = ~i_33_ & n395;
  assign n738 = ~n736 & n737;
  assign n739 = n734 & ~n738;
  assign n740 = n728 & n739;
  assign n741 = ~i_32_ & ~n740;
  assign n742 = n56 & n278;
  assign n743 = n59 & n742;
  assign n744 = ~n226 & ~n743;
  assign n745 = n90 & ~n744;
  assign n746 = ~n505 & ~n745;
  assign n747 = n287 & ~n746;
  assign n748 = ~n253 & n533;
  assign n749 = n118 & n748;
  assign n750 = ~i_12_ & n715;
  assign n751 = ~n714 & ~n750;
  assign n752 = n519 & ~n751;
  assign n753 = ~n710 & ~n752;
  assign n754 = n437 & ~n753;
  assign n755 = n222 & n395;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n749 & n756;
  assign n758 = ~n747 & n757;
  assign n759 = ~i_33_ & ~n758;
  assign n760 = ~i_35_ & n559;
  assign n761 = ~n168 & ~n476;
  assign n762 = n760 & ~n761;
  assign n763 = n154 & n231;
  assign n764 = n227 & n513;
  assign n765 = n311 & ~n322;
  assign n766 = n457 & n540;
  assign n767 = n194 & n766;
  assign n768 = n765 & n767;
  assign n769 = ~n764 & ~n768;
  assign n770 = ~n763 & n769;
  assign n771 = ~n762 & n770;
  assign n772 = n101 & ~n610;
  assign n773 = ~i_33_ & n731;
  assign n774 = n234 & n297;
  assign n775 = ~i_27_ & n77;
  assign n776 = n774 & n775;
  assign n777 = n773 & n776;
  assign n778 = i_33_ & ~n729;
  assign n779 = n126 & ~n778;
  assign n780 = n243 & n255;
  assign n781 = n765 & n780;
  assign n782 = n91 & n781;
  assign n783 = ~n779 & ~n782;
  assign n784 = ~n777 & n783;
  assign n785 = ~n772 & n784;
  assign n786 = i_34_ & ~n785;
  assign n787 = n559 & n715;
  assign n788 = n565 & n760;
  assign n789 = ~i_8_ & ~i_33_;
  assign n790 = n712 & n789;
  assign n791 = n82 & n790;
  assign n792 = ~n788 & ~n791;
  assign n793 = n382 & ~n792;
  assign n794 = ~n787 & ~n793;
  assign n795 = n130 & n664;
  assign n796 = n96 & n795;
  assign n797 = ~n794 & n796;
  assign n798 = ~n786 & ~n797;
  assign n799 = n771 & n798;
  assign n800 = ~n759 & n799;
  assign n801 = ~n741 & n800;
  assign n802 = i_37_ & ~n801;
  assign n803 = n232 & n506;
  assign n804 = n91 & ~n225;
  assign n805 = n96 & n804;
  assign n806 = n647 & n805;
  assign n807 = ~n803 & ~n806;
  assign n808 = n559 & ~n807;
  assign n809 = ~i_24_ & ~i_30_;
  assign n810 = n261 & n809;
  assign n811 = n647 & n810;
  assign n812 = n550 & n811;
  assign n813 = ~i_30_ & n774;
  assign n814 = ~n222 & ~n813;
  assign n815 = n624 & ~n814;
  assign n816 = ~n812 & ~n815;
  assign n817 = ~n808 & n816;
  assign n818 = n90 & ~n817;
  assign n819 = n90 & n647;
  assign n820 = ~n536 & ~n819;
  assign n821 = n444 & ~n820;
  assign n822 = n608 & n821;
  assign n823 = n581 & n781;
  assign n824 = ~n822 & ~n823;
  assign n825 = n387 & ~n820;
  assign n826 = n262 & n613;
  assign n827 = ~n825 & ~n826;
  assign n828 = n149 & ~n827;
  assign n829 = n77 & n302;
  assign n830 = n53 & n335;
  assign n831 = n829 & n830;
  assign n832 = n508 & n789;
  assign n833 = n71 & n832;
  assign n834 = n79 & n833;
  assign n835 = ~n831 & ~n834;
  assign n836 = i_34_ & ~n835;
  assign n837 = ~n828 & ~n836;
  assign n838 = ~i_30_ & ~n837;
  assign n839 = n340 & n631;
  assign n840 = ~n838 & ~n839;
  assign n841 = n824 & n840;
  assign n842 = ~n818 & n841;
  assign n843 = n518 & n593;
  assign n844 = ~n667 & ~n843;
  assign n845 = n62 & ~n844;
  assign n846 = ~i_33_ & n593;
  assign n847 = n83 & n846;
  assign n848 = ~n845 & ~n847;
  assign n849 = n520 & ~n848;
  assign n850 = n195 & n288;
  assign n851 = n165 & n850;
  assign n852 = n61 & ~n820;
  assign n853 = n804 & n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = ~n849 & n854;
  assign n856 = ~i_32_ & ~n855;
  assign n857 = n387 & n773;
  assign n858 = n230 & n857;
  assign n859 = ~i_29_ & n559;
  assign n860 = n805 & n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = n508 & ~n861;
  assign n863 = ~n467 & ~n862;
  assign n864 = n158 & ~n863;
  assign n865 = ~n856 & ~n864;
  assign n866 = n842 & n865;
  assign n867 = ~n802 & n866;
  assign o_1_ = ~n705 | ~n867;
  assign n869 = n123 & n223;
  assign n870 = ~n95 & n220;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n514 & n871;
  assign n873 = n580 & ~n872;
  assign n874 = ~i_30_ & n89;
  assign n875 = i_8_ & i_32_;
  assign n876 = ~i_7_ & ~n875;
  assign n877 = n874 & n876;
  assign n878 = n178 & n653;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~n302 & ~n879;
  assign n881 = ~n873 & ~n880;
  assign n882 = ~i_24_ & i_38_;
  assign n883 = ~n881 & n882;
  assign n884 = ~n378 & ~n883;
  assign n885 = ~i_25_ & n89;
  assign n886 = i_38_ & n206;
  assign n887 = ~i_35_ & n886;
  assign n888 = ~i_10_ & ~i_24_;
  assign n889 = i_9_ & n888;
  assign n890 = n887 & n889;
  assign n891 = i_38_ & ~n871;
  assign n892 = ~i_35_ & i_38_;
  assign n893 = n51 & n892;
  assign n894 = n223 & n893;
  assign n895 = ~n891 & ~n894;
  assign n896 = ~i_24_ & ~n895;
  assign n897 = ~n890 & ~n896;
  assign n898 = n885 & ~n897;
  assign n899 = ~n49 & ~n56;
  assign n900 = ~n302 & n893;
  assign n901 = ~n899 & n900;
  assign n902 = ~i_30_ & n892;
  assign n903 = i_9_ & ~i_10_;
  assign n904 = n789 & n903;
  assign n905 = n902 & n904;
  assign n906 = i_31_ & ~n310;
  assign n907 = ~n905 & ~n906;
  assign n908 = ~n901 & n907;
  assign n909 = ~i_29_ & ~n908;
  assign n910 = ~n310 & ~n340;
  assign n911 = ~i_23_ & ~n910;
  assign n912 = i_22_ & ~n911;
  assign n913 = ~i_8_ & i_9_;
  assign n914 = ~i_10_ & n913;
  assign n915 = n892 & n914;
  assign n916 = ~n893 & ~n915;
  assign n917 = ~i_25_ & n731;
  assign n918 = ~n916 & n917;
  assign n919 = ~n912 & ~n918;
  assign n920 = ~n909 & n919;
  assign n921 = n77 & ~n920;
  assign n922 = ~i_33_ & n892;
  assign n923 = n78 & n340;
  assign n924 = n223 & n386;
  assign n925 = n504 & n924;
  assign n926 = ~n923 & ~n925;
  assign n927 = n922 & ~n926;
  assign n928 = ~n921 & ~n927;
  assign n929 = ~n898 & n928;
  assign n930 = n884 & n929;
  assign n931 = i_34_ & ~n930;
  assign n932 = ~i_26_ & n89;
  assign n933 = ~i_24_ & ~i_25_;
  assign n934 = n53 & n223;
  assign n935 = i_11_ & ~i_13_;
  assign n936 = ~n67 & n935;
  assign n937 = ~n899 & n913;
  assign n938 = n936 & n937;
  assign n939 = ~n934 & ~n938;
  assign n940 = ~i_30_ & n51;
  assign n941 = n939 & ~n940;
  assign n942 = n892 & ~n941;
  assign n943 = ~i_32_ & n892;
  assign n944 = ~n899 & n903;
  assign n945 = n943 & n944;
  assign n946 = i_38_ & n123;
  assign n947 = ~n893 & ~n946;
  assign n948 = n653 & ~n947;
  assign n949 = ~n945 & ~n948;
  assign n950 = ~n942 & n949;
  assign n951 = n933 & ~n950;
  assign n952 = i_38_ & n457;
  assign n953 = ~n891 & ~n952;
  assign n954 = ~i_24_ & ~n953;
  assign n955 = ~i_24_ & ~n899;
  assign n956 = n915 & n955;
  assign n957 = ~n890 & ~n956;
  assign n958 = ~n954 & n957;
  assign n959 = ~i_33_ & ~n958;
  assign n960 = ~i_31_ & n922;
  assign n961 = n924 & n960;
  assign n962 = ~n959 & ~n961;
  assign n963 = ~n951 & n962;
  assign n964 = n932 & ~n963;
  assign n965 = ~n931 & ~n964;
  assign n966 = ~i_22_ & n130;
  assign n967 = n144 & n966;
  assign n968 = n922 & n967;
  assign n969 = ~i_28_ & n966;
  assign n970 = ~i_25_ & n969;
  assign n971 = n902 & n970;
  assign n972 = ~n968 & ~n971;
  assign n973 = ~i_3_ & ~i_13_;
  assign n974 = ~n66 & n973;
  assign n975 = i_12_ & n974;
  assign n976 = ~i_13_ & i_18_;
  assign n977 = ~n66 & n976;
  assign n978 = i_2_ & ~i_12_;
  assign n979 = n977 & ~n978;
  assign n980 = ~n975 & ~n979;
  assign n981 = n913 & ~n980;
  assign n982 = ~n972 & n981;
  assign n983 = ~i_32_ & n968;
  assign n984 = n886 & n970;
  assign n985 = ~i_35_ & n984;
  assign n986 = ~n983 & ~n985;
  assign n987 = ~i_10_ & ~n978;
  assign n988 = ~n986 & n987;
  assign n989 = ~i_33_ & i_38_;
  assign n990 = n966 & n989;
  assign n991 = n180 & n990;
  assign n992 = ~n984 & ~n991;
  assign n993 = ~i_7_ & ~n992;
  assign n994 = i_12_ & n993;
  assign n995 = ~i_25_ & n932;
  assign n996 = i_34_ & n580;
  assign n997 = ~n995 & ~n996;
  assign n998 = n887 & ~n997;
  assign n999 = ~i_35_ & n250;
  assign n1000 = ~i_25_ & n999;
  assign n1001 = ~i_26_ & n760;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = i_38_ & n874;
  assign n1004 = ~n1002 & n1003;
  assign n1005 = ~n998 & ~n1004;
  assign n1006 = i_18_ & n935;
  assign n1007 = ~n974 & ~n1006;
  assign n1008 = ~n1005 & ~n1007;
  assign n1009 = ~i_24_ & n1008;
  assign n1010 = ~n994 & ~n1009;
  assign n1011 = n72 & n974;
  assign n1012 = ~n972 & n1011;
  assign n1013 = i_12_ & ~i_24_;
  assign n1014 = ~i_22_ & n1013;
  assign n1015 = ~i_26_ & ~i_28_;
  assign n1016 = ~n302 & n1015;
  assign n1017 = n952 & n1016;
  assign n1018 = n1014 & n1017;
  assign n1019 = n943 & n1016;
  assign n1020 = n809 & n1019;
  assign n1021 = ~i_22_ & n1020;
  assign n1022 = ~n980 & n1021;
  assign n1023 = ~n1018 & ~n1022;
  assign n1024 = ~n1012 & n1023;
  assign n1025 = n1010 & n1024;
  assign n1026 = ~n988 & n1025;
  assign n1027 = i_9_ & ~n1026;
  assign n1028 = ~n982 & ~n1027;
  assign n1029 = n933 & n1015;
  assign n1030 = n255 & n1029;
  assign n1031 = ~n302 & n386;
  assign n1032 = n932 & n1031;
  assign n1033 = n89 & n150;
  assign n1034 = n559 & n1033;
  assign n1035 = ~n1032 & ~n1034;
  assign n1036 = ~i_30_ & ~n1035;
  assign n1037 = ~n1030 & ~n1036;
  assign n1038 = n903 & ~n1037;
  assign n1039 = n51 & ~n899;
  assign n1040 = ~i_24_ & n932;
  assign n1041 = ~i_25_ & n1040;
  assign n1042 = ~n970 & ~n1041;
  assign n1043 = n1039 & ~n1042;
  assign n1044 = n914 & n995;
  assign n1045 = ~n53 & ~n1044;
  assign n1046 = ~i_28_ & i_34_;
  assign n1047 = ~i_29_ & n1046;
  assign n1048 = ~n932 & ~n1047;
  assign n1049 = ~n302 & ~n1048;
  assign n1050 = n955 & n1049;
  assign n1051 = ~n1045 & n1050;
  assign n1052 = ~n1043 & ~n1051;
  assign n1053 = ~n973 & ~n976;
  assign n1054 = i_19_ & ~i_24_;
  assign n1055 = ~i_25_ & n1054;
  assign n1056 = ~n1048 & n1055;
  assign n1057 = ~i_22_ & n1016;
  assign n1058 = n1054 & n1057;
  assign n1059 = ~n130 & ~n150;
  assign n1060 = n580 & ~n1059;
  assign n1061 = ~n66 & n1060;
  assign n1062 = n933 & n1047;
  assign n1063 = i_11_ & n1062;
  assign n1064 = ~n1061 & ~n1063;
  assign n1065 = ~n1058 & n1064;
  assign n1066 = ~n1056 & n1065;
  assign n1067 = n937 & ~n1066;
  assign n1068 = ~n1053 & n1067;
  assign n1069 = n1052 & ~n1068;
  assign n1070 = ~n1038 & n1069;
  assign n1071 = n892 & ~n1070;
  assign n1072 = ~n894 & n953;
  assign n1073 = n1041 & ~n1072;
  assign n1074 = n123 & ~n899;
  assign n1075 = ~n458 & ~n1074;
  assign n1076 = n990 & ~n1075;
  assign n1077 = ~n317 & ~n340;
  assign n1078 = n146 & n1077;
  assign n1079 = ~n322 & ~n1078;
  assign n1080 = i_22_ & ~n1079;
  assign n1081 = ~n151 & n1080;
  assign n1082 = ~n1076 & ~n1081;
  assign n1083 = ~i_28_ & ~n1082;
  assign n1084 = ~n1073 & ~n1083;
  assign n1085 = ~n1071 & n1084;
  assign n1086 = i_27_ & n137;
  assign n1087 = n966 & n1086;
  assign n1088 = ~i_25_ & n892;
  assign n1089 = n53 & n1088;
  assign n1090 = ~i_33_ & ~n947;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~i_30_ & n1040;
  assign n1093 = ~n1091 & n1092;
  assign n1094 = ~n310 & n1033;
  assign n1095 = ~n206 & n1094;
  assign n1096 = ~n1093 & ~n1095;
  assign n1097 = ~n1087 & n1096;
  assign n1098 = n130 & n922;
  assign n1099 = n150 & n1088;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n504 & ~n1100;
  assign n1102 = n960 & n1033;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n875 & ~n1103;
  assign n1105 = i_38_ & n760;
  assign n1106 = n969 & n1105;
  assign n1107 = ~i_31_ & n1106;
  assign n1108 = ~n969 & ~n1040;
  assign n1109 = n1089 & ~n1108;
  assign n1110 = ~n1107 & ~n1109;
  assign n1111 = ~n1104 & n1110;
  assign n1112 = n653 & ~n1111;
  assign n1113 = n1097 & ~n1112;
  assign n1114 = n885 & ~n1059;
  assign n1115 = ~n970 & ~n1114;
  assign n1116 = ~n1060 & n1115;
  assign n1117 = n943 & ~n1116;
  assign n1118 = ~n1106 & ~n1117;
  assign n1119 = ~i_2_ & i_9_;
  assign n1120 = n55 & n1119;
  assign n1121 = n977 & n1120;
  assign n1122 = i_3_ & ~n49;
  assign n1123 = i_9_ & ~i_13_;
  assign n1124 = n68 & n1123;
  assign n1125 = ~n899 & n1124;
  assign n1126 = ~n1122 & n1125;
  assign n1127 = ~n1121 & ~n1126;
  assign n1128 = ~n1118 & ~n1127;
  assign n1129 = ~n350 & n1077;
  assign n1130 = ~i_28_ & n1129;
  assign n1131 = ~n1128 & ~n1130;
  assign n1132 = ~n148 & ~n193;
  assign n1133 = n322 & ~n1132;
  assign n1134 = n914 & n1014;
  assign n1135 = ~i_22_ & n888;
  assign n1136 = n72 & n1135;
  assign n1137 = i_9_ & n1136;
  assign n1138 = ~n1134 & ~n1137;
  assign n1139 = ~i_26_ & n144;
  assign n1140 = ~n1138 & n1139;
  assign n1141 = n1088 & n1140;
  assign n1142 = ~n95 & n989;
  assign n1143 = ~i_32_ & n1040;
  assign n1144 = n118 & n1143;
  assign n1145 = n1142 & n1144;
  assign n1146 = ~n315 & ~n1145;
  assign n1147 = ~n1141 & n1146;
  assign n1148 = ~n1133 & n1147;
  assign n1149 = n1131 & n1148;
  assign n1150 = n1113 & n1149;
  assign n1151 = ~i_3_ & n1119;
  assign n1152 = n1020 & n1151;
  assign n1153 = ~i_13_ & ~i_22_;
  assign n1154 = n1152 & n1153;
  assign n1155 = i_19_ & n1154;
  assign n1156 = n1150 & ~n1155;
  assign n1157 = n1085 & n1156;
  assign n1158 = n1028 & n1157;
  assign n1159 = n936 & n1018;
  assign n1160 = n952 & n1058;
  assign n1161 = n976 & n1160;
  assign n1162 = ~n974 & ~n977;
  assign n1163 = ~i_31_ & n1029;
  assign n1164 = n887 & n1163;
  assign n1165 = n145 & n1098;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = ~i_22_ & ~n1166;
  assign n1168 = n51 & ~n972;
  assign n1169 = ~n993 & ~n1168;
  assign n1170 = ~n1167 & n1169;
  assign n1171 = ~n1162 & ~n1170;
  assign n1172 = ~n1161 & ~n1171;
  assign n1173 = i_12_ & ~n1172;
  assign n1174 = ~n1159 & ~n1173;
  assign n1175 = i_10_ & ~n1174;
  assign n1176 = i_12_ & n95;
  assign n1177 = ~i_3_ & n1176;
  assign n1178 = n1160 & n1177;
  assign n1179 = ~n302 & n1047;
  assign n1180 = n956 & n1179;
  assign n1181 = i_9_ & i_12_;
  assign n1182 = n1168 & n1181;
  assign n1183 = n346 & n513;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = i_18_ & n1054;
  assign n1186 = n1123 & n1185;
  assign n1187 = ~n1005 & n1186;
  assign n1188 = n1184 & ~n1187;
  assign n1189 = ~n1180 & n1188;
  assign n1190 = ~i_35_ & n1039;
  assign n1191 = ~n514 & ~n1190;
  assign n1192 = ~n1108 & ~n1191;
  assign n1193 = n944 & n1143;
  assign n1194 = ~n1140 & ~n1193;
  assign n1195 = ~i_35_ & ~n1194;
  assign n1196 = ~n1192 & ~n1195;
  assign n1197 = n989 & ~n1196;
  assign n1198 = n85 & ~n947;
  assign n1199 = n1016 & n1198;
  assign n1200 = n1019 & n1120;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = n1135 & ~n1201;
  assign n1203 = n177 & n692;
  assign n1204 = n902 & n1031;
  assign n1205 = n1124 & n1204;
  assign n1206 = ~n1048 & n1205;
  assign n1207 = ~n1203 & ~n1206;
  assign n1208 = ~n1202 & n1207;
  assign n1209 = ~n1197 & n1208;
  assign n1210 = n1189 & n1209;
  assign n1211 = ~n1178 & n1210;
  assign n1212 = ~n1175 & n1211;
  assign n1213 = n1158 & n1212;
  assign n1214 = n965 & n1213;
  assign n1215 = i_13_ & n1199;
  assign n1216 = n134 & ~n899;
  assign n1217 = ~i_35_ & n938;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n1016 & ~n1218;
  assign n1220 = ~i_31_ & n1015;
  assign n1221 = n223 & n760;
  assign n1222 = n1220 & n1221;
  assign n1223 = ~n1219 & ~n1222;
  assign n1224 = i_38_ & ~n1223;
  assign n1225 = n162 & n1220;
  assign n1226 = n1105 & n1225;
  assign n1227 = n49 & n1019;
  assign n1228 = n903 & n1227;
  assign n1229 = i_29_ & n1046;
  assign n1230 = ~n422 & n1229;
  assign n1231 = ~n1228 & ~n1230;
  assign n1232 = ~n1226 & n1231;
  assign n1233 = ~n1224 & n1232;
  assign n1234 = ~n1215 & n1233;
  assign n1235 = ~i_22_ & ~n1234;
  assign n1236 = n945 & n1179;
  assign n1237 = ~n934 & ~n940;
  assign n1238 = n922 & ~n1237;
  assign n1239 = ~i_23_ & ~n1238;
  assign n1240 = ~i_29_ & ~n1239;
  assign n1241 = ~i_16_ & ~i_27_;
  assign n1242 = ~n340 & ~n1241;
  assign n1243 = ~n1240 & ~n1242;
  assign n1244 = ~n690 & n1046;
  assign n1245 = ~n1243 & n1244;
  assign n1246 = ~n1236 & ~n1245;
  assign n1247 = ~n1235 & n1246;
  assign n1248 = ~i_24_ & ~n1247;
  assign n1249 = n223 & n1089;
  assign n1250 = i_29_ & ~n316;
  assign n1251 = ~i_31_ & n943;
  assign n1252 = ~n915 & ~n1251;
  assign n1253 = ~n899 & ~n1252;
  assign n1254 = n162 & ~n947;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = n895 & n1255;
  assign n1257 = ~n302 & ~n1256;
  assign n1258 = ~n1250 & ~n1257;
  assign n1259 = ~n1249 & n1258;
  assign n1260 = n193 & ~n1259;
  assign n1261 = ~n1166 & n1181;
  assign n1262 = n935 & n1152;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n318 & ~n422;
  assign n1265 = ~i_2_ & n1164;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n1263 & n1266;
  assign n1268 = ~n1260 & n1267;
  assign n1269 = ~i_22_ & ~n1268;
  assign n1270 = n653 & n876;
  assign n1271 = ~n1216 & ~n1270;
  assign n1272 = n885 & ~n1271;
  assign n1273 = i_30_ & ~n223;
  assign n1274 = n580 & n653;
  assign n1275 = n1273 & ~n1274;
  assign n1276 = ~n1074 & n1275;
  assign n1277 = ~n302 & n876;
  assign n1278 = ~n1276 & n1277;
  assign n1279 = n89 & n1278;
  assign n1280 = ~n1272 & ~n1279;
  assign n1281 = n146 & ~n1280;
  assign n1282 = n809 & ~n1002;
  assign n1283 = n130 & n1221;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = n504 & ~n1284;
  assign n1286 = n458 & n970;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = n362 & n932;
  assign n1289 = ~n1216 & ~n1288;
  assign n1290 = ~n1048 & ~n1289;
  assign n1291 = n223 & n999;
  assign n1292 = n504 & n1291;
  assign n1293 = ~n1290 & ~n1292;
  assign n1294 = n933 & ~n1293;
  assign n1295 = ~n406 & n580;
  assign n1296 = n1216 & n1295;
  assign n1297 = n514 & ~n1115;
  assign n1298 = ~n1074 & ~n1297;
  assign n1299 = ~n1116 & ~n1298;
  assign n1300 = ~n1296 & ~n1299;
  assign n1301 = ~n1294 & n1300;
  assign n1302 = n1287 & n1301;
  assign n1303 = ~n1281 & n1302;
  assign n1304 = i_38_ & ~n1303;
  assign n1305 = ~n1269 & ~n1304;
  assign n1306 = ~n1248 & n1305;
  assign o_2_ = ~n1214 | ~n1306;
endmodule


