// Benchmark "alu4_cl" written by ABC on Tue May 16 16:07:44 2017

module alu4_cl ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    o, p, q, r, s, t, u, v  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output o, p, q, r, s, t, u, v;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
    n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n473, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n638, n639, n640,
    n641, n642, n643;
  assign n23 = i & ~j;
  assign n24 = ~k & n23;
  assign n25 = ~n & n24;
  assign n26 = ~a & e;
  assign n27 = a & e;
  assign n28 = ~a & ~n26;
  assign n29 = ~n27 & ~n28;
  assign n30 = ~i & j;
  assign n31 = n & n30;
  assign n32 = ~j & ~n;
  assign n33 = l & n32;
  assign n34 = k & ~l;
  assign n35 = i & j;
  assign n36 = n34 & n35;
  assign n37 = i & k;
  assign n38 = n33 & n37;
  assign n39 = n31 & ~n34;
  assign n40 = ~n36 & ~n39;
  assign n41 = ~n38 & n40;
  assign n42 = ~i & ~k;
  assign n43 = ~n & n42;
  assign n44 = n33 & n43;
  assign n45 = ~l & n43;
  assign n46 = ~n44 & ~n45;
  assign n47 = ~i & k;
  assign n48 = i & ~k;
  assign n49 = ~l & n48;
  assign n50 = ~n47 & ~n49;
  assign n51 = ~j & n50;
  assign n52 = n25 & ~n50;
  assign n53 = k & n;
  assign n54 = n51 & n53;
  assign n55 = ~n52 & ~n54;
  assign n56 = ~k & l;
  assign n57 = n35 & n56;
  assign n58 = ~l & n30;
  assign n59 = ~n57 & ~n58;
  assign n60 = ~n42 & ~n59;
  assign n61 = n & n60;
  assign n62 = ~i & ~j;
  assign n63 = l & n62;
  assign n64 = k & l;
  assign n65 = ~n35 & n64;
  assign n66 = ~n63 & ~n65;
  assign n67 = n & ~n66;
  assign n68 = n35 & n61;
  assign n69 = n34 & n62;
  assign n70 = ~k & n67;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n68 & n71;
  assign n73 = n29 & n41;
  assign n74 = n31 & n73;
  assign n75 = ~a & ~n46;
  assign n76 = n29 & ~n55;
  assign n77 = n27 & ~n72;
  assign n78 = a & ~n55;
  assign n79 = ~e & ~n41;
  assign n80 = ~n78 & ~n79;
  assign n81 = ~n77 & n80;
  assign n82 = ~n76 & n81;
  assign n83 = ~n75 & n82;
  assign n84 = ~n74 & n83;
  assign n85 = ~n42 & ~n64;
  assign n86 = k & ~n;
  assign n87 = ~n85 & n86;
  assign n88 = n & n34;
  assign n89 = k & n35;
  assign n90 = n88 & n89;
  assign n91 = n35 & n88;
  assign n92 = a & ~n84;
  assign n93 = n62 & n88;
  assign n94 = n23 & n88;
  assign n95 = ~i & l;
  assign n96 = n & n95;
  assign n97 = j & n96;
  assign n98 = n91 & n92;
  assign n99 = n84 & n93;
  assign n100 = n27 & n94;
  assign n101 = a & n97;
  assign n102 = ~n84 & n97;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~n100 & n103;
  assign n105 = ~n99 & n104;
  assign n106 = ~n98 & n105;
  assign n107 = n & n24;
  assign n108 = ~l & n;
  assign n109 = ~n34 & ~n35;
  assign n110 = n108 & n109;
  assign n111 = n & n89;
  assign n112 = ~n85 & n111;
  assign n113 = ~n84 & ~n106;
  assign n114 = ~n67 & n113;
  assign n115 = ~n90 & n114;
  assign n116 = a & ~n27;
  assign n117 = n107 & n116;
  assign n118 = a & n84;
  assign n119 = n67 & n118;
  assign n120 = ~a & ~n84;
  assign n121 = n67 & n120;
  assign n122 = ~n84 & n110;
  assign n123 = a & n110;
  assign n124 = ~a & n112;
  assign n125 = n61 & n84;
  assign n126 = n90 & n106;
  assign n127 = n93 & n106;
  assign n128 = ~a & n93;
  assign n129 = n26 & n107;
  assign n130 = n84 & n94;
  assign n131 = ~n129 & ~n130;
  assign n132 = ~n128 & n131;
  assign n133 = ~n127 & n132;
  assign n134 = ~n126 & n133;
  assign n135 = ~n125 & n134;
  assign n136 = ~n124 & n135;
  assign n137 = ~n123 & n136;
  assign n138 = ~n122 & n137;
  assign n139 = ~n121 & n138;
  assign n140 = ~n119 & n139;
  assign n141 = ~n117 & n140;
  assign n142 = ~n115 & n141;
  assign n143 = n32 & ~n50;
  assign n144 = j & ~n;
  assign n145 = n95 & n144;
  assign n146 = n32 & ~n85;
  assign n147 = n34 & n55;
  assign n148 = n51 & n147;
  assign n149 = l & ~n;
  assign n150 = ~n24 & n149;
  assign n151 = n34 & ~n50;
  assign n152 = n144 & n151;
  assign n153 = ~k & n35;
  assign n154 = n108 & n153;
  assign n155 = k & n95;
  assign n156 = n32 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = ~n & ~n84;
  assign n159 = n29 & n158;
  assign n160 = ~n25 & n159;
  assign n161 = n29 & n33;
  assign n162 = ~n87 & n161;
  assign n163 = ~m & n;
  assign n164 = n142 & n163;
  assign n165 = n84 & n143;
  assign n166 = n26 & n145;
  assign n167 = a & n87;
  assign n168 = ~n84 & n146;
  assign n169 = ~e & n148;
  assign n170 = n27 & n150;
  assign n171 = ~n29 & n152;
  assign n172 = m & ~n142;
  assign n173 = n157 & ~n172;
  assign n174 = ~n171 & n173;
  assign n175 = ~n170 & n174;
  assign n176 = ~n169 & n175;
  assign n177 = ~n168 & n176;
  assign n178 = ~n167 & n177;
  assign n179 = ~n166 & n178;
  assign n180 = ~n165 & n179;
  assign n181 = ~n164 & n180;
  assign n182 = ~n162 & n181;
  assign o = n160 | ~n182;
  assign n184 = b & f;
  assign n185 = ~b & ~f;
  assign n186 = ~n184 & ~n185;
  assign n187 = b & ~f;
  assign n188 = ~b & f;
  assign n189 = n26 & ~n187;
  assign n190 = ~n188 & ~n189;
  assign n191 = ~j & n88;
  assign n192 = n72 & ~n191;
  assign n193 = a & ~n42;
  assign n194 = n96 & n193;
  assign n195 = ~n31 & n194;
  assign n196 = ~n26 & n41;
  assign n197 = n186 & n196;
  assign n198 = n31 & n197;
  assign n199 = n41 & ~n190;
  assign n200 = ~n186 & n199;
  assign n201 = n31 & n200;
  assign n202 = ~b & ~n46;
  assign n203 = n184 & ~n192;
  assign n204 = ~n55 & ~n185;
  assign n205 = ~f & ~n41;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n203 & n206;
  assign n208 = ~n202 & n207;
  assign n209 = ~n201 & n208;
  assign n210 = ~n198 & n209;
  assign n211 = ~n195 & n210;
  assign n212 = ~m & ~n142;
  assign n213 = ~b & n211;
  assign n214 = ~n42 & n84;
  assign n215 = ~k & n97;
  assign n216 = b & ~n211;
  assign n217 = n91 & n216;
  assign n218 = n97 & ~n213;
  assign n219 = n94 & n184;
  assign n220 = n93 & n211;
  assign n221 = ~n219 & ~n220;
  assign n222 = ~n218 & n221;
  assign n223 = ~n217 & n222;
  assign n224 = n184 & n215;
  assign n225 = n94 & n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = n223 & ~n226;
  assign n228 = ~n223 & n226;
  assign n229 = ~n227 & ~n228;
  assign n230 = n34 & ~n55;
  assign n231 = a & ~n106;
  assign n232 = ~n223 & ~n231;
  assign n233 = n223 & n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = n & ~n59;
  assign n236 = n92 & ~n213;
  assign n237 = ~n216 & ~n236;
  assign n238 = ~a & ~b;
  assign n239 = n84 & n211;
  assign n240 = n27 & n215;
  assign n241 = n94 & n106;
  assign n242 = ~n240 & ~n241;
  assign n243 = ~n106 & ~n242;
  assign n244 = ~n84 & ~n242;
  assign n245 = ~n211 & ~n226;
  assign n246 = ~n244 & ~n245;
  assign n247 = n106 & n223;
  assign n248 = n231 & n234;
  assign n249 = b & ~n234;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n27 & ~n184;
  assign n252 = ~n67 & n251;
  assign n253 = ~n229 & n252;
  assign n254 = ~n214 & n253;
  assign n255 = ~n213 & n254;
  assign n256 = ~n90 & n255;
  assign n257 = b & n234;
  assign n258 = ~n230 & n257;
  assign n259 = n108 & n258;
  assign n260 = ~n61 & n259;
  assign n261 = n27 & n107;
  assign n262 = ~n186 & n261;
  assign n263 = ~n108 & n262;
  assign n264 = a & ~n213;
  assign n265 = n112 & n264;
  assign n266 = n67 & n92;
  assign n267 = n216 & n266;
  assign n268 = n67 & n213;
  assign n269 = n92 & n268;
  assign n270 = n107 & n186;
  assign n271 = n108 & n270;
  assign n272 = ~n211 & ~n214;
  assign n273 = n235 & n272;
  assign n274 = n67 & n237;
  assign n275 = ~n213 & n274;
  assign n276 = ~n27 & n107;
  assign n277 = n186 & n276;
  assign n278 = n112 & n238;
  assign n279 = n61 & n239;
  assign n280 = n239 & n243;
  assign n281 = n230 & n246;
  assign n282 = n90 & n247;
  assign n283 = n93 & n250;
  assign n284 = ~n282 & ~n283;
  assign n285 = ~n281 & n284;
  assign n286 = ~n280 & n285;
  assign n287 = ~n279 & n286;
  assign n288 = ~n278 & n287;
  assign n289 = ~n277 & n288;
  assign n290 = ~n275 & n289;
  assign n291 = ~n273 & n290;
  assign n292 = ~n271 & n291;
  assign n293 = ~n269 & n292;
  assign n294 = ~n267 & n293;
  assign n295 = ~n265 & n294;
  assign n296 = ~n263 & n295;
  assign n297 = ~n260 & n296;
  assign n298 = ~n256 & n297;
  assign n299 = ~n & ~n211;
  assign n300 = n186 & n299;
  assign n301 = ~n25 & n300;
  assign n302 = n33 & n186;
  assign n303 = ~n87 & n302;
  assign n304 = n145 & n188;
  assign n305 = n143 & n211;
  assign n306 = b & n87;
  assign n307 = n146 & ~n211;
  assign n308 = ~f & n148;
  assign n309 = n150 & n184;
  assign n310 = n152 & ~n186;
  assign n311 = n212 & n298;
  assign n312 = ~n212 & ~n298;
  assign n313 = n157 & ~n312;
  assign n314 = ~n311 & n313;
  assign n315 = ~n310 & n314;
  assign n316 = ~n309 & n315;
  assign n317 = ~n308 & n316;
  assign n318 = ~n307 & n317;
  assign n319 = ~n306 & n318;
  assign n320 = ~n305 & n319;
  assign n321 = ~n304 & n320;
  assign n322 = ~n303 & n321;
  assign p = n301 | ~n322;
  assign n324 = ~c & ~g;
  assign n325 = c & g;
  assign n326 = c & ~g;
  assign n327 = c & n190;
  assign n328 = ~g & n190;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~n326 & n329;
  assign n331 = n41 & ~n325;
  assign n332 = n190 & n331;
  assign n333 = ~n324 & n332;
  assign n334 = n31 & n333;
  assign n335 = b & ~n42;
  assign n336 = n96 & n335;
  assign n337 = ~n31 & n336;
  assign n338 = n41 & n325;
  assign n339 = n330 & n338;
  assign n340 = n31 & n339;
  assign n341 = n324 & n330;
  assign n342 = n31 & n341;
  assign n343 = ~c & ~n46;
  assign n344 = ~n192 & n325;
  assign n345 = ~n55 & ~n324;
  assign n346 = ~g & ~n41;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n344 & n347;
  assign n349 = ~n343 & n348;
  assign n350 = ~n342 & n349;
  assign n351 = ~n340 & n350;
  assign n352 = ~n337 & n351;
  assign n353 = ~n334 & n352;
  assign n354 = n212 & ~n298;
  assign n355 = c & ~n353;
  assign n356 = ~c & n353;
  assign n357 = n91 & n355;
  assign n358 = n97 & ~n356;
  assign n359 = n94 & n325;
  assign n360 = n93 & n353;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n358 & n361;
  assign n363 = ~n357 & n362;
  assign n364 = n215 & n325;
  assign n365 = n94 & n363;
  assign n366 = ~n364 & ~n365;
  assign n367 = n363 & n366;
  assign n368 = ~n363 & ~n366;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n353 & ~n366;
  assign n371 = n353 & n366;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n223 & n243;
  assign n374 = ~n223 & ~n226;
  assign n375 = ~n373 & ~n374;
  assign n376 = n239 & n353;
  assign n377 = n27 & ~n185;
  assign n378 = ~n184 & ~n377;
  assign n379 = ~n324 & ~n378;
  assign n380 = ~n325 & ~n379;
  assign n381 = n59 & ~n62;
  assign n382 = n250 & ~n363;
  assign n383 = ~n250 & n363;
  assign n384 = ~n382 & ~n383;
  assign n385 = n211 & n214;
  assign n386 = ~n237 & ~n356;
  assign n387 = ~n355 & ~n386;
  assign n388 = n247 & n363;
  assign n389 = ~c & n238;
  assign n390 = n246 & n375;
  assign n391 = n372 & n390;
  assign n392 = ~n67 & n391;
  assign n393 = n369 & n392;
  assign n394 = ~n111 & n393;
  assign n395 = c & ~n238;
  assign n396 = n111 & n395;
  assign n397 = n376 & n396;
  assign n398 = n107 & ~n378;
  assign n399 = n324 & n398;
  assign n400 = ~n110 & n399;
  assign n401 = n107 & ~n380;
  assign n402 = n110 & n401;
  assign n403 = n111 & ~n247;
  assign n404 = n355 & n403;
  assign n405 = n67 & ~n237;
  assign n406 = n355 & n405;
  assign n407 = n356 & ~n384;
  assign n408 = ~n381 & n407;
  assign n409 = n372 & ~n385;
  assign n410 = n235 & n409;
  assign n411 = n356 & n405;
  assign n412 = n67 & n387;
  assign n413 = ~n356 & n412;
  assign n414 = n107 & n380;
  assign n415 = ~n324 & n414;
  assign n416 = n107 & n325;
  assign n417 = ~n378 & n416;
  assign n418 = c & n384;
  assign n419 = n93 & n418;
  assign n420 = n61 & n376;
  assign n421 = n110 & ~n356;
  assign n422 = n90 & n388;
  assign n423 = n111 & n389;
  assign n424 = ~n246 & ~n372;
  assign n425 = ~n369 & ~n375;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n423 & n426;
  assign n428 = ~n422 & n427;
  assign n429 = ~n421 & n428;
  assign n430 = ~n420 & n429;
  assign n431 = ~n419 & n430;
  assign n432 = ~n417 & n431;
  assign n433 = ~n415 & n432;
  assign n434 = ~n413 & n433;
  assign n435 = ~n411 & n434;
  assign n436 = ~n410 & n435;
  assign n437 = ~n408 & n436;
  assign n438 = ~n406 & n437;
  assign n439 = ~n404 & n438;
  assign n440 = ~n402 & n439;
  assign n441 = ~n400 & n440;
  assign n442 = ~n397 & n441;
  assign n443 = ~n394 & n442;
  assign n444 = ~n & ~n353;
  assign n445 = ~n324 & n444;
  assign n446 = ~n143 & n445;
  assign n447 = ~n324 & ~n325;
  assign n448 = n33 & n447;
  assign n449 = ~n87 & n448;
  assign n450 = n143 & n353;
  assign n451 = g & n145;
  assign n452 = c & n87;
  assign n453 = n146 & n324;
  assign n454 = ~g & n148;
  assign n455 = n150 & n325;
  assign n456 = n152 & n324;
  assign n457 = n152 & n325;
  assign n458 = n354 & n443;
  assign n459 = ~n354 & ~n443;
  assign n460 = n157 & ~n459;
  assign n461 = ~n458 & n460;
  assign n462 = ~n457 & n461;
  assign n463 = ~n456 & n462;
  assign n464 = ~n455 & n463;
  assign n465 = ~n454 & n464;
  assign n466 = ~n453 & n465;
  assign n467 = ~n452 & n466;
  assign n468 = ~n451 & n467;
  assign n469 = ~n450 & n468;
  assign n470 = ~n449 & n469;
  assign q = n446 | ~n470;
  assign t = d & h;
  assign n473 = ~d & ~h;
  assign s = t | n473;
  assign n475 = c & n;
  assign n476 = ~n50 & n475;
  assign n477 = n62 & n476;
  assign n478 = n72 & n477;
  assign n479 = n60 & s;
  assign n480 = n88 & n479;
  assign n481 = n330 & n480;
  assign n482 = n60 & ~s;
  assign n483 = n88 & n482;
  assign n484 = ~n330 & n483;
  assign n485 = ~d & n43;
  assign n486 = ~n381 & n485;
  assign n487 = ~n72 & t;
  assign n488 = ~n55 & t;
  assign n489 = ~n55 & ~s;
  assign n490 = ~h & ~n41;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~n488 & n491;
  assign n493 = ~n487 & n492;
  assign n494 = ~n486 & n493;
  assign n495 = ~n484 & n494;
  assign n496 = ~n481 & n495;
  assign n497 = ~n478 & n496;
  assign n498 = n354 & ~n443;
  assign n499 = d & ~n497;
  assign n500 = ~d & n497;
  assign n501 = n91 & n499;
  assign n502 = n97 & ~n500;
  assign n503 = n94 & t;
  assign n504 = n93 & n497;
  assign n505 = ~n503 & ~n504;
  assign n506 = ~n502 & n505;
  assign n507 = ~n501 & n506;
  assign n508 = n215 & t;
  assign n509 = n94 & n507;
  assign n510 = ~n508 & ~n509;
  assign n511 = n497 & n510;
  assign n512 = ~n497 & ~n510;
  assign n513 = ~n511 & ~n512;
  assign n514 = n507 & n510;
  assign n515 = ~n507 & ~n510;
  assign n516 = ~n514 & ~n515;
  assign n517 = ~n366 & ~n372;
  assign n518 = n246 & ~n517;
  assign n519 = ~n367 & ~n375;
  assign n520 = ~n368 & ~n519;
  assign n521 = ~d & n507;
  assign n522 = d & ~n507;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n250 & n384;
  assign n525 = c & ~n384;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n499 & ~n500;
  assign n528 = ~d & n;
  assign n529 = ~n85 & n528;
  assign n530 = n389 & n529;
  assign n531 = n88 & n507;
  assign n532 = n388 & n531;
  assign n533 = ~n530 & ~n532;
  assign n534 = n518 & n520;
  assign n535 = ~n67 & n534;
  assign n536 = n516 & n535;
  assign n537 = n513 & n536;
  assign n538 = ~n90 & n537;
  assign n539 = ~n380 & s;
  assign n540 = n107 & n539;
  assign n541 = ~n110 & n540;
  assign n542 = n61 & ~n513;
  assign n543 = n376 & n542;
  assign n544 = n107 & ~s;
  assign n545 = n110 & n544;
  assign n546 = ~n389 & n523;
  assign n547 = n112 & n546;
  assign n548 = ~n353 & n513;
  assign n549 = n61 & n548;
  assign n550 = n90 & n516;
  assign n551 = ~n388 & n550;
  assign n552 = ~n385 & n513;
  assign n553 = n235 & n552;
  assign n554 = n93 & n526;
  assign n555 = n523 & n554;
  assign n556 = n93 & ~n526;
  assign n557 = n527 & n556;
  assign n558 = n412 & n527;
  assign n559 = n67 & ~n387;
  assign n560 = ~n527 & n559;
  assign n561 = n380 & ~s;
  assign n562 = n107 & n561;
  assign n563 = n110 & n523;
  assign n564 = ~n513 & ~n518;
  assign n565 = n89 & ~n533;
  assign n566 = ~n516 & ~n520;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n564 & n567;
  assign n569 = ~n563 & n568;
  assign n570 = ~n562 & n569;
  assign n571 = ~n560 & n570;
  assign n572 = ~n558 & n571;
  assign n573 = ~n557 & n572;
  assign n574 = ~n555 & n573;
  assign n575 = ~n553 & n574;
  assign n576 = ~n551 & n575;
  assign n577 = ~n549 & n576;
  assign n578 = ~n547 & n577;
  assign n579 = ~n545 & n578;
  assign n580 = ~n543 & n579;
  assign n581 = ~n541 & n580;
  assign n582 = ~n538 & n581;
  assign n583 = ~n & ~s;
  assign n584 = ~n497 & n583;
  assign n585 = ~n143 & n584;
  assign n586 = n33 & ~s;
  assign n587 = ~n87 & n586;
  assign n588 = n143 & n497;
  assign n589 = h & n145;
  assign n590 = d & n87;
  assign n591 = n146 & ~n497;
  assign n592 = ~h & n148;
  assign n593 = n150 & t;
  assign n594 = n498 & n582;
  assign n595 = ~n498 & ~n582;
  assign n596 = n157 & ~n595;
  assign n597 = ~n594 & n596;
  assign n598 = n152 & s;
  assign n599 = n597 & ~n598;
  assign n600 = ~n593 & n599;
  assign n601 = ~n592 & n600;
  assign n602 = ~n591 & n601;
  assign n603 = ~n590 & n602;
  assign n604 = ~n589 & n603;
  assign n605 = ~n588 & n604;
  assign n606 = ~n587 & n605;
  assign r = n585 | ~n606;
  assign n608 = n & n85;
  assign n609 = n582 & n608;
  assign n610 = ~n89 & n609;
  assign n611 = ~n107 & n610;
  assign n612 = ~n235 & n611;
  assign n613 = n85 & n235;
  assign n614 = n511 & n613;
  assign n615 = n376 & n614;
  assign n616 = n & ~n85;
  assign n617 = n582 & n616;
  assign n618 = ~n511 & n617;
  assign n619 = d & n497;
  assign n620 = ~n507 & n619;
  assign n621 = ~n67 & n620;
  assign n622 = ~s & n582;
  assign n623 = n107 & n622;
  assign n624 = n50 & t;
  assign n625 = n107 & n624;
  assign n626 = d & ~n387;
  assign n627 = n67 & n626;
  assign n628 = n498 & ~n582;
  assign n629 = n518 & ~n565;
  assign n630 = ~n628 & n629;
  assign n631 = ~n627 & n630;
  assign n632 = ~n625 & n631;
  assign n633 = ~n623 & n632;
  assign n634 = ~n621 & n633;
  assign n635 = ~n618 & n634;
  assign n636 = ~n615 & n635;
  assign u = n612 | ~n636;
  assign n638 = ~n29 & s;
  assign n639 = ~n186 & n638;
  assign n640 = n324 & n639;
  assign n641 = n325 & s;
  assign n642 = ~n29 & n641;
  assign n643 = ~n186 & n642;
  assign v = n640 | n643;
endmodule


