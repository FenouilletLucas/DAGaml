// Benchmark "i3" written by ABC on Tue May 16 16:07:50 2017

module i3 ( 
    \V132(5) , \V28(13) , \V126(1) , \V88(21) , \V132(4) , \V28(12) ,
    \V126(0) , \V88(20) , \V28(15) , \V28(14) , \V132(1) , \V132(0) ,
    \V28(11) , \V88(27) , \V28(10) , \V88(0) , \V88(26) , \V88(1) ,
    \V88(29) , \V88(2) , \V88(28) , \V88(3) , \V88(4) , \V28(17) ,
    \V88(5) , \V120(31) , \V28(16) , \V88(6) , \V120(30) , \V56(13) ,
    \V28(19) , \V88(7) , \V56(12) , \V28(18) , \V88(8) , \V56(15) ,
    \V28(23) , \V88(9) , \V88(31) , \V56(14) , \V28(22) , \V88(30) ,
    \V28(25) , \V28(24) , \V56(11) , \V56(10) , \V28(21) , \V28(20) ,
    \V120(27) , \V120(26) , \V120(29) , \V56(17) , \V120(28) , \V120(3) ,
    \V56(0) , \V56(16) , \V120(2) , \V56(1) , \V56(19) , \V28(27) ,
    \V120(5) , \V56(2) , \V56(18) , \V28(26) , \V120(4) , \V56(3) ,
    \V56(23) , \V56(4) , \V56(22) , \V56(5) , \V56(25) , \V120(1) ,
    \V56(6) , \V56(24) , \V120(21) , \V120(0) , \V56(7) , \V120(20) ,
    \V56(8) , \V120(23) , \V56(9) , \V56(21) , \V120(22) , \V56(20) ,
    \V120(25) , \V120(24) , \V120(7) , \V120(17) , \V120(6) , \V120(16) ,
    \V120(9) , \V120(19) , \V120(8) , \V56(27) , \V120(18) , \V56(26) ,
    \V88(13) , \V28(0) , \V88(12) , \V28(1) , \V88(15) , \V120(11) ,
    \V28(2) , \V88(14) , \V120(10) , \V28(3) , \V120(13) , \V28(4) ,
    \V120(12) , \V28(5) , \V88(11) , \V120(15) , \V28(6) , \V88(10) ,
    \V120(14) , \V28(7) , \V28(8) , \V28(9) , \V88(17) , \V88(16) ,
    \V88(19) , \V88(18) , \V126(3) , \V88(23) , \V126(2) , \V88(22) ,
    \V126(5) , \V88(25) , \V126(4) , \V88(24) , \V132(3) , \V132(2) ,
    \V138(3) , \V138(2) , \V134(1) , \V134(0) , \V138(1) , \V138(0)   );
  input  \V132(5) , \V28(13) , \V126(1) , \V88(21) , \V132(4) ,
    \V28(12) , \V126(0) , \V88(20) , \V28(15) , \V28(14) , \V132(1) ,
    \V132(0) , \V28(11) , \V88(27) , \V28(10) , \V88(0) , \V88(26) ,
    \V88(1) , \V88(29) , \V88(2) , \V88(28) , \V88(3) , \V88(4) ,
    \V28(17) , \V88(5) , \V120(31) , \V28(16) , \V88(6) , \V120(30) ,
    \V56(13) , \V28(19) , \V88(7) , \V56(12) , \V28(18) , \V88(8) ,
    \V56(15) , \V28(23) , \V88(9) , \V88(31) , \V56(14) , \V28(22) ,
    \V88(30) , \V28(25) , \V28(24) , \V56(11) , \V56(10) , \V28(21) ,
    \V28(20) , \V120(27) , \V120(26) , \V120(29) , \V56(17) , \V120(28) ,
    \V120(3) , \V56(0) , \V56(16) , \V120(2) , \V56(1) , \V56(19) ,
    \V28(27) , \V120(5) , \V56(2) , \V56(18) , \V28(26) , \V120(4) ,
    \V56(3) , \V56(23) , \V56(4) , \V56(22) , \V56(5) , \V56(25) ,
    \V120(1) , \V56(6) , \V56(24) , \V120(21) , \V120(0) , \V56(7) ,
    \V120(20) , \V56(8) , \V120(23) , \V56(9) , \V56(21) , \V120(22) ,
    \V56(20) , \V120(25) , \V120(24) , \V120(7) , \V120(17) , \V120(6) ,
    \V120(16) , \V120(9) , \V120(19) , \V120(8) , \V56(27) , \V120(18) ,
    \V56(26) , \V88(13) , \V28(0) , \V88(12) , \V28(1) , \V88(15) ,
    \V120(11) , \V28(2) , \V88(14) , \V120(10) , \V28(3) , \V120(13) ,
    \V28(4) , \V120(12) , \V28(5) , \V88(11) , \V120(15) , \V28(6) ,
    \V88(10) , \V120(14) , \V28(7) , \V28(8) , \V28(9) , \V88(17) ,
    \V88(16) , \V88(19) , \V88(18) , \V126(3) , \V88(23) , \V126(2) ,
    \V88(22) , \V126(5) , \V88(25) , \V126(4) , \V88(24) , \V132(3) ,
    \V132(2) ;
  output \V138(3) , \V138(2) , \V134(1) , \V134(0) , \V138(1) , \V138(0) ;
  wire n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263;
  assign n139 = ~\V126(1)  & ~\V132(1) ;
  assign n140 = ~\V126(0)  & ~\V132(0) ;
  assign n141 = ~\V120(30)  & ~\V88(30) ;
  assign n142 = ~\V120(31)  & ~\V88(31) ;
  assign n143 = ~\V88(29)  & ~\V120(29) ;
  assign n144 = ~\V88(27)  & ~\V120(27) ;
  assign n145 = ~\V88(26)  & ~\V120(26) ;
  assign n146 = ~\V88(28)  & ~\V120(28) ;
  assign n147 = ~\V120(23)  & ~\V88(23) ;
  assign n148 = ~\V120(22)  & ~\V88(22) ;
  assign n149 = ~\V120(24)  & ~\V88(24) ;
  assign n150 = ~\V120(25)  & ~\V88(25) ;
  assign n151 = ~\V126(3)  & ~\V132(3) ;
  assign n152 = ~\V126(2)  & ~\V132(2) ;
  assign n153 = ~\V132(4)  & ~\V126(4) ;
  assign n154 = ~\V132(5)  & ~\V126(5) ;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n152 & n155;
  assign n157 = ~n151 & n156;
  assign n158 = ~n150 & n157;
  assign n159 = ~n149 & n158;
  assign n160 = ~n148 & n159;
  assign n161 = ~n147 & n160;
  assign n162 = ~n146 & n161;
  assign n163 = ~n145 & n162;
  assign n164 = ~n144 & n163;
  assign n165 = ~n143 & n164;
  assign n166 = ~n142 & n165;
  assign n167 = ~n141 & n166;
  assign n168 = ~n140 & n167;
  assign \V138(3)  = ~n139 & n168;
  assign n170 = ~\V120(17)  & ~\V88(17) ;
  assign n171 = ~\V120(16)  & ~\V88(16) ;
  assign n172 = ~\V88(14)  & ~\V120(14) ;
  assign n173 = ~\V88(15)  & ~\V120(15) ;
  assign n174 = ~\V88(13)  & ~\V120(13) ;
  assign n175 = ~\V120(11)  & ~\V88(11) ;
  assign n176 = ~\V120(10)  & ~\V88(10) ;
  assign n177 = ~\V88(12)  & ~\V120(12) ;
  assign n178 = ~\V88(7)  & ~\V120(7) ;
  assign n179 = ~\V88(6)  & ~\V120(6) ;
  assign n180 = ~\V88(8)  & ~\V120(8) ;
  assign n181 = ~\V88(9)  & ~\V120(9) ;
  assign n182 = ~\V120(19)  & ~\V88(19) ;
  assign n183 = ~\V120(18)  & ~\V88(18) ;
  assign n184 = ~\V88(20)  & ~\V120(20) ;
  assign n185 = ~\V88(21)  & ~\V120(21) ;
  assign n186 = ~n184 & ~n185;
  assign n187 = ~n183 & n186;
  assign n188 = ~n182 & n187;
  assign n189 = ~n181 & n188;
  assign n190 = ~n180 & n189;
  assign n191 = ~n179 & n190;
  assign n192 = ~n178 & n191;
  assign n193 = ~n177 & n192;
  assign n194 = ~n176 & n193;
  assign n195 = ~n175 & n194;
  assign n196 = ~n174 & n195;
  assign n197 = ~n173 & n196;
  assign n198 = ~n172 & n197;
  assign n199 = ~n171 & n198;
  assign \V138(2)  = ~n170 & n199;
  assign \V134(1)  = \V56(1)  | \V28(1) ;
  assign \V134(0)  = \V56(0)  | \V28(0) ;
  assign n203 = ~\V88(1)  & ~\V120(1) ;
  assign n204 = ~\V88(0)  & ~\V120(0) ;
  assign n205 = ~\V28(26)  & ~\V56(26) ;
  assign n206 = ~\V28(27)  & ~\V56(27) ;
  assign n207 = ~\V28(25)  & ~\V56(25) ;
  assign n208 = ~\V28(23)  & ~\V56(23) ;
  assign n209 = ~\V28(22)  & ~\V56(22) ;
  assign n210 = ~\V28(24)  & ~\V56(24) ;
  assign n211 = ~\V28(19)  & ~\V56(19) ;
  assign n212 = ~\V28(18)  & ~\V56(18) ;
  assign n213 = ~\V28(20)  & ~\V56(20) ;
  assign n214 = ~\V28(21)  & ~\V56(21) ;
  assign n215 = ~\V88(3)  & ~\V120(3) ;
  assign n216 = ~\V88(2)  & ~\V120(2) ;
  assign n217 = ~\V88(4)  & ~\V120(4) ;
  assign n218 = ~\V88(5)  & ~\V120(5) ;
  assign n219 = ~n217 & ~n218;
  assign n220 = ~n216 & n219;
  assign n221 = ~n215 & n220;
  assign n222 = ~n214 & n221;
  assign n223 = ~n213 & n222;
  assign n224 = ~n212 & n223;
  assign n225 = ~n211 & n224;
  assign n226 = ~n210 & n225;
  assign n227 = ~n209 & n226;
  assign n228 = ~n208 & n227;
  assign n229 = ~n207 & n228;
  assign n230 = ~n206 & n229;
  assign n231 = ~n205 & n230;
  assign n232 = ~n204 & n231;
  assign \V138(1)  = ~n203 & n232;
  assign n234 = ~\V28(13)  & ~\V56(13) ;
  assign n235 = ~\V28(12)  & ~\V56(12) ;
  assign n236 = ~\V28(10)  & ~\V56(10) ;
  assign n237 = ~\V28(11)  & ~\V56(11) ;
  assign n238 = ~\V56(9)  & ~\V28(9) ;
  assign n239 = ~\V56(7)  & ~\V28(7) ;
  assign n240 = ~\V56(6)  & ~\V28(6) ;
  assign n241 = ~\V56(8)  & ~\V28(8) ;
  assign n242 = ~\V56(3)  & ~\V28(3) ;
  assign n243 = ~\V56(2)  & ~\V28(2) ;
  assign n244 = ~\V56(4)  & ~\V28(4) ;
  assign n245 = ~\V56(5)  & ~\V28(5) ;
  assign n246 = ~\V28(15)  & ~\V56(15) ;
  assign n247 = ~\V28(14)  & ~\V56(14) ;
  assign n248 = ~\V28(16)  & ~\V56(16) ;
  assign n249 = ~\V28(17)  & ~\V56(17) ;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n247 & n250;
  assign n252 = ~n246 & n251;
  assign n253 = ~n245 & n252;
  assign n254 = ~n244 & n253;
  assign n255 = ~n243 & n254;
  assign n256 = ~n242 & n255;
  assign n257 = ~n241 & n256;
  assign n258 = ~n240 & n257;
  assign n259 = ~n239 & n258;
  assign n260 = ~n238 & n259;
  assign n261 = ~n237 & n260;
  assign n262 = ~n236 & n261;
  assign n263 = ~n235 & n262;
  assign \V138(0)  = ~n234 & n263;
endmodule


