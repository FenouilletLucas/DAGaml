// Benchmark "TOP" written by ABC on Sun Apr 24 20:32:57 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
    n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342;
  assign n23 = i_5_ & ~i_9_;
  assign n24 = ~i_5_ & ~i_10_;
  assign n25 = i_0_ & ~n24;
  assign n26 = ~n23 & n25;
  assign n27 = i_6_ & i_9_;
  assign n28 = ~i_6_ & i_10_;
  assign n29 = ~n27 & ~n28;
  assign n30 = i_1_ & ~n29;
  assign n31 = ~n26 & ~n30;
  assign n32 = i_8_ & ~i_9_;
  assign n33 = ~i_8_ & ~i_10_;
  assign n34 = i_3_ & ~n33;
  assign n35 = ~n32 & n34;
  assign n36 = ~i_7_ & ~i_10_;
  assign n37 = i_7_ & ~i_9_;
  assign n38 = ~n36 & ~n37;
  assign n39 = i_2_ & n38;
  assign n40 = ~n35 & ~n39;
  assign o_0_ = ~n31 | ~n40;
  assign n42 = i_4_ & ~i_13_;
  assign n43 = ~i_8_ & i_11_;
  assign n44 = i_8_ & i_12_;
  assign n45 = ~i_3_ & ~n44;
  assign n46 = ~n43 & n45;
  assign n47 = ~n35 & ~n46;
  assign n48 = ~n42 & n47;
  assign n49 = n42 & ~n47;
  assign o_1_ = ~n48 & ~n49;
  assign n51 = i_0_ & i_2_;
  assign n52 = i_1_ & n51;
  assign n53 = ~n46 & n52;
  assign n54 = ~n38 & ~n53;
  assign n55 = ~i_1_ & ~i_6_;
  assign n56 = i_6_ & n51;
  assign n57 = i_2_ & i_5_;
  assign n58 = ~n56 & ~n57;
  assign n59 = i_12_ & ~n58;
  assign n60 = ~n55 & n59;
  assign n61 = ~i_5_ & ~i_6_;
  assign n62 = i_1_ & ~i_5_;
  assign n63 = i_0_ & ~i_6_;
  assign n64 = ~n62 & ~n63;
  assign n65 = ~n61 & n64;
  assign n66 = i_2_ & ~n65;
  assign n67 = i_11_ & n66;
  assign n68 = ~n60 & ~n67;
  assign n69 = ~n52 & n68;
  assign n70 = ~n54 & ~n69;
  assign n71 = ~i_7_ & n43;
  assign n72 = n61 & n71;
  assign n73 = ~n70 & ~n72;
  assign n74 = ~i_7_ & ~n64;
  assign n75 = i_0_ & i_1_;
  assign n76 = ~i_7_ & n75;
  assign n77 = ~n66 & ~n76;
  assign n78 = ~n74 & n77;
  assign n79 = ~i_8_ & ~n78;
  assign n80 = i_7_ & ~n66;
  assign n81 = n65 & ~n75;
  assign n82 = i_3_ & ~n81;
  assign n83 = ~n80 & n82;
  assign n84 = ~n79 & ~n83;
  assign n85 = i_11_ & ~n84;
  assign n86 = i_7_ & i_8_;
  assign n87 = i_5_ & n86;
  assign n88 = i_6_ & n87;
  assign n89 = i_3_ & i_6_;
  assign n90 = n57 & n89;
  assign n91 = ~i_11_ & ~n90;
  assign n92 = ~n88 & n91;
  assign n93 = i_8_ & ~n55;
  assign n94 = ~n58 & n93;
  assign n95 = i_3_ & i_7_;
  assign n96 = ~i_0_ & ~i_1_;
  assign n97 = n86 & ~n96;
  assign n98 = ~n95 & ~n97;
  assign n99 = ~i_0_ & ~i_5_;
  assign n100 = ~n55 & ~n99;
  assign n101 = ~n98 & n100;
  assign n102 = ~n94 & ~n101;
  assign n103 = i_3_ & n56;
  assign n104 = i_1_ & i_2_;
  assign n105 = i_5_ & n104;
  assign n106 = i_3_ & n105;
  assign n107 = ~n103 & ~n106;
  assign n108 = n102 & n107;
  assign n109 = n92 & n108;
  assign n110 = i_12_ & ~n109;
  assign n111 = i_5_ & i_12_;
  assign n112 = ~i_5_ & i_11_;
  assign n113 = ~n111 & ~n112;
  assign n114 = ~i_0_ & n113;
  assign n115 = ~n31 & ~n114;
  assign n116 = ~n110 & ~n115;
  assign n117 = ~n85 & n116;
  assign o_2_ = ~n73 | ~n117;
  assign n119 = i_1_ & i_6_;
  assign n120 = i_0_ & i_5_;
  assign n121 = ~i_3_ & ~n120;
  assign n122 = ~n119 & n121;
  assign n123 = ~i_7_ & n122;
  assign n124 = ~i_1_ & ~i_3_;
  assign n125 = ~i_2_ & ~i_5_;
  assign n126 = n124 & n125;
  assign n127 = ~n123 & ~n126;
  assign n128 = n33 & ~n127;
  assign n129 = ~i_6_ & ~i_8_;
  assign n130 = ~i_10_ & n129;
  assign n131 = ~i_2_ & ~i_3_;
  assign n132 = ~n120 & n131;
  assign n133 = n130 & n132;
  assign n134 = ~n23 & ~n99;
  assign n135 = ~n100 & ~n134;
  assign n136 = ~n133 & ~n135;
  assign n137 = ~i_1_ & ~i_2_;
  assign n138 = ~i_0_ & n137;
  assign n139 = ~i_3_ & ~i_8_;
  assign n140 = i_7_ & ~n139;
  assign n141 = n138 & ~n140;
  assign n142 = ~i_8_ & n37;
  assign n143 = i_1_ & ~i_6_;
  assign n144 = i_0_ & ~i_5_;
  assign n145 = ~i_3_ & ~n144;
  assign n146 = ~n143 & n145;
  assign n147 = n142 & n146;
  assign n148 = ~n141 & ~n147;
  assign n149 = n136 & n148;
  assign n150 = ~n128 & n149;
  assign n151 = ~i_11_ & ~n150;
  assign n152 = i_5_ & i_6_;
  assign n153 = ~i_3_ & i_4_;
  assign n154 = n37 & n153;
  assign n155 = n152 & n154;
  assign n156 = ~i_9_ & n152;
  assign n157 = ~i_2_ & n153;
  assign n158 = n156 & n157;
  assign n159 = ~i_1_ & n153;
  assign n160 = i_5_ & n37;
  assign n161 = n159 & n160;
  assign n162 = ~n158 & ~n161;
  assign n163 = ~i_2_ & i_5_;
  assign n164 = i_4_ & ~i_9_;
  assign n165 = i_3_ & ~i_8_;
  assign n166 = n164 & ~n165;
  assign n167 = n163 & n166;
  assign n168 = ~i_1_ & n167;
  assign n169 = n162 & ~n168;
  assign n170 = ~n155 & n169;
  assign n171 = i_4_ & n33;
  assign n172 = n137 & n171;
  assign n173 = ~n119 & n153;
  assign n174 = n36 & n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = ~i_5_ & ~n175;
  assign n177 = n170 & ~n176;
  assign n178 = ~i_6_ & ~i_7_;
  assign n179 = n171 & n178;
  assign n180 = ~i_2_ & ~i_6_;
  assign n181 = ~i_1_ & ~i_7_;
  assign n182 = ~n180 & ~n181;
  assign n183 = n171 & ~n182;
  assign n184 = ~i_2_ & ~i_10_;
  assign n185 = n173 & n184;
  assign n186 = ~n183 & ~n185;
  assign n187 = ~n179 & n186;
  assign n188 = ~i_5_ & ~n187;
  assign n189 = n177 & ~n188;
  assign n190 = ~n151 & n189;
  assign n191 = ~i_2_ & i_6_;
  assign n192 = ~i_0_ & ~i_3_;
  assign n193 = n164 & n192;
  assign n194 = n191 & n193;
  assign n195 = i_8_ & n164;
  assign n196 = n137 & n195;
  assign n197 = i_6_ & n37;
  assign n198 = ~i_6_ & n36;
  assign n199 = ~n197 & ~n198;
  assign n200 = n153 & ~n199;
  assign n201 = ~i_2_ & i_4_;
  assign n202 = i_6_ & n32;
  assign n203 = ~n130 & ~n202;
  assign n204 = n201 & ~n203;
  assign n205 = ~n200 & ~n204;
  assign n206 = ~n196 & n205;
  assign n207 = ~i_7_ & i_8_;
  assign n208 = i_4_ & n36;
  assign n209 = ~n195 & ~n208;
  assign n210 = ~n207 & ~n209;
  assign n211 = ~n154 & ~n210;
  assign n212 = ~i_1_ & ~n211;
  assign n213 = n206 & ~n212;
  assign n214 = ~i_0_ & ~n213;
  assign n215 = ~n194 & ~n214;
  assign n216 = n33 & n138;
  assign n217 = ~i_10_ & n192;
  assign n218 = ~n182 & n217;
  assign n219 = ~n216 & ~n218;
  assign n220 = i_4_ & ~n219;
  assign n221 = n215 & ~n220;
  assign n222 = i_7_ & ~i_12_;
  assign n223 = ~i_7_ & ~i_11_;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~i_10_ & ~n224;
  assign n226 = n180 & n225;
  assign n227 = i_6_ & i_7_;
  assign n228 = n195 & n227;
  assign n229 = ~n226 & ~n228;
  assign n230 = ~i_9_ & ~i_11_;
  assign n231 = ~i_7_ & n230;
  assign n232 = ~i_12_ & n37;
  assign n233 = ~n231 & ~n232;
  assign n234 = n191 & ~n233;
  assign n235 = ~n179 & ~n234;
  assign n236 = n229 & n235;
  assign n237 = ~i_0_ & ~n236;
  assign n238 = n184 & ~n233;
  assign n239 = ~i_10_ & n164;
  assign n240 = ~n238 & ~n239;
  assign n241 = ~n237 & n240;
  assign n242 = n96 & n131;
  assign n243 = i_7_ & ~n143;
  assign n244 = ~n191 & ~n243;
  assign n245 = n32 & ~n244;
  assign n246 = i_5_ & n245;
  assign n247 = ~n242 & ~n246;
  assign n248 = i_4_ & ~n247;
  assign n249 = ~n143 & n163;
  assign n250 = ~n233 & n249;
  assign n251 = i_6_ & ~i_12_;
  assign n252 = ~i_6_ & ~i_11_;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n25 & ~n253;
  assign n255 = ~i_1_ & n254;
  assign n256 = ~n250 & ~n255;
  assign n257 = ~n119 & n125;
  assign n258 = n225 & n257;
  assign n259 = ~i_9_ & ~i_10_;
  assign n260 = n46 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = n256 & n261;
  assign n263 = ~n248 & n262;
  assign n264 = n241 & n263;
  assign n265 = ~i_10_ & n207;
  assign n266 = n122 & n265;
  assign n267 = ~i_3_ & n137;
  assign n268 = n32 & n267;
  assign n269 = i_0_ & ~n268;
  assign n270 = i_5_ & ~n269;
  assign n271 = ~i_3_ & i_8_;
  assign n272 = ~i_7_ & ~n271;
  assign n273 = n138 & ~n272;
  assign n274 = ~n270 & ~n273;
  assign n275 = n145 & n245;
  assign n276 = ~i_1_ & i_6_;
  assign n277 = n23 & n276;
  assign n278 = ~n275 & ~n277;
  assign n279 = n274 & n278;
  assign n280 = ~n266 & n279;
  assign n281 = ~i_12_ & ~n280;
  assign n282 = n264 & ~n281;
  assign n283 = n221 & n282;
  assign o_3_ = ~n190 | ~n283;
  assign n285 = ~i_12_ & ~i_13_;
  assign n286 = n202 & n285;
  assign n287 = i_7_ & n286;
  assign n288 = ~i_9_ & ~i_13_;
  assign n289 = ~i_11_ & n288;
  assign n290 = ~i_8_ & n227;
  assign n291 = n289 & n290;
  assign n292 = ~n287 & ~n291;
  assign n293 = ~i_3_ & ~n292;
  assign n294 = n55 & n289;
  assign n295 = ~i_13_ & n164;
  assign n296 = i_6_ & n86;
  assign n297 = n295 & n296;
  assign n298 = ~n294 & ~n297;
  assign n299 = i_1_ & i_9_;
  assign n300 = i_6_ & n299;
  assign n301 = n37 & n191;
  assign n302 = n285 & n301;
  assign n303 = ~n300 & ~n302;
  assign n304 = i_9_ & i_12_;
  assign n305 = ~n153 & n304;
  assign n306 = n296 & n305;
  assign n307 = i_5_ & ~i_13_;
  assign n308 = ~n23 & ~n307;
  assign n309 = ~n306 & ~n308;
  assign n310 = n303 & n309;
  assign n311 = n298 & n310;
  assign n312 = i_2_ & i_7_;
  assign n313 = i_3_ & i_8_;
  assign n314 = i_4_ & ~n313;
  assign n315 = i_11_ & ~n314;
  assign n316 = ~n312 & ~n315;
  assign n317 = ~n252 & n304;
  assign n318 = ~n316 & n317;
  assign n319 = n311 & ~n318;
  assign n320 = ~n293 & n319;
  assign n321 = ~i_13_ & ~n44;
  assign n322 = n36 & n252;
  assign n323 = n321 & n322;
  assign n324 = ~i_3_ & n323;
  assign n325 = ~i_10_ & ~i_13_;
  assign n326 = n223 & n325;
  assign n327 = n180 & n326;
  assign n328 = i_4_ & n325;
  assign n329 = ~i_8_ & n178;
  assign n330 = n328 & n329;
  assign n331 = ~n327 & ~n330;
  assign n332 = i_10_ & i_11_;
  assign n333 = ~i_4_ & n332;
  assign n334 = ~i_12_ & ~n329;
  assign n335 = n333 & ~n334;
  assign n336 = ~i_11_ & ~i_13_;
  assign n337 = n55 & n336;
  assign n338 = n276 & n285;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~i_10_ & ~n339;
  assign n341 = ~i_5_ & ~i_13_;
  assign n342 = ~n143 & n341;
  assign n343 = ~n24 & ~n342;
  assign n344 = ~n340 & ~n343;
  assign n345 = ~n335 & n344;
  assign n346 = n331 & n345;
  assign n347 = ~n324 & n346;
  assign n348 = ~n320 & ~n347;
  assign n349 = ~n157 & n304;
  assign n350 = n332 & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = ~i_13_ & ~n240;
  assign n353 = i_8_ & n152;
  assign n354 = n295 & n353;
  assign n355 = ~i_13_ & n171;
  assign n356 = ~i_11_ & n325;
  assign n357 = ~i_12_ & n356;
  assign n358 = ~n355 & ~n357;
  assign n359 = n61 & ~n358;
  assign n360 = ~i_12_ & n288;
  assign n361 = n152 & n360;
  assign n362 = ~i_11_ & n361;
  assign n363 = ~n359 & ~n362;
  assign n364 = ~n354 & n363;
  assign n365 = ~i_2_ & ~n364;
  assign n366 = ~n43 & n321;
  assign n367 = n259 & n366;
  assign n368 = ~i_3_ & ~n367;
  assign n369 = i_7_ & i_9_;
  assign n370 = i_10_ & i_12_;
  assign n371 = n369 & n370;
  assign n372 = i_6_ & n371;
  assign n373 = ~i_7_ & n332;
  assign n374 = i_9_ & n373;
  assign n375 = i_3_ & ~n374;
  assign n376 = ~n89 & ~n375;
  assign n377 = ~n372 & ~n376;
  assign n378 = ~n368 & ~n377;
  assign n379 = n23 & n86;
  assign n380 = n42 & n379;
  assign n381 = ~i_7_ & ~i_8_;
  assign n382 = ~i_5_ & n381;
  assign n383 = n328 & n382;
  assign n384 = ~n380 & ~n383;
  assign n385 = ~n361 & n384;
  assign n386 = ~i_1_ & ~n385;
  assign n387 = i_9_ & i_10_;
  assign n388 = i_1_ & n387;
  assign n389 = i_0_ & ~n388;
  assign n390 = i_7_ & n152;
  assign n391 = n288 & n390;
  assign n392 = n198 & n341;
  assign n393 = ~n391 & ~n392;
  assign n394 = n153 & ~n393;
  assign n395 = n389 & ~n394;
  assign n396 = ~n386 & n395;
  assign n397 = ~n378 & n396;
  assign n398 = ~n365 & n397;
  assign n399 = ~n352 & n398;
  assign n400 = n351 & n399;
  assign n401 = ~i_11_ & i_12_;
  assign n402 = ~i_4_ & n401;
  assign n403 = i_2_ & i_8_;
  assign n404 = ~n95 & ~n403;
  assign n405 = i_1_ & ~n404;
  assign n406 = n402 & n405;
  assign n407 = ~n296 & ~n406;
  assign n408 = ~i_11_ & n304;
  assign n409 = i_3_ & n408;
  assign n410 = i_11_ & ~i_12_;
  assign n411 = ~i_13_ & n410;
  assign n412 = ~i_3_ & n411;
  assign n413 = i_11_ & n295;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~i_9_ & ~n414;
  assign n416 = ~n409 & ~n415;
  assign n417 = ~n402 & n416;
  assign n418 = ~n407 & ~n417;
  assign n419 = ~n276 & ~n301;
  assign n420 = n411 & ~n419;
  assign n421 = i_6_ & n312;
  assign n422 = n408 & n421;
  assign n423 = ~i_11_ & i_13_;
  assign n424 = ~n422 & ~n423;
  assign n425 = ~i_11_ & n300;
  assign n426 = n424 & ~n425;
  assign n427 = ~n420 & n426;
  assign n428 = ~n418 & n427;
  assign n429 = ~i_5_ & ~n428;
  assign n430 = ~i_4_ & n410;
  assign n431 = i_3_ & ~i_12_;
  assign n432 = n332 & n431;
  assign n433 = ~n430 & ~n432;
  assign n434 = i_1_ & n433;
  assign n435 = n57 & n129;
  assign n436 = i_3_ & i_5_;
  assign n437 = n178 & n436;
  assign n438 = ~n435 & ~n437;
  assign n439 = n430 & ~n438;
  assign n440 = i_12_ & n325;
  assign n441 = ~i_3_ & ~i_11_;
  assign n442 = ~i_4_ & ~n441;
  assign n443 = n440 & ~n442;
  assign n444 = ~i_1_ & ~n443;
  assign n445 = n381 & ~n444;
  assign n446 = i_5_ & n445;
  assign n447 = ~n439 & ~n446;
  assign n448 = ~n434 & ~n447;
  assign n449 = ~i_5_ & i_6_;
  assign n450 = ~n404 & n449;
  assign n451 = n62 & n86;
  assign n452 = ~n450 & ~n451;
  assign n453 = n402 & ~n452;
  assign n454 = ~n448 & ~n453;
  assign n455 = ~n429 & n454;
  assign n456 = ~i_0_ & n455;
  assign n457 = ~n400 & ~n456;
  assign n458 = n51 & ~n153;
  assign n459 = n304 & n353;
  assign n460 = n458 & n459;
  assign n461 = ~i_8_ & i_10_;
  assign n462 = i_3_ & n461;
  assign n463 = i_12_ & n462;
  assign n464 = n144 & n463;
  assign n465 = i_11_ & n464;
  assign n466 = ~n460 & ~n465;
  assign n467 = n144 & ~n251;
  assign n468 = n373 & n467;
  assign n469 = i_2_ & n468;
  assign n470 = n466 & ~n469;
  assign n471 = i_8_ & i_9_;
  assign n472 = ~i_7_ & n471;
  assign n473 = n436 & n472;
  assign n474 = ~i_4_ & i_5_;
  assign n475 = i_2_ & i_3_;
  assign n476 = ~i_0_ & n475;
  assign n477 = i_9_ & n381;
  assign n478 = ~n476 & ~n477;
  assign n479 = n474 & ~n478;
  assign n480 = ~n473 & ~n479;
  assign n481 = ~i_6_ & i_11_;
  assign n482 = ~i_12_ & n481;
  assign n483 = ~n480 & n482;
  assign n484 = i_0_ & n137;
  assign n485 = n232 & n307;
  assign n486 = ~n153 & ~n223;
  assign n487 = ~i_5_ & n325;
  assign n488 = ~n486 & n487;
  assign n489 = ~i_3_ & i_5_;
  assign n490 = n295 & n489;
  assign n491 = ~n488 & ~n490;
  assign n492 = ~n485 & n491;
  assign n493 = n484 & ~n492;
  assign n494 = ~n483 & ~n493;
  assign n495 = i_10_ & n86;
  assign n496 = ~n476 & ~n495;
  assign n497 = n402 & ~n496;
  assign n498 = n408 & n476;
  assign n499 = i_11_ & ~i_13_;
  assign n500 = ~i_9_ & n499;
  assign n501 = ~i_0_ & n201;
  assign n502 = n500 & n501;
  assign n503 = n288 & n410;
  assign n504 = ~i_0_ & n131;
  assign n505 = n503 & n504;
  assign n506 = ~n502 & ~n505;
  assign n507 = ~n498 & n506;
  assign n508 = i_8_ & ~n507;
  assign n509 = ~n497 & ~n508;
  assign n510 = n449 & ~n509;
  assign n511 = n75 & ~n153;
  assign n512 = n87 & n511;
  assign n513 = i_10_ & n56;
  assign n514 = ~n512 & ~n513;
  assign n515 = n304 & ~n514;
  assign n516 = n227 & n304;
  assign n517 = i_2_ & n299;
  assign n518 = ~n516 & ~n517;
  assign n519 = i_3_ & ~i_4_;
  assign n520 = n120 & n519;
  assign n521 = ~n518 & n520;
  assign n522 = i_2_ & n63;
  assign n523 = i_11_ & n387;
  assign n524 = n522 & n523;
  assign n525 = ~n521 & ~n524;
  assign n526 = ~n515 & n525;
  assign n527 = ~n510 & n526;
  assign n528 = n494 & n527;
  assign n529 = n470 & n528;
  assign n530 = ~n457 & n529;
  assign n531 = i_2_ & i_10_;
  assign n532 = i_6_ & ~i_7_;
  assign n533 = n401 & n532;
  assign n534 = n75 & n165;
  assign n535 = ~n76 & ~n534;
  assign n536 = ~n533 & n535;
  assign n537 = n531 & ~n536;
  assign n538 = n139 & n356;
  assign n539 = ~n355 & ~n538;
  assign n540 = n484 & ~n539;
  assign n541 = ~n76 & ~n522;
  assign n542 = i_3_ & n333;
  assign n543 = ~n541 & n542;
  assign n544 = ~i_7_ & ~n313;
  assign n545 = ~i_0_ & n104;
  assign n546 = ~i_11_ & n545;
  assign n547 = i_9_ & n546;
  assign n548 = ~n544 & n547;
  assign n549 = ~n543 & ~n548;
  assign n550 = ~n540 & n549;
  assign n551 = ~n191 & ~n227;
  assign n552 = n193 & ~n551;
  assign n553 = n187 & ~n552;
  assign n554 = n499 & ~n553;
  assign n555 = n159 & n500;
  assign n556 = ~i_0_ & n555;
  assign n557 = n138 & n411;
  assign n558 = ~n556 & ~n557;
  assign n559 = i_7_ & ~n558;
  assign n560 = ~i_10_ & n285;
  assign n561 = i_8_ & n560;
  assign n562 = ~n328 & ~n561;
  assign n563 = i_0_ & n131;
  assign n564 = ~n562 & n563;
  assign n565 = ~i_6_ & n564;
  assign n566 = ~n559 & ~n565;
  assign n567 = ~n554 & n566;
  assign n568 = n550 & n567;
  assign n569 = ~n537 & n568;
  assign n570 = i_2_ & ~i_8_;
  assign n571 = i_10_ & ~i_11_;
  assign n572 = i_3_ & n571;
  assign n573 = n570 & n572;
  assign n574 = ~i_6_ & n571;
  assign n575 = ~n573 & ~n574;
  assign n576 = i_1_ & ~n575;
  assign n577 = ~i_2_ & i_8_;
  assign n578 = ~n414 & n577;
  assign n579 = n96 & n578;
  assign n580 = ~i_5_ & ~n579;
  assign n581 = ~n576 & n580;
  assign n582 = n259 & n411;
  assign n583 = n271 & n582;
  assign n584 = n42 & n259;
  assign n585 = i_11_ & n584;
  assign n586 = ~n583 & ~n585;
  assign n587 = i_0_ & n124;
  assign n588 = ~i_7_ & ~n562;
  assign n589 = n587 & n588;
  assign n590 = ~i_8_ & n104;
  assign n591 = n333 & n590;
  assign n592 = i_0_ & n591;
  assign n593 = ~n589 & ~n592;
  assign n594 = n586 & n593;
  assign n595 = n581 & n594;
  assign n596 = n265 & n412;
  assign n597 = n184 & n499;
  assign n598 = n222 & n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = ~n119 & ~n599;
  assign n601 = ~i_0_ & i_1_;
  assign n602 = n409 & n601;
  assign n603 = n96 & n415;
  assign n604 = ~n602 & ~n603;
  assign n605 = n86 & ~n604;
  assign n606 = ~n600 & ~n605;
  assign n607 = ~i_5_ & ~n606;
  assign n608 = n595 & ~n607;
  assign n609 = n569 & n608;
  assign n610 = i_4_ & n440;
  assign n611 = n192 & n610;
  assign n612 = i_2_ & ~i_12_;
  assign n613 = n332 & n612;
  assign n614 = ~i_0_ & n613;
  assign n615 = ~n611 & ~n614;
  assign n616 = ~i_6_ & ~n615;
  assign n617 = n410 & n519;
  assign n618 = ~i_12_ & n531;
  assign n619 = ~n617 & ~n618;
  assign n620 = n601 & ~n619;
  assign n621 = i_12_ & ~i_13_;
  assign n622 = ~i_11_ & n621;
  assign n623 = n138 & n622;
  assign n624 = ~n620 & ~n623;
  assign n625 = ~n616 & n624;
  assign n626 = ~i_7_ & ~n625;
  assign n627 = ~i_12_ & n545;
  assign n628 = n43 & n627;
  assign n629 = n75 & ~n404;
  assign n630 = ~n103 & ~n629;
  assign n631 = n304 & ~n630;
  assign n632 = ~n628 & ~n631;
  assign n633 = ~i_4_ & ~n632;
  assign n634 = ~n626 & ~n633;
  assign n635 = n219 & ~n245;
  assign n636 = n621 & ~n635;
  assign n637 = i_8_ & n484;
  assign n638 = n288 & n637;
  assign n639 = ~n636 & ~n638;
  assign n640 = i_4_ & ~n639;
  assign n641 = n440 & n501;
  assign n642 = ~i_12_ & n332;
  assign n643 = n476 & n642;
  assign n644 = i_12_ & n356;
  assign n645 = n504 & n644;
  assign n646 = ~n643 & ~n645;
  assign n647 = ~n641 & n646;
  assign n648 = n129 & ~n647;
  assign n649 = n139 & n622;
  assign n650 = ~n138 & ~n259;
  assign n651 = n649 & ~n650;
  assign n652 = n369 & n612;
  assign n653 = n481 & n652;
  assign n654 = n37 & n42;
  assign n655 = n587 & n654;
  assign n656 = ~n653 & ~n655;
  assign n657 = i_5_ & n656;
  assign n658 = ~n651 & n657;
  assign n659 = ~n648 & n658;
  assign n660 = ~n640 & n659;
  assign n661 = n433 & ~n443;
  assign n662 = n329 & ~n661;
  assign n663 = i_12_ & ~n337;
  assign n664 = ~n327 & n663;
  assign n665 = ~n285 & ~n664;
  assign n666 = ~n662 & ~n665;
  assign n667 = ~i_0_ & ~n666;
  assign n668 = n51 & ~n544;
  assign n669 = ~n251 & ~n668;
  assign n670 = n299 & ~n669;
  assign n671 = i_10_ & ~i_12_;
  assign n672 = n165 & n545;
  assign n673 = ~i_0_ & n143;
  assign n674 = ~n672 & ~n673;
  assign n675 = n671 & ~n674;
  assign n676 = ~n670 & ~n675;
  assign n677 = i_6_ & n295;
  assign n678 = n563 & n677;
  assign n679 = n139 & n289;
  assign n680 = n271 & n360;
  assign n681 = ~n679 & ~n680;
  assign n682 = n484 & ~n681;
  assign n683 = ~n678 & ~n682;
  assign n684 = n676 & n683;
  assign n685 = ~n667 & n684;
  assign n686 = n660 & n685;
  assign n687 = n634 & n686;
  assign n688 = ~n609 & ~n687;
  assign n689 = n142 & n336;
  assign n690 = n489 & n689;
  assign n691 = ~n143 & n690;
  assign n692 = i_12_ & n691;
  assign n693 = n231 & n249;
  assign n694 = n170 & ~n693;
  assign n695 = n621 & ~n694;
  assign n696 = ~n692 & ~n695;
  assign n697 = ~i_5_ & n519;
  assign n698 = n75 & n531;
  assign n699 = ~n546 & ~n698;
  assign n700 = n697 & ~n699;
  assign n701 = n87 & n587;
  assign n702 = n353 & n563;
  assign n703 = ~n701 & ~n702;
  assign n704 = n360 & ~n703;
  assign n705 = ~n700 & ~n704;
  assign n706 = ~i_5_ & n153;
  assign n707 = n499 & n706;
  assign n708 = i_5_ & n153;
  assign n709 = n621 & n708;
  assign n710 = ~n707 & ~n709;
  assign n711 = n138 & ~n710;
  assign n712 = n111 & n584;
  assign n713 = i_3_ & n449;
  assign n714 = i_7_ & n461;
  assign n715 = n713 & n714;
  assign n716 = n401 & n715;
  assign n717 = ~n712 & ~n716;
  assign n718 = ~n711 & n717;
  assign n719 = n705 & n718;
  assign n720 = i_5_ & n519;
  assign n721 = i_9_ & n313;
  assign n722 = ~n38 & ~n721;
  assign n723 = ~i_11_ & ~n722;
  assign n724 = ~n720 & ~n723;
  assign n725 = n627 & ~n724;
  assign n726 = ~n165 & ~n519;
  assign n727 = n144 & n178;
  assign n728 = ~n726 & n727;
  assign n729 = n382 & n511;
  assign n730 = ~i_8_ & n61;
  assign n731 = n458 & n730;
  assign n732 = ~n729 & ~n731;
  assign n733 = ~n728 & n732;
  assign n734 = n332 & ~n733;
  assign n735 = n563 & n730;
  assign n736 = n382 & n587;
  assign n737 = ~n735 & ~n736;
  assign n738 = n356 & ~n737;
  assign n739 = ~n734 & ~n738;
  assign n740 = ~n725 & n739;
  assign n741 = n719 & n740;
  assign n742 = n696 & n741;
  assign n743 = i_12_ & n499;
  assign n744 = ~n221 & n743;
  assign n745 = n742 & ~n744;
  assign n746 = ~n688 & n745;
  assign o_4_ = ~n530 | ~n746;
  assign n748 = i_3_ & n143;
  assign n749 = i_10_ & n381;
  assign n750 = n748 & n749;
  assign n751 = ~n38 & n159;
  assign n752 = ~n196 & ~n751;
  assign n753 = n621 & ~n752;
  assign n754 = ~i_3_ & ~i_6_;
  assign n755 = ~n312 & n754;
  assign n756 = n561 & n755;
  assign n757 = ~n753 & ~n756;
  assign n758 = ~n750 & n757;
  assign n759 = i_11_ & ~n758;
  assign n760 = ~i_11_ & n369;
  assign n761 = i_2_ & n760;
  assign n762 = i_2_ & ~n32;
  assign n763 = n411 & ~n475;
  assign n764 = ~n762 & n763;
  assign n765 = ~n519 & ~n721;
  assign n766 = n401 & ~n765;
  assign n767 = i_8_ & n413;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n764 & n768;
  assign n770 = i_7_ & ~n769;
  assign n771 = ~n423 & ~n770;
  assign n772 = ~n761 & n771;
  assign n773 = ~i_6_ & ~n772;
  assign n774 = ~i_2_ & ~i_7_;
  assign n775 = n44 & ~n774;
  assign n776 = ~i_4_ & n252;
  assign n777 = n775 & n776;
  assign n778 = n532 & ~n619;
  assign n779 = ~n777 & ~n778;
  assign n780 = n381 & ~n661;
  assign n781 = ~i_12_ & i_13_;
  assign n782 = n622 & n774;
  assign n783 = n430 & n570;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~n781 & n784;
  assign n786 = ~n780 & n785;
  assign n787 = i_6_ & ~n786;
  assign n788 = ~i_1_ & ~n787;
  assign n789 = n779 & n788;
  assign n790 = ~n773 & n789;
  assign n791 = n205 & n240;
  assign n792 = n236 & n791;
  assign n793 = ~i_13_ & ~n792;
  assign n794 = i_6_ & i_11_;
  assign n795 = n472 & n794;
  assign n796 = n375 & ~n795;
  assign n797 = ~n371 & n796;
  assign n798 = ~n287 & ~n323;
  assign n799 = i_6_ & n689;
  assign n800 = n798 & ~n799;
  assign n801 = n368 & n800;
  assign n802 = ~n797 & ~n801;
  assign n803 = ~i_13_ & ~n71;
  assign n804 = ~n29 & ~n42;
  assign n805 = ~n803 & n804;
  assign n806 = n304 & n794;
  assign n807 = n370 & n481;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~i_4_ & ~n808;
  assign n810 = ~i_9_ & ~n178;
  assign n811 = ~n421 & ~n531;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n809 & ~n812;
  assign n814 = i_1_ & ~n306;
  assign n815 = n813 & n814;
  assign n816 = ~n805 & n815;
  assign n817 = ~n802 & n816;
  assign n818 = ~n793 & n817;
  assign n819 = ~n790 & ~n818;
  assign n820 = n104 & n462;
  assign n821 = ~i_6_ & ~n591;
  assign n822 = ~n820 & n821;
  assign n823 = ~i_1_ & n475;
  assign n824 = ~i_11_ & n471;
  assign n825 = n823 & n824;
  assign n826 = i_1_ & n519;
  assign n827 = n373 & n826;
  assign n828 = ~n825 & ~n827;
  assign n829 = ~n573 & n828;
  assign n830 = n822 & n829;
  assign n831 = n586 & n830;
  assign n832 = n157 & n499;
  assign n833 = ~n578 & ~n832;
  assign n834 = ~i_1_ & ~n833;
  assign n835 = ~i_11_ & n463;
  assign n836 = ~n555 & ~n835;
  assign n837 = i_7_ & ~n836;
  assign n838 = i_1_ & n131;
  assign n839 = n43 & ~n312;
  assign n840 = ~n838 & ~n839;
  assign n841 = n328 & ~n840;
  assign n842 = ~n837 & ~n841;
  assign n843 = ~n834 & n842;
  assign n844 = n831 & n843;
  assign n845 = ~n312 & ~n531;
  assign n846 = n159 & n845;
  assign n847 = ~n239 & ~n846;
  assign n848 = ~n172 & n847;
  assign n849 = n621 & ~n848;
  assign n850 = ~n104 & ~n612;
  assign n851 = n721 & ~n850;
  assign n852 = i_6_ & ~n652;
  assign n853 = ~n851 & n852;
  assign n854 = n37 & n649;
  assign n855 = n44 & n654;
  assign n856 = n671 & n823;
  assign n857 = n267 & n622;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~i_8_ & ~n858;
  assign n860 = ~n855 & ~n859;
  assign n861 = ~n854 & n860;
  assign n862 = n853 & n861;
  assign n863 = ~n849 & n862;
  assign n864 = ~n844 & ~n863;
  assign n865 = n574 & n775;
  assign n866 = i_2_ & ~n45;
  assign n867 = n30 & n866;
  assign n868 = ~n253 & n823;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n865 & n869;
  assign n871 = ~i_4_ & ~n870;
  assign n872 = n130 & n336;
  assign n873 = ~n286 & ~n872;
  assign n874 = ~n677 & n873;
  assign n875 = n838 & ~n874;
  assign n876 = n516 & n826;
  assign n877 = n714 & n748;
  assign n878 = i_12_ & n877;
  assign n879 = ~n876 & ~n878;
  assign n880 = n431 & n795;
  assign n881 = ~n37 & n574;
  assign n882 = i_2_ & n881;
  assign n883 = ~n880 & ~n882;
  assign n884 = n879 & n883;
  assign n885 = ~n875 & n884;
  assign n886 = ~n871 & n885;
  assign n887 = ~n864 & n886;
  assign n888 = ~n819 & n887;
  assign o_5_ = n759 | ~n888;
  assign n890 = ~n430 & ~n610;
  assign n891 = ~i_8_ & ~n890;
  assign n892 = ~i_13_ & ~n519;
  assign n893 = ~i_12_ & ~n892;
  assign n894 = ~n649 & ~n893;
  assign n895 = ~n891 & n894;
  assign n896 = ~i_2_ & ~n895;
  assign n897 = n42 & n475;
  assign n898 = i_8_ & n897;
  assign n899 = ~n157 & ~n195;
  assign n900 = n621 & ~n899;
  assign n901 = ~n898 & ~n900;
  assign n902 = i_7_ & n901;
  assign n903 = ~n896 & n902;
  assign n904 = ~n195 & n572;
  assign n905 = ~i_8_ & n897;
  assign n906 = ~i_2_ & ~i_11_;
  assign n907 = ~n721 & n892;
  assign n908 = n906 & ~n907;
  assign n909 = ~n905 & ~n908;
  assign n910 = ~n904 & n909;
  assign n911 = i_11_ & ~n471;
  assign n912 = n328 & n911;
  assign n913 = n402 & n577;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~i_7_ & n914;
  assign n916 = n910 & n915;
  assign n917 = n833 & n916;
  assign n918 = ~n903 & ~n917;
  assign n919 = i_9_ & n86;
  assign n920 = ~i_2_ & n714;
  assign n921 = ~n919 & ~n920;
  assign n922 = n431 & ~n921;
  assign n923 = ~n918 & ~n922;
  assign n924 = ~n588 & ~n654;
  assign n925 = ~i_3_ & ~n924;
  assign n926 = i_7_ & ~n681;
  assign n927 = ~n584 & ~n926;
  assign n928 = i_3_ & n387;
  assign n929 = n230 & n560;
  assign n930 = ~i_3_ & n929;
  assign n931 = ~n928 & ~n930;
  assign n932 = n38 & ~n42;
  assign n933 = ~n366 & n932;
  assign n934 = ~i_7_ & n538;
  assign n935 = ~n933 & ~n934;
  assign n936 = n931 & n935;
  assign n937 = n927 & n936;
  assign n938 = ~n925 & n937;
  assign n939 = i_2_ & ~n938;
  assign n940 = n39 & n519;
  assign n941 = ~n939 & ~n940;
  assign o_6_ = ~n923 | ~n941;
  assign n943 = ~i_2_ & n75;
  assign n944 = i_6_ & n381;
  assign n945 = n413 & n489;
  assign n946 = n288 & n720;
  assign n947 = n571 & n946;
  assign n948 = ~n945 & ~n947;
  assign n949 = n944 & ~n948;
  assign n950 = i_3_ & n61;
  assign n951 = n714 & n781;
  assign n952 = n950 & n951;
  assign n953 = ~i_7_ & n423;
  assign n954 = n471 & n953;
  assign n955 = i_5_ & n89;
  assign n956 = n954 & n955;
  assign n957 = ~n952 & ~n956;
  assign n958 = i_6_ & n489;
  assign n959 = n423 & n477;
  assign n960 = n958 & n959;
  assign n961 = n671 & n720;
  assign n962 = n288 & n290;
  assign n963 = n961 & n962;
  assign n964 = ~n960 & ~n963;
  assign n965 = ~i_3_ & n61;
  assign n966 = n495 & n781;
  assign n967 = n965 & n966;
  assign n968 = n964 & ~n967;
  assign n969 = n957 & n968;
  assign n970 = ~n949 & n969;
  assign n971 = n943 & ~n970;
  assign n972 = n293 & n474;
  assign n973 = i_3_ & i_4_;
  assign n974 = n288 & n973;
  assign n975 = n88 & n974;
  assign n976 = n290 & n945;
  assign n977 = ~n975 & ~n976;
  assign n978 = i_10_ & n697;
  assign n979 = ~i_5_ & n973;
  assign n980 = n325 & n979;
  assign n981 = ~n978 & ~n980;
  assign n982 = n329 & ~n981;
  assign n983 = i_10_ & n781;
  assign n984 = n207 & n983;
  assign n985 = n965 & n984;
  assign n986 = n369 & n423;
  assign n987 = ~i_8_ & n986;
  assign n988 = n958 & n987;
  assign n989 = ~n985 & ~n988;
  assign n990 = ~n982 & n989;
  assign n991 = n977 & n990;
  assign n992 = n749 & n950;
  assign n993 = n919 & n955;
  assign n994 = ~n928 & ~n993;
  assign n995 = ~n992 & n994;
  assign n996 = i_13_ & ~n995;
  assign n997 = ~i_3_ & ~i_4_;
  assign n998 = ~i_5_ & n997;
  assign n999 = n323 & n998;
  assign n1000 = ~i_4_ & ~n931;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~n996 & n1001;
  assign n1003 = n991 & n1002;
  assign n1004 = ~n972 & n1003;
  assign n1005 = n52 & ~n1004;
  assign n1006 = ~n971 & ~n1005;
  assign n1007 = i_9_ & ~n72;
  assign n1008 = n75 & n475;
  assign n1009 = ~n71 & ~n1008;
  assign n1010 = ~n81 & ~n1009;
  assign n1011 = n325 & n1010;
  assign n1012 = ~n1007 & n1011;
  assign n1013 = i_3_ & n198;
  assign n1014 = i_2_ & n130;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = n500 & ~n1015;
  assign n1017 = ~n89 & ~n93;
  assign n1018 = n37 & ~n1017;
  assign n1019 = i_2_ & n202;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = n440 & ~n1020;
  assign n1022 = ~n1016 & ~n1021;
  assign n1023 = i_0_ & ~n1022;
  assign n1024 = n242 & n743;
  assign n1025 = ~n55 & n621;
  assign n1026 = ~n28 & n1025;
  assign n1027 = n379 & n1026;
  assign n1028 = ~n1024 & ~n1027;
  assign n1029 = ~n1023 & n1028;
  assign n1030 = ~n1012 & n1029;
  assign n1031 = i_4_ & ~n1030;
  assign n1032 = n1006 & ~n1031;
  assign n1033 = i_5_ & n754;
  assign n1034 = n984 & n1033;
  assign n1035 = n329 & n961;
  assign n1036 = n500 & n706;
  assign n1037 = n290 & n1036;
  assign n1038 = ~n1035 & ~n1037;
  assign n1039 = ~n165 & n449;
  assign n1040 = n986 & n1039;
  assign n1041 = ~n271 & n1040;
  assign n1042 = n381 & n983;
  assign n1043 = ~i_6_ & n436;
  assign n1044 = n1042 & n1043;
  assign n1045 = ~n1041 & ~n1044;
  assign n1046 = n1038 & n1045;
  assign n1047 = ~n1034 & n1046;
  assign n1048 = n545 & ~n1047;
  assign n1049 = n730 & n953;
  assign n1050 = i_10_ & n1049;
  assign n1051 = ~n1048 & ~n1050;
  assign n1052 = ~i_2_ & n601;
  assign n1053 = i_8_ & n532;
  assign n1054 = n1052 & n1053;
  assign n1055 = n296 & n545;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = i_2_ & n96;
  assign n1058 = ~i_6_ & n86;
  assign n1059 = n1057 & n1058;
  assign n1060 = n1056 & ~n1059;
  assign n1061 = n112 & n974;
  assign n1062 = ~n1060 & n1061;
  assign n1063 = i_5_ & n973;
  assign n1064 = ~i_4_ & n489;
  assign n1065 = ~i_12_ & n1064;
  assign n1066 = ~n1063 & ~n1065;
  assign n1067 = ~i_1_ & n51;
  assign n1068 = n1058 & n1067;
  assign n1069 = n943 & n1053;
  assign n1070 = n178 & n637;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1068 & n1071;
  assign n1073 = n500 & ~n1072;
  assign n1074 = ~n1066 & n1073;
  assign n1075 = ~n1062 & ~n1074;
  assign n1076 = n353 & n652;
  assign n1077 = n826 & n1076;
  assign n1078 = n1075 & ~n1077;
  assign n1079 = n1051 & n1078;
  assign n1080 = ~i_4_ & n271;
  assign n1081 = ~n541 & n1080;
  assign n1082 = n403 & n998;
  assign n1083 = ~n276 & n1082;
  assign n1084 = ~n1081 & ~n1083;
  assign n1085 = n582 & ~n1084;
  assign n1086 = i_7_ & n129;
  assign n1087 = n945 & n1086;
  assign n1088 = ~n253 & n946;
  assign n1089 = n713 & n781;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n749 & ~n1090;
  assign n1092 = n423 & n919;
  assign n1093 = n1043 & n1092;
  assign n1094 = n987 & n1033;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~i_3_ & n449;
  assign n1097 = n984 & n1096;
  assign n1098 = n1095 & ~n1097;
  assign n1099 = ~n1091 & n1098;
  assign n1100 = ~n1087 & n1099;
  assign n1101 = n1067 & ~n1100;
  assign n1102 = n944 & n1057;
  assign n1103 = n129 & n601;
  assign n1104 = ~n774 & n1103;
  assign n1105 = ~n312 & n1104;
  assign n1106 = ~n1102 & ~n1105;
  assign n1107 = n325 & ~n1106;
  assign n1108 = ~n962 & ~n1107;
  assign n1109 = n1064 & ~n1108;
  assign n1110 = n401 & n1109;
  assign n1111 = ~n1101 & ~n1110;
  assign n1112 = ~n1085 & n1111;
  assign n1113 = n1079 & n1112;
  assign n1114 = n499 & n671;
  assign n1115 = n697 & n1114;
  assign n1116 = n1086 & n1115;
  assign n1117 = n336 & n720;
  assign n1118 = n304 & n1117;
  assign n1119 = n1053 & n1118;
  assign n1120 = i_8_ & n178;
  assign n1121 = n411 & n998;
  assign n1122 = ~n1061 & ~n1121;
  assign n1123 = n1120 & ~n1122;
  assign n1124 = ~n1119 & ~n1123;
  assign n1125 = n296 & n709;
  assign n1126 = n950 & n954;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = n329 & n707;
  assign n1129 = n1127 & ~n1128;
  assign n1130 = n1124 & n1129;
  assign n1131 = n290 & n474;
  assign n1132 = n622 & n1131;
  assign n1133 = ~n1049 & ~n1132;
  assign n1134 = ~i_3_ & ~n1133;
  assign n1135 = ~n271 & ~n462;
  assign n1136 = n390 & ~n1135;
  assign n1137 = ~n441 & ~n1136;
  assign n1138 = n781 & ~n1137;
  assign n1139 = ~n1134 & ~n1138;
  assign n1140 = n1130 & n1139;
  assign n1141 = ~n1116 & n1140;
  assign n1142 = n138 & ~n1141;
  assign n1143 = n950 & n1092;
  assign n1144 = n571 & n621;
  assign n1145 = n720 & n1144;
  assign n1146 = n329 & n1145;
  assign n1147 = ~n1143 & ~n1146;
  assign n1148 = n944 & n1115;
  assign n1149 = n1147 & ~n1148;
  assign n1150 = n955 & n1042;
  assign n1151 = n1036 & n1086;
  assign n1152 = n965 & n987;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1150 & n1153;
  assign n1155 = n1058 & n1118;
  assign n1156 = n958 & n984;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = n1154 & n1157;
  assign n1159 = n1149 & n1158;
  assign n1160 = n1057 & ~n1159;
  assign n1161 = n966 & n1033;
  assign n1162 = n944 & n1036;
  assign n1163 = n951 & n1043;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = n959 & n1096;
  assign n1166 = n713 & n954;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = n1164 & n1167;
  assign n1169 = ~n1161 & n1168;
  assign n1170 = n1052 & ~n1169;
  assign n1171 = n329 & n945;
  assign n1172 = n959 & n1033;
  assign n1173 = n713 & n951;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n954 & n1043;
  assign n1176 = n966 & n1096;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = n1174 & n1177;
  assign n1179 = ~n1171 & n1178;
  assign n1180 = n484 & ~n1179;
  assign n1181 = ~n1170 & ~n1180;
  assign n1182 = ~n1160 & n1181;
  assign n1183 = ~n1142 & n1182;
  assign n1184 = ~n107 & n983;
  assign n1185 = n341 & n617;
  assign n1186 = n184 & n1058;
  assign n1187 = n1185 & n1186;
  assign n1188 = ~n1184 & ~n1187;
  assign n1189 = n52 & n296;
  assign n1190 = ~i_6_ & n1057;
  assign n1191 = n138 & n532;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = n1144 & ~n1192;
  assign n1194 = n644 & n1052;
  assign n1195 = n1120 & n1194;
  assign n1196 = ~n1193 & ~n1195;
  assign n1197 = ~n1189 & n1196;
  assign n1198 = n720 & ~n1197;
  assign n1199 = n531 & n826;
  assign n1200 = n113 & n1199;
  assign n1201 = ~n1198 & ~n1200;
  assign n1202 = n1188 & n1201;
  assign n1203 = i_13_ & n571;
  assign n1204 = i_3_ & n74;
  assign n1205 = n61 & n475;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n79 & n1206;
  assign n1208 = n1203 & ~n1207;
  assign n1209 = i_9_ & ~n1208;
  assign n1210 = n1202 & n1209;
  assign n1211 = i_7_ & n75;
  assign n1212 = ~n56 & ~n1211;
  assign n1213 = ~i_4_ & n139;
  assign n1214 = ~n1212 & n1213;
  assign n1215 = ~n55 & n1064;
  assign n1216 = n570 & n1215;
  assign n1217 = ~n1214 & ~n1216;
  assign n1218 = n644 & ~n1217;
  assign n1219 = n137 & n1086;
  assign n1220 = n520 & n1219;
  assign n1221 = n697 & n1052;
  assign n1222 = n290 & n1221;
  assign n1223 = ~n1220 & ~n1222;
  assign n1224 = n1114 & ~n1223;
  assign n1225 = n36 & n499;
  assign n1226 = n62 & n973;
  assign n1227 = n1225 & n1226;
  assign n1228 = n944 & n1145;
  assign n1229 = ~i_2_ & n1228;
  assign n1230 = ~n1227 & ~n1229;
  assign n1231 = ~n1224 & n1230;
  assign n1232 = ~n1218 & n1231;
  assign n1233 = ~i_9_ & n1232;
  assign n1234 = ~n1210 & ~n1233;
  assign n1235 = n1183 & ~n1234;
  assign n1236 = n1113 & n1235;
  assign n1237 = n191 & n441;
  assign n1238 = ~n144 & n1237;
  assign n1239 = ~n88 & ~n1238;
  assign n1240 = i_9_ & ~n1239;
  assign n1241 = i_11_ & n102;
  assign n1242 = n387 & ~n1241;
  assign n1243 = n146 & n760;
  assign n1244 = ~i_0_ & ~n244;
  assign n1245 = ~n249 & ~n1244;
  assign n1246 = n824 & ~n1245;
  assign n1247 = ~n1243 & ~n1246;
  assign n1248 = ~n1242 & n1247;
  assign n1249 = ~i_2_ & n965;
  assign n1250 = ~n178 & n182;
  assign n1251 = ~i_0_ & ~n1250;
  assign n1252 = ~n257 & ~n1251;
  assign n1253 = ~i_8_ & ~n1252;
  assign n1254 = ~n123 & ~n1253;
  assign n1255 = ~n1249 & n1254;
  assign n1256 = n571 & ~n1255;
  assign n1257 = n1248 & ~n1256;
  assign n1258 = ~n1240 & n1257;
  assign n1259 = n781 & ~n1258;
  assign n1260 = ~i_9_ & n973;
  assign n1261 = n1211 & n1260;
  assign n1262 = ~n105 & ~n1261;
  assign n1263 = n164 & ~n1262;
  assign n1264 = ~n139 & n1263;
  assign n1265 = n156 & n973;
  assign n1266 = i_2_ & n1265;
  assign n1267 = ~n1264 & ~n1266;
  assign n1268 = n138 & n290;
  assign n1269 = ~n197 & ~n1268;
  assign n1270 = n1106 & n1269;
  assign n1271 = n1063 & ~n1270;
  assign n1272 = n545 & n1120;
  assign n1273 = n1052 & n1058;
  assign n1274 = n1053 & n1057;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = ~n1272 & n1275;
  assign n1277 = n708 & ~n1276;
  assign n1278 = ~n1271 & ~n1277;
  assign n1279 = n1053 & n1067;
  assign n1280 = n227 & n637;
  assign n1281 = n943 & n1058;
  assign n1282 = n52 & n1120;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1280 & n1283;
  assign n1285 = ~n1279 & n1284;
  assign n1286 = n706 & ~n1285;
  assign n1287 = n290 & n484;
  assign n1288 = n943 & n1086;
  assign n1289 = n944 & n1067;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1287 & n1290;
  assign n1292 = n979 & ~n1291;
  assign n1293 = ~n1286 & ~n1292;
  assign n1294 = n1278 & n1293;
  assign n1295 = n1267 & n1294;
  assign n1296 = n440 & ~n1295;
  assign n1297 = n177 & ~n239;
  assign n1298 = n215 & n1297;
  assign n1299 = n743 & ~n1298;
  assign n1300 = ~n1296 & ~n1299;
  assign n1301 = ~n1259 & n1300;
  assign n1302 = ~n186 & n743;
  assign n1303 = n943 & n1120;
  assign n1304 = ~n1068 & ~n1303;
  assign n1305 = n356 & ~n1304;
  assign n1306 = n560 & n1067;
  assign n1307 = ~n546 & ~n1306;
  assign n1308 = n296 & ~n1307;
  assign n1309 = n251 & n1057;
  assign n1310 = ~n36 & n499;
  assign n1311 = ~n33 & n1310;
  assign n1312 = n1309 & n1311;
  assign n1313 = ~n1308 & ~n1312;
  assign n1314 = n484 & n644;
  assign n1315 = n1053 & n1314;
  assign n1316 = n560 & n943;
  assign n1317 = ~n557 & ~n1316;
  assign n1318 = n1058 & ~n1317;
  assign n1319 = ~n1315 & ~n1318;
  assign n1320 = n1313 & n1319;
  assign n1321 = ~n1305 & n1320;
  assign n1322 = i_9_ & n519;
  assign n1323 = ~n1321 & n1322;
  assign n1324 = n644 & ~n1291;
  assign n1325 = n503 & ~n1060;
  assign n1326 = n207 & n325;
  assign n1327 = n482 & n1326;
  assign n1328 = ~n1325 & ~n1327;
  assign n1329 = ~n1324 & n1328;
  assign n1330 = n997 & ~n1329;
  assign n1331 = ~i_6_ & n475;
  assign n1332 = ~n590 & ~n1331;
  assign n1333 = n585 & ~n1332;
  assign n1334 = ~i_7_ & n820;
  assign n1335 = n776 & n1334;
  assign n1336 = ~n1333 & ~n1335;
  assign n1337 = ~n1330 & n1336;
  assign n1338 = ~n1323 & n1337;
  assign n1339 = ~n1302 & n1338;
  assign n1340 = ~i_5_ & ~n1339;
  assign n1341 = n1301 & ~n1340;
  assign n1342 = n1236 & n1341;
  assign o_7_ = ~n1032 | ~n1342;
endmodule


