// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:22 2016

module TOP ( 
    Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_,
    Poutreg_59_, Poutreg_58_, Poutreg_57_, Poutreg_56_, Poutreg_55_,
    Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_,
    Poutreg_49_, Poutreg_48_, Poutreg_47_, Poutreg_46_, Poutreg_45_,
    Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_,
    Poutreg_39_, Poutreg_38_, Poutreg_37_, Poutreg_36_, Poutreg_35_,
    Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_,
    Poutreg_29_, Poutreg_28_, Poutreg_27_, Poutreg_26_, Poutreg_25_,
    Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_,
    Poutreg_19_, Poutreg_18_, Poutreg_17_, Poutreg_16_, Poutreg_15_,
    Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_,
    Poutreg_9_, Poutreg_8_, Poutreg_7_, Poutreg_6_, Poutreg_5_, Poutreg_4_,
    Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_,
    Pinreg_55_, Pinreg_54_, Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_,
    Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_,
    Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_,
    Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, Pinreg_33_, Pinreg_32_,
    Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_,
    Pinreg_25_, Pinreg_24_, Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_,
    Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_,
    Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_,
    Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, Pinreg_3_, Pinreg_2_,
    Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_,
    Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, Pdata_in_3_, Pdata_in_2_,
    Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_,
    Pdata_59_, Pdata_58_, Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_,
    Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_,
    Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_,
    Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, Pdata_37_, Pdata_36_,
    Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_,
    Pdata_29_, Pdata_28_, Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_,
    Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_,
    Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_,
    Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, Pdata_7_, Pdata_6_, Pdata_5_,
    Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_,
    PD_21_, PD_20_, PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_,
    PD_12_, PD_11_, PD_10_, PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_,
    PD_3_, PD_2_, PD_1_, PD_0_, PC_27_, PC_26_, PC_25_, PC_24_, PC_23_,
    PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, PC_17_, PC_16_, PC_15_, PC_14_,
    PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, PC_7_, PC_6_, PC_5_,
    PC_4_, PC_3_, PC_2_, PC_1_, PC_0_,
    Poutreg_new_63_, Poutreg_new_62_, Poutreg_new_61_, Poutreg_new_60_,
    Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_,
    Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_,
    Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_,
    Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_,
    Poutreg_new_43_, Poutreg_new_42_, Poutreg_new_41_, Poutreg_new_40_,
    Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_,
    Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_,
    Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_,
    Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_,
    Poutreg_new_23_, Poutreg_new_22_, Poutreg_new_21_, Poutreg_new_20_,
    Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_,
    Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_,
    Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_,
    Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_,
    Poutreg_new_3_, Poutreg_new_2_, Poutreg_new_1_, Poutreg_new_0_,
    Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_,
    Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_,
    Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_,
    Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_,
    Pinreg_new_39_, Pinreg_new_38_, Pinreg_new_37_, Pinreg_new_36_,
    Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_,
    Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_,
    Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_,
    Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_,
    Pinreg_new_19_, Pinreg_new_18_, Pinreg_new_17_, Pinreg_new_16_,
    Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_,
    Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_,
    Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_,
    Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_,
    Pencrypt_mode_new_0_, Pdata_new_63_, Pdata_new_62_, Pdata_new_61_,
    Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_,
    Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_,
    Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_,
    Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_,
    Pdata_new_44_, Pdata_new_43_, Pdata_new_42_, Pdata_new_41_,
    Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_,
    Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_,
    Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_,
    Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_,
    Pdata_new_24_, Pdata_new_23_, Pdata_new_22_, Pdata_new_21_,
    Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_,
    Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_,
    Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_,
    Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_,
    Pdata_new_3_, Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_,
    Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_,
    PD_new_25_, PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_,
    PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, PD_new_14_,
    PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_,
    PD_new_7_, PD_new_6_, PD_new_5_, PD_new_4_, PD_new_3_, PD_new_2_,
    PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_,
    PC_new_23_, PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_,
    PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, PC_new_12_,
    PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_,
    PC_new_5_, PC_new_4_, PC_new_3_, PC_new_2_, PC_new_1_, PC_new_0_  );
  input  Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_,
    Poutreg_59_, Poutreg_58_, Poutreg_57_, Poutreg_56_, Poutreg_55_,
    Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_,
    Poutreg_49_, Poutreg_48_, Poutreg_47_, Poutreg_46_, Poutreg_45_,
    Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_,
    Poutreg_39_, Poutreg_38_, Poutreg_37_, Poutreg_36_, Poutreg_35_,
    Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_,
    Poutreg_29_, Poutreg_28_, Poutreg_27_, Poutreg_26_, Poutreg_25_,
    Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_,
    Poutreg_19_, Poutreg_18_, Poutreg_17_, Poutreg_16_, Poutreg_15_,
    Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_,
    Poutreg_9_, Poutreg_8_, Poutreg_7_, Poutreg_6_, Poutreg_5_, Poutreg_4_,
    Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_,
    Pinreg_55_, Pinreg_54_, Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_,
    Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_,
    Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_,
    Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, Pinreg_33_, Pinreg_32_,
    Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_,
    Pinreg_25_, Pinreg_24_, Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_,
    Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_,
    Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_,
    Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, Pinreg_3_, Pinreg_2_,
    Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_,
    Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, Pdata_in_3_, Pdata_in_2_,
    Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_,
    Pdata_59_, Pdata_58_, Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_,
    Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_,
    Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_,
    Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, Pdata_37_, Pdata_36_,
    Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_,
    Pdata_29_, Pdata_28_, Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_,
    Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_,
    Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_,
    Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, Pdata_7_, Pdata_6_, Pdata_5_,
    Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_,
    PD_21_, PD_20_, PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_,
    PD_12_, PD_11_, PD_10_, PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_,
    PD_3_, PD_2_, PD_1_, PD_0_, PC_27_, PC_26_, PC_25_, PC_24_, PC_23_,
    PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, PC_17_, PC_16_, PC_15_, PC_14_,
    PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, PC_7_, PC_6_, PC_5_,
    PC_4_, PC_3_, PC_2_, PC_1_, PC_0_;
  output Poutreg_new_63_, Poutreg_new_62_, Poutreg_new_61_, Poutreg_new_60_,
    Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_,
    Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_,
    Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_,
    Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_,
    Poutreg_new_43_, Poutreg_new_42_, Poutreg_new_41_, Poutreg_new_40_,
    Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_,
    Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_,
    Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_,
    Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_,
    Poutreg_new_23_, Poutreg_new_22_, Poutreg_new_21_, Poutreg_new_20_,
    Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_,
    Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_,
    Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_,
    Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_,
    Poutreg_new_3_, Poutreg_new_2_, Poutreg_new_1_, Poutreg_new_0_,
    Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_,
    Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_,
    Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_,
    Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_,
    Pinreg_new_39_, Pinreg_new_38_, Pinreg_new_37_, Pinreg_new_36_,
    Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_,
    Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_,
    Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_,
    Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_,
    Pinreg_new_19_, Pinreg_new_18_, Pinreg_new_17_, Pinreg_new_16_,
    Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_,
    Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_,
    Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_,
    Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_,
    Pencrypt_mode_new_0_, Pdata_new_63_, Pdata_new_62_, Pdata_new_61_,
    Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_,
    Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_,
    Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_,
    Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_,
    Pdata_new_44_, Pdata_new_43_, Pdata_new_42_, Pdata_new_41_,
    Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_,
    Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_,
    Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_,
    Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_,
    Pdata_new_24_, Pdata_new_23_, Pdata_new_22_, Pdata_new_21_,
    Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_,
    Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_,
    Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_,
    Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_,
    Pdata_new_3_, Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_,
    Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_,
    PD_new_25_, PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_,
    PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, PD_new_14_,
    PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_,
    PD_new_7_, PD_new_6_, PD_new_5_, PD_new_4_, PD_new_3_, PD_new_2_,
    PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_,
    PC_new_23_, PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_,
    PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, PC_new_12_,
    PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_,
    PC_new_5_, PC_new_4_, PC_new_3_, PC_new_2_, PC_new_1_, PC_new_0_;
  wire n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n608, n609,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n724, n725, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n763, n764, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n873, n874, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n914, n915, n916, n917,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1020, n1021, n1022,
    n1023, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1055, n1056, n1057, n1058, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1101, n1102, n1103, n1104, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1224, n1225, n1226, n1227, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1335, n1336, n1337, n1338, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1375, n1376, n1377, n1378, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1416, n1417, n1418, n1419, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1448, n1449, n1450, n1451, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1481, n1482, n1483, n1484, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1592, n1593, n1594, n1595, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1623, n1624, n1625, n1626, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1656, n1657, n1658, n1659, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1701, n1702, n1703, n1704, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1735, n1736, n1737, n1738,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1769, n1770,
    n1771, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1881, n1882,
    n1883, n1884, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1922, n1923, n1924,
    n1925, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1960, n1961, n1962, n1963, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2005, n2006, n2007, n2008,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2030,
    n2031, n2032, n2033, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2061, n2062,
    n2063, n2064, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2092, n2093, n2094,
    n2095, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2126,
    n2127, n2128, n2129, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2159, n2160, n2161, n2162, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2190,
    n2191, n2192, n2193, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2223, n2224, n2225, n2226, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2254,
    n2255, n2256, n2257, n2259, n2260, n2262, n2263, n2265, n2266, n2268,
    n2269, n2271, n2272, n2274, n2275, n2277, n2278, n2280, n2281, n2283,
    n2284, n2286, n2287, n2289, n2290, n2292, n2293, n2295, n2296, n2298,
    n2299, n2301, n2302, n2304, n2305, n2307, n2308, n2310, n2311, n2313,
    n2314, n2316, n2317, n2319, n2320, n2322, n2323, n2325, n2326, n2328,
    n2329, n2331, n2332, n2334, n2335, n2337, n2338, n2340, n2341, n2343,
    n2344, n2346, n2347, n2349, n2350, n2352, n2353, n2355, n2356, n2358,
    n2359, n2361, n2362, n2364, n2365, n2367, n2368, n2370, n2371, n2373,
    n2374, n2376, n2377, n2379, n2380, n2382, n2383, n2385, n2386, n2388,
    n2389, n2391, n2392, n2394, n2395, n2397, n2398, n2400, n2401, n2403,
    n2404, n2406, n2407, n2409, n2410, n2412, n2413, n2415, n2416, n2418,
    n2419, n2421, n2422, n2424, n2425, n2427, n2428, n2430, n2431, n2433,
    n2434, n2436, n2437, n2439, n2440, n2442, n2443, n2445, n2446, n2448,
    n2449, n2451, n2452, n2454, n2455, n2457, n2458, n2460, n2461, n2463,
    n2464, n2466, n2467, n2469, n2470, n2472, n2473, n2475, n2476, n2478,
    n2479, n2481, n2482, n2484, n2485, n2487, n2488, n2490, n2491, n2493,
    n2494, n2496, n2497, n2499, n2500, n2502, n2503, n2505, n2506, n2508,
    n2509, n2511, n2512, n2514, n2515, n2517, n2518, n2520, n2521, n2523,
    n2524, n2526, n2527, n2529, n2530, n2532, n2533, n2535, n2536, n2538,
    n2539, n2541, n2542, n2544, n2545, n2547, n2548, n2550, n2551, n2553,
    n2554, n2556, n2557, n2559, n2560, n2562, n2563, n2565, n2566, n2568,
    n2569, n2571, n2572, n2574, n2575, n2577, n2578, n2580, n2581, n2583,
    n2584, n2586, n2587, n2589, n2590, n2592, n2593, n2595, n2596, n2598,
    n2599, n2601, n2602, n2604, n2605, n2607, n2608, n2610, n2611, n2613,
    n2614, n2616, n2617, n2619, n2620, n2622, n2623, n2625, n2626, n2628,
    n2629, n2630, n2631, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3201, n3202,
    n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
    n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381;
  assign n502 = Poutreg_63_ & ~Pcount_0_;
  assign n503 = Pcount_1_ & Pcount_0_;
  assign n504 = Pcount_2_ & n503;
  assign n505 = Pcount_3_ & n504;
  assign n506 = Pdata_52_ & ~PD_26_;
  assign n507 = ~Pdata_52_ & PD_26_;
  assign n508 = ~n506 & ~n507;
  assign n509 = Pdata_48_ & ~PD_23_;
  assign n510 = ~Pdata_48_ & PD_23_;
  assign n511 = ~n509 & ~n510;
  assign n512 = n508 & n511;
  assign n513 = Pdata_49_ & ~PD_2_;
  assign n514 = ~Pdata_49_ & PD_2_;
  assign n515 = ~n513 & ~n514;
  assign n516 = Pdata_47_ & ~PD_12_;
  assign n517 = ~Pdata_47_ & PD_12_;
  assign n518 = ~n516 & ~n517;
  assign n519 = Pdata_51_ & ~PD_18_;
  assign n520 = ~Pdata_51_ & PD_18_;
  assign n521 = ~n519 & ~n520;
  assign n522 = Pdata_50_ & ~PD_8_;
  assign n523 = ~Pdata_50_ & PD_8_;
  assign n524 = ~n522 & ~n523;
  assign n525 = n521 & ~n524;
  assign n526 = n518 & n525;
  assign n527 = ~n515 & n526;
  assign n528 = ~n521 & ~n524;
  assign n529 = n515 & n528;
  assign n530 = ~n518 & n529;
  assign n531 = ~n527 & ~n530;
  assign n532 = n512 & ~n531;
  assign n533 = ~n518 & n521;
  assign n534 = ~n528 & ~n533;
  assign n535 = ~n518 & ~n524;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n508 & ~n511;
  assign n538 = n518 & n524;
  assign n539 = ~n535 & ~n538;
  assign n540 = n537 & n539;
  assign n541 = ~n536 & ~n540;
  assign n542 = n508 & ~n511;
  assign n543 = ~n534 & ~n542;
  assign n544 = ~n541 & ~n543;
  assign n545 = n518 & ~n521;
  assign n546 = ~n533 & ~n545;
  assign n547 = n524 & ~n546;
  assign n548 = ~n508 & n511;
  assign n549 = n547 & n548;
  assign n550 = ~n544 & ~n549;
  assign n551 = n515 & ~n550;
  assign n552 = ~n532 & ~n551;
  assign n553 = ~n515 & n518;
  assign n554 = n512 & n553;
  assign n555 = n521 & n524;
  assign n556 = n554 & n555;
  assign n557 = ~n521 & n524;
  assign n558 = n553 & n557;
  assign n559 = ~n530 & ~n558;
  assign n560 = n548 & ~n559;
  assign n561 = ~n515 & ~n518;
  assign n562 = n512 & n561;
  assign n563 = n525 & n562;
  assign n564 = ~n560 & ~n563;
  assign n565 = ~n556 & n564;
  assign n566 = n552 & n565;
  assign n567 = ~n525 & ~n557;
  assign n568 = n537 & n567;
  assign n569 = n515 & ~n545;
  assign n570 = n568 & ~n569;
  assign n571 = n508 & n561;
  assign n572 = n555 & n571;
  assign n573 = n537 & n555;
  assign n574 = ~n518 & n573;
  assign n575 = ~n572 & ~n574;
  assign n576 = ~n570 & n575;
  assign n577 = ~n554 & n576;
  assign n578 = n548 & n561;
  assign n579 = ~n542 & ~n548;
  assign n580 = n515 & ~n579;
  assign n581 = n518 & n580;
  assign n582 = ~n578 & ~n581;
  assign n583 = n525 & ~n582;
  assign n584 = n542 & n561;
  assign n585 = n528 & n584;
  assign n586 = n557 & n578;
  assign n587 = ~n585 & ~n586;
  assign n588 = n518 & n555;
  assign n589 = n548 & n588;
  assign n590 = n515 & n589;
  assign n591 = n526 & n542;
  assign n592 = ~n515 & n591;
  assign n593 = ~n590 & ~n592;
  assign n594 = n587 & n593;
  assign n595 = n512 & ~n533;
  assign n596 = n569 & n595;
  assign n597 = ~n584 & ~n596;
  assign n598 = n524 & ~n597;
  assign n599 = n594 & ~n598;
  assign n600 = ~n583 & n599;
  assign n601 = n577 & n600;
  assign n602 = n566 & n601;
  assign n603 = Pdata_24_ & ~n602;
  assign n604 = ~Pdata_24_ & n602;
  assign n605 = ~n603 & ~n604;
  assign n606 = n505 & n605;
  assign Poutreg_new_63_ = n502 | n606;
  assign n608 = Poutreg_62_ & ~Pcount_0_;
  assign n609 = Pdata_56_ & n505;
  assign Poutreg_new_62_ = n608 | n609;
  assign n611 = Poutreg_61_ & ~Pcount_0_;
  assign n612 = Pdata_63_ & ~PC_13_;
  assign n613 = ~Pdata_63_ & PC_13_;
  assign n614 = ~n612 & ~n613;
  assign n615 = Pdata_35_ & ~PC_0_;
  assign n616 = ~Pdata_35_ & PC_0_;
  assign n617 = ~n615 & ~n616;
  assign n618 = Pdata_36_ & ~PC_4_;
  assign n619 = ~Pdata_36_ & PC_4_;
  assign n620 = ~n618 & ~n619;
  assign n621 = n617 & ~n620;
  assign n622 = Pdata_34_ & ~PC_23_;
  assign n623 = ~Pdata_34_ & PC_23_;
  assign n624 = ~n622 & ~n623;
  assign n625 = Pdata_32_ & ~PC_16_;
  assign n626 = ~Pdata_32_ & PC_16_;
  assign n627 = ~n625 & ~n626;
  assign n628 = Pdata_33_ & ~PC_10_;
  assign n629 = ~Pdata_33_ & PC_10_;
  assign n630 = ~n628 & ~n629;
  assign n631 = n627 & ~n630;
  assign n632 = ~n624 & n631;
  assign n633 = n621 & n632;
  assign n634 = n614 & n633;
  assign n635 = n617 & n627;
  assign n636 = n630 & n635;
  assign n637 = n614 & ~n624;
  assign n638 = n636 & n637;
  assign n639 = n620 & n638;
  assign n640 = ~n634 & ~n639;
  assign n641 = ~n614 & ~n617;
  assign n642 = ~n624 & ~n627;
  assign n643 = n641 & n642;
  assign n644 = ~n620 & ~n643;
  assign n645 = ~n620 & ~n630;
  assign n646 = n624 & n635;
  assign n647 = ~n614 & ~n630;
  assign n648 = n646 & n647;
  assign n649 = ~n645 & ~n648;
  assign n650 = ~n644 & ~n649;
  assign n651 = n614 & n624;
  assign n652 = n620 & n630;
  assign n653 = ~n645 & ~n652;
  assign n654 = ~n617 & n627;
  assign n655 = n653 & n654;
  assign n656 = n651 & n655;
  assign n657 = n617 & ~n627;
  assign n658 = n620 & ~n657;
  assign n659 = ~n620 & ~n635;
  assign n660 = ~n614 & n624;
  assign n661 = n630 & n660;
  assign n662 = ~n659 & n661;
  assign n663 = ~n658 & n662;
  assign n664 = ~n656 & ~n663;
  assign n665 = ~n650 & n664;
  assign n666 = n640 & n665;
  assign n667 = n632 & n641;
  assign n668 = ~n638 & ~n667;
  assign n669 = ~n620 & ~n668;
  assign n670 = n614 & n630;
  assign n671 = ~n617 & n620;
  assign n672 = n642 & n671;
  assign n673 = ~n647 & n672;
  assign n674 = ~n670 & n673;
  assign n675 = ~n669 & ~n674;
  assign n676 = n666 & n675;
  assign n677 = n620 & n624;
  assign n678 = n627 & ~n641;
  assign n679 = n677 & n678;
  assign n680 = ~n617 & ~n620;
  assign n681 = n637 & ~n680;
  assign n682 = ~n627 & n681;
  assign n683 = ~n621 & ~n671;
  assign n684 = ~n627 & n660;
  assign n685 = ~n683 & n684;
  assign n686 = ~n682 & ~n685;
  assign n687 = ~n679 & n686;
  assign n688 = n630 & ~n687;
  assign n689 = n624 & n627;
  assign n690 = ~n683 & n689;
  assign n691 = ~n624 & n657;
  assign n692 = ~n690 & ~n691;
  assign n693 = n647 & ~n692;
  assign n694 = ~n637 & ~n660;
  assign n695 = n620 & n694;
  assign n696 = n636 & n695;
  assign n697 = n614 & n645;
  assign n698 = n646 & n697;
  assign n699 = ~n614 & n630;
  assign n700 = ~n624 & n699;
  assign n701 = ~n627 & n680;
  assign n702 = n700 & n701;
  assign n703 = ~n698 & ~n702;
  assign n704 = ~n696 & n703;
  assign n705 = ~n693 & n704;
  assign n706 = ~n627 & n651;
  assign n707 = n627 & ~n694;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n631 & n680;
  assign n710 = ~n708 & n709;
  assign n711 = n614 & n620;
  assign n712 = n624 & ~n630;
  assign n713 = n657 & n712;
  assign n714 = n711 & n713;
  assign n715 = ~n710 & ~n714;
  assign n716 = n705 & n715;
  assign n717 = ~n688 & n716;
  assign n718 = n676 & n717;
  assign n719 = Pdata_16_ & ~n718;
  assign n720 = ~Pdata_16_ & n718;
  assign n721 = ~n719 & ~n720;
  assign n722 = n505 & n721;
  assign Poutreg_new_61_ = n611 | n722;
  assign n724 = Poutreg_60_ & ~Pcount_0_;
  assign n725 = Pdata_48_ & n505;
  assign Poutreg_new_60_ = n724 | n725;
  assign n727 = Poutreg_59_ & ~Pcount_0_;
  assign n728 = n617 & n620;
  assign n729 = ~n627 & ~n728;
  assign n730 = n627 & n683;
  assign n731 = n700 & ~n730;
  assign n732 = ~n729 & n731;
  assign n733 = ~n620 & n713;
  assign n734 = ~n627 & n670;
  assign n735 = ~n683 & n734;
  assign n736 = n660 & n680;
  assign n737 = n627 & n736;
  assign n738 = ~n735 & ~n737;
  assign n739 = ~n733 & n738;
  assign n740 = ~n732 & n739;
  assign n741 = n637 & n645;
  assign n742 = ~n677 & ~n741;
  assign n743 = ~n627 & ~n742;
  assign n744 = n632 & n711;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n617 & ~n745;
  assign n747 = ~n614 & n671;
  assign n748 = n614 & n728;
  assign n749 = ~n747 & ~n748;
  assign n750 = n632 & ~n749;
  assign n751 = n630 & n701;
  assign n752 = ~n694 & n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = n704 & n753;
  assign n755 = ~n746 & n754;
  assign n756 = n666 & n755;
  assign n757 = n740 & n756;
  assign n758 = Pdata_8_ & ~n757;
  assign n759 = ~Pdata_8_ & n757;
  assign n760 = ~n758 & ~n759;
  assign n761 = n505 & n760;
  assign Poutreg_new_59_ = n727 | n761;
  assign n763 = Poutreg_58_ & ~Pcount_0_;
  assign n764 = Pdata_40_ & n505;
  assign Poutreg_new_58_ = n763 | n764;
  assign n766 = Poutreg_57_ & ~Pcount_0_;
  assign n767 = Pdata_47_ & ~PC_12_;
  assign n768 = ~Pdata_47_ & PC_12_;
  assign n769 = ~n767 & ~n768;
  assign n770 = Pdata_48_ & ~PC_1_;
  assign n771 = ~Pdata_48_ & PC_1_;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n769 & ~n772;
  assign n774 = Pdata_46_ & ~PC_19_;
  assign n775 = ~Pdata_46_ & PC_19_;
  assign n776 = ~n774 & ~n775;
  assign n777 = Pdata_44_ & ~PC_6_;
  assign n778 = ~Pdata_44_ & PC_6_;
  assign n779 = ~n777 & ~n778;
  assign n780 = Pdata_45_ & ~PC_26_;
  assign n781 = ~Pdata_45_ & PC_26_;
  assign n782 = ~n780 & ~n781;
  assign n783 = Pdata_43_ & ~PC_15_;
  assign n784 = ~Pdata_43_ & PC_15_;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n782 & n785;
  assign n787 = n772 & n786;
  assign n788 = n779 & n787;
  assign n789 = ~n776 & n788;
  assign n790 = n769 & n789;
  assign n791 = n782 & ~n785;
  assign n792 = ~n772 & n776;
  assign n793 = n776 & ~n779;
  assign n794 = ~n792 & ~n793;
  assign n795 = n791 & ~n794;
  assign n796 = ~n790 & ~n795;
  assign n797 = ~n773 & ~n796;
  assign n798 = ~n779 & ~n782;
  assign n799 = ~n776 & n785;
  assign n800 = ~n769 & n799;
  assign n801 = n798 & n800;
  assign n802 = n769 & ~n779;
  assign n803 = n776 & n802;
  assign n804 = n791 & n803;
  assign n805 = ~n801 & ~n804;
  assign n806 = n772 & ~n805;
  assign n807 = ~n786 & ~n791;
  assign n808 = ~n769 & n779;
  assign n809 = ~n807 & n808;
  assign n810 = n792 & n809;
  assign n811 = ~n806 & ~n810;
  assign n812 = ~n791 & ~n799;
  assign n813 = n776 & ~n782;
  assign n814 = n779 & ~n813;
  assign n815 = n812 & n814;
  assign n816 = n769 & n772;
  assign n817 = ~n773 & ~n816;
  assign n818 = n815 & n817;
  assign n819 = n811 & ~n818;
  assign n820 = n776 & n782;
  assign n821 = n773 & n785;
  assign n822 = ~n779 & n821;
  assign n823 = n820 & n822;
  assign n824 = ~n769 & ~n785;
  assign n825 = n792 & n824;
  assign n826 = n798 & n825;
  assign n827 = n815 & n816;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n823 & n828;
  assign n830 = n779 & ~n782;
  assign n831 = n776 & n830;
  assign n832 = n772 & n824;
  assign n833 = n831 & n832;
  assign n834 = n773 & ~n785;
  assign n835 = ~n776 & n782;
  assign n836 = ~n779 & n835;
  assign n837 = n834 & n836;
  assign n838 = ~n833 & ~n837;
  assign n839 = n769 & ~n772;
  assign n840 = n779 & n782;
  assign n841 = n799 & n840;
  assign n842 = n839 & n841;
  assign n843 = n787 & n803;
  assign n844 = ~n842 & ~n843;
  assign n845 = n838 & n844;
  assign n846 = n829 & n845;
  assign n847 = n819 & n846;
  assign n848 = ~n772 & ~n802;
  assign n849 = n769 & n785;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~n824 & n850;
  assign n852 = n835 & n851;
  assign n853 = n830 & n834;
  assign n854 = ~n779 & n816;
  assign n855 = n807 & n854;
  assign n856 = ~n853 & ~n855;
  assign n857 = n776 & ~n856;
  assign n858 = n785 & n803;
  assign n859 = ~n800 & ~n858;
  assign n860 = ~n772 & ~n782;
  assign n861 = n800 & n840;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n859 & ~n862;
  assign n864 = ~n857 & ~n863;
  assign n865 = ~n852 & n864;
  assign n866 = n847 & n865;
  assign n867 = ~n797 & n866;
  assign n868 = Pdata_0_ & ~n867;
  assign n869 = ~Pdata_0_ & n867;
  assign n870 = ~n868 & ~n869;
  assign n871 = n505 & n870;
  assign Poutreg_new_57_ = n766 | n871;
  assign n873 = Poutreg_56_ & ~Pcount_0_;
  assign n874 = Pdata_32_ & n505;
  assign Poutreg_new_56_ = n873 | n874;
  assign n876 = n776 & n840;
  assign n877 = n821 & n876;
  assign n878 = n845 & ~n877;
  assign n879 = ~n789 & n878;
  assign n880 = ~n776 & n802;
  assign n881 = n786 & n880;
  assign n882 = ~n772 & n881;
  assign n883 = n816 & n841;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n776 & n798;
  assign n886 = n834 & n885;
  assign n887 = n832 & n836;
  assign n888 = ~n886 & ~n887;
  assign n889 = n884 & n888;
  assign n890 = n772 & n840;
  assign n891 = ~n779 & n792;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n831 & n892;
  assign n894 = n769 & ~n893;
  assign n895 = ~n785 & n894;
  assign n896 = n889 & ~n895;
  assign n897 = ~n822 & n856;
  assign n898 = ~n776 & ~n897;
  assign n899 = ~n769 & n793;
  assign n900 = n786 & n899;
  assign n901 = ~n898 & ~n900;
  assign n902 = n896 & n901;
  assign n903 = n819 & n902;
  assign n904 = n879 & n903;
  assign n905 = Pdata_25_ & ~n904;
  assign n906 = ~Pdata_25_ & n904;
  assign n907 = ~n905 & ~n906;
  assign n908 = n505 & n907;
  assign n909 = Pcount_0_ & ~n505;
  assign n910 = Poutreg_63_ & n909;
  assign n911 = Poutreg_55_ & ~Pcount_0_;
  assign n912 = ~n910 & ~n911;
  assign Poutreg_new_55_ = n908 | ~n912;
  assign n914 = Poutreg_62_ & n909;
  assign n915 = Poutreg_54_ & ~Pcount_0_;
  assign n916 = Pdata_57_ & n505;
  assign n917 = ~n915 & ~n916;
  assign Poutreg_new_54_ = n914 | ~n917;
  assign n919 = Pdata_36_ & ~PC_27_;
  assign n920 = ~Pdata_36_ & PC_27_;
  assign n921 = ~n919 & ~n920;
  assign n922 = Pdata_35_ & ~PC_2_;
  assign n923 = ~Pdata_35_ & PC_2_;
  assign n924 = ~n922 & ~n923;
  assign n925 = n921 & ~n924;
  assign n926 = Pdata_38_ & ~PC_5_;
  assign n927 = ~Pdata_38_ & PC_5_;
  assign n928 = ~n926 & ~n927;
  assign n929 = Pdata_39_ & ~PC_20_;
  assign n930 = ~Pdata_39_ & PC_20_;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n928 & ~n931;
  assign n933 = Pdata_40_ & ~PC_9_;
  assign n934 = ~Pdata_40_ & PC_9_;
  assign n935 = ~n933 & ~n934;
  assign n936 = Pdata_37_ & ~PC_14_;
  assign n937 = ~Pdata_37_ & PC_14_;
  assign n938 = ~n936 & ~n937;
  assign n939 = n935 & n938;
  assign n940 = n932 & n939;
  assign n941 = n925 & n940;
  assign n942 = n928 & n931;
  assign n943 = ~n935 & n942;
  assign n944 = ~n924 & n938;
  assign n945 = n943 & n944;
  assign n946 = ~n921 & n945;
  assign n947 = ~n941 & ~n946;
  assign n948 = ~n921 & n924;
  assign n949 = ~n935 & ~n938;
  assign n950 = ~n928 & n931;
  assign n951 = n949 & n950;
  assign n952 = n948 & n951;
  assign n953 = n935 & ~n938;
  assign n954 = n921 & n924;
  assign n955 = n928 & ~n931;
  assign n956 = n954 & n955;
  assign n957 = n953 & n956;
  assign n958 = ~n952 & ~n957;
  assign n959 = n947 & n958;
  assign n960 = n938 & n954;
  assign n961 = n943 & n960;
  assign n962 = n932 & ~n935;
  assign n963 = n960 & n962;
  assign n964 = ~n921 & ~n924;
  assign n965 = ~n935 & n950;
  assign n966 = n938 & n965;
  assign n967 = n964 & n966;
  assign n968 = n925 & n950;
  assign n969 = n948 & n955;
  assign n970 = ~n968 & ~n969;
  assign n971 = n939 & ~n970;
  assign n972 = ~n967 & ~n971;
  assign n973 = ~n963 & n972;
  assign n974 = ~n961 & n973;
  assign n975 = n959 & n974;
  assign n976 = n953 & n964;
  assign n977 = n932 & n976;
  assign n978 = ~n939 & ~n949;
  assign n979 = ~n935 & n955;
  assign n980 = n925 & n979;
  assign n981 = n942 & n954;
  assign n982 = ~n980 & ~n981;
  assign n983 = ~n978 & ~n982;
  assign n984 = ~n977 & ~n983;
  assign n985 = ~n931 & n949;
  assign n986 = ~n966 & ~n985;
  assign n987 = ~n921 & ~n986;
  assign n988 = ~n921 & n942;
  assign n989 = ~n956 & ~n988;
  assign n990 = n939 & ~n989;
  assign n991 = ~n987 & ~n990;
  assign n992 = n984 & n991;
  assign n993 = n932 & n978;
  assign n994 = n942 & n949;
  assign n995 = ~n993 & ~n994;
  assign n996 = n925 & ~n995;
  assign n997 = ~n924 & ~n928;
  assign n998 = ~n950 & ~n964;
  assign n999 = n953 & ~n998;
  assign n1000 = ~n997 & n999;
  assign n1001 = ~n996 & ~n1000;
  assign n1002 = n921 & n945;
  assign n1003 = n960 & n979;
  assign n1004 = n940 & n948;
  assign n1005 = n953 & n968;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1003 & n1006;
  assign n1008 = ~n1002 & n1007;
  assign n1009 = n1001 & n1008;
  assign n1010 = n992 & n1009;
  assign n1011 = n975 & n1010;
  assign n1012 = Pdata_17_ & ~n1011;
  assign n1013 = ~Pdata_17_ & n1011;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = n505 & n1014;
  assign n1016 = Poutreg_61_ & n909;
  assign n1017 = Poutreg_53_ & ~Pcount_0_;
  assign n1018 = ~n1016 & ~n1017;
  assign Poutreg_new_53_ = n1015 | ~n1018;
  assign n1020 = Poutreg_60_ & n909;
  assign n1021 = Poutreg_52_ & ~Pcount_0_;
  assign n1022 = Pdata_49_ & n505;
  assign n1023 = ~n1021 & ~n1022;
  assign Poutreg_new_52_ = n1020 | ~n1023;
  assign n1025 = n791 & n802;
  assign n1026 = n785 & n808;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~n820 & ~n1027;
  assign n1029 = n807 & n899;
  assign n1030 = n772 & ~n1029;
  assign n1031 = ~n1028 & n1030;
  assign n1032 = n807 & n880;
  assign n1033 = ~n900 & ~n1032;
  assign n1034 = ~n772 & n1033;
  assign n1035 = ~n1031 & ~n1034;
  assign n1036 = ~n785 & n876;
  assign n1037 = n831 & n839;
  assign n1038 = n834 & n835;
  assign n1039 = n800 & n830;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = ~n1037 & n1040;
  assign n1042 = ~n1036 & n1041;
  assign n1043 = ~n1035 & n1042;
  assign n1044 = n811 & n889;
  assign n1045 = n846 & n1044;
  assign n1046 = n1043 & n1045;
  assign n1047 = Pdata_9_ & ~n1046;
  assign n1048 = ~Pdata_9_ & n1046;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = n505 & n1049;
  assign n1051 = Poutreg_59_ & n909;
  assign n1052 = Poutreg_51_ & ~Pcount_0_;
  assign n1053 = ~n1051 & ~n1052;
  assign Poutreg_new_51_ = n1050 | ~n1053;
  assign n1055 = Poutreg_58_ & n909;
  assign n1056 = Pdata_41_ & n505;
  assign n1057 = Poutreg_50_ & ~Pcount_0_;
  assign n1058 = ~n1056 & ~n1057;
  assign Poutreg_new_50_ = n1055 | ~n1058;
  assign n1060 = n932 & n935;
  assign n1061 = ~n979 & ~n1060;
  assign n1062 = ~n921 & ~n1061;
  assign n1063 = ~n965 & ~n1062;
  assign n1064 = n944 & ~n1063;
  assign n1065 = n975 & ~n1064;
  assign n1066 = n951 & n964;
  assign n1067 = n932 & n954;
  assign n1068 = ~n938 & ~n1067;
  assign n1069 = ~n924 & n955;
  assign n1070 = n921 & n1069;
  assign n1071 = ~n1067 & ~n1070;
  assign n1072 = ~n1068 & ~n1071;
  assign n1073 = ~n978 & n1072;
  assign n1074 = n984 & ~n1073;
  assign n1075 = ~n1066 & n1074;
  assign n1076 = n939 & n950;
  assign n1077 = n995 & ~n1076;
  assign n1078 = n948 & ~n1077;
  assign n1079 = ~n950 & ~n955;
  assign n1080 = n976 & ~n1079;
  assign n1081 = ~n1078 & ~n1080;
  assign n1082 = ~n924 & ~n942;
  assign n1083 = ~n962 & n1082;
  assign n1084 = n921 & ~n938;
  assign n1085 = n931 & n935;
  assign n1086 = n924 & ~n1085;
  assign n1087 = ~n979 & n1086;
  assign n1088 = n1084 & ~n1087;
  assign n1089 = ~n1083 & n1088;
  assign n1090 = n1081 & ~n1089;
  assign n1091 = n1075 & n1090;
  assign n1092 = n1065 & n1091;
  assign n1093 = ~Pdata_1_ & ~n1092;
  assign n1094 = Pdata_1_ & n1092;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = n505 & ~n1095;
  assign n1097 = Poutreg_57_ & n909;
  assign n1098 = Poutreg_49_ & ~Pcount_0_;
  assign n1099 = ~n1097 & ~n1098;
  assign Poutreg_new_49_ = n1096 | ~n1099;
  assign n1101 = Poutreg_56_ & n909;
  assign n1102 = Pdata_33_ & n505;
  assign n1103 = Poutreg_48_ & ~Pcount_0_;
  assign n1104 = ~n1102 & ~n1103;
  assign Poutreg_new_48_ = n1101 | ~n1104;
  assign n1106 = Pdata_63_ & ~PD_0_;
  assign n1107 = ~Pdata_63_ & PD_0_;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = Pdata_62_ & ~PD_7_;
  assign n1110 = ~Pdata_62_ & PD_7_;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = Pdata_60_ & ~PD_13_;
  assign n1113 = ~Pdata_60_ & PD_13_;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = Pdata_61_ & ~PD_21_;
  assign n1116 = ~Pdata_61_ & PD_21_;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = n1114 & ~n1117;
  assign n1119 = n1111 & n1118;
  assign n1120 = ~n1108 & n1119;
  assign n1121 = Pdata_32_ & ~PD_3_;
  assign n1122 = ~Pdata_32_ & PD_3_;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = Pdata_59_ & ~PD_17_;
  assign n1125 = ~Pdata_59_ & PD_17_;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = n1123 & ~n1126;
  assign n1128 = n1120 & n1127;
  assign n1129 = ~n1117 & n1123;
  assign n1130 = n1111 & n1126;
  assign n1131 = n1108 & n1130;
  assign n1132 = n1129 & n1131;
  assign n1133 = n1108 & ~n1114;
  assign n1134 = ~n1117 & ~n1126;
  assign n1135 = ~n1111 & n1134;
  assign n1136 = ~n1129 & ~n1135;
  assign n1137 = n1133 & ~n1136;
  assign n1138 = ~n1132 & ~n1137;
  assign n1139 = ~n1114 & n1117;
  assign n1140 = n1130 & n1139;
  assign n1141 = ~n1108 & ~n1114;
  assign n1142 = n1111 & n1141;
  assign n1143 = ~n1126 & n1142;
  assign n1144 = n1117 & n1126;
  assign n1145 = n1133 & n1144;
  assign n1146 = ~n1143 & ~n1145;
  assign n1147 = ~n1108 & ~n1111;
  assign n1148 = n1126 & n1147;
  assign n1149 = n1118 & n1148;
  assign n1150 = n1146 & ~n1149;
  assign n1151 = ~n1140 & n1150;
  assign n1152 = ~n1123 & ~n1151;
  assign n1153 = n1123 & n1148;
  assign n1154 = ~n1143 & ~n1153;
  assign n1155 = n1117 & ~n1154;
  assign n1156 = ~n1111 & ~n1123;
  assign n1157 = n1111 & n1117;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = n1108 & n1114;
  assign n1160 = ~n1129 & n1159;
  assign n1161 = n1158 & n1160;
  assign n1162 = ~n1126 & n1161;
  assign n1163 = ~n1155 & ~n1162;
  assign n1164 = ~n1152 & n1163;
  assign n1165 = n1138 & n1164;
  assign n1166 = ~n1108 & n1114;
  assign n1167 = n1117 & n1166;
  assign n1168 = ~n1126 & n1156;
  assign n1169 = n1167 & n1168;
  assign n1170 = n1111 & ~n1126;
  assign n1171 = n1117 & n1159;
  assign n1172 = n1170 & n1171;
  assign n1173 = n1123 & n1172;
  assign n1174 = ~n1169 & ~n1173;
  assign n1175 = ~n1114 & ~n1117;
  assign n1176 = n1153 & n1175;
  assign n1177 = n1108 & n1126;
  assign n1178 = n1118 & n1177;
  assign n1179 = n1156 & n1178;
  assign n1180 = ~n1176 & ~n1179;
  assign n1181 = n1174 & n1180;
  assign n1182 = n1111 & ~n1123;
  assign n1183 = ~n1111 & n1123;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = n1135 & n1166;
  assign n1186 = n1144 & n1159;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = n1184 & ~n1187;
  assign n1189 = n1139 & n1147;
  assign n1190 = n1127 & n1189;
  assign n1191 = ~n1188 & ~n1190;
  assign n1192 = n1181 & n1191;
  assign n1193 = n1117 & ~n1123;
  assign n1194 = ~n1129 & ~n1193;
  assign n1195 = n1133 & n1170;
  assign n1196 = n1130 & n1167;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1194 & ~n1197;
  assign n1199 = n1123 & n1126;
  assign n1200 = n1120 & n1199;
  assign n1201 = ~n1198 & ~n1200;
  assign n1202 = n1134 & n1159;
  assign n1203 = n1183 & n1202;
  assign n1204 = ~n1108 & n1175;
  assign n1205 = ~n1123 & n1130;
  assign n1206 = n1204 & n1205;
  assign n1207 = ~n1203 & ~n1206;
  assign n1208 = n1168 & n1171;
  assign n1209 = n1139 & n1153;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = n1207 & n1210;
  assign n1212 = n1201 & n1211;
  assign n1213 = n1192 & n1212;
  assign n1214 = n1165 & n1213;
  assign n1215 = ~n1128 & n1214;
  assign n1216 = Pdata_26_ & ~n1215;
  assign n1217 = ~Pdata_26_ & n1215;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n505 & n1218;
  assign n1220 = Poutreg_55_ & n909;
  assign n1221 = Poutreg_47_ & ~Pcount_0_;
  assign n1222 = ~n1220 & ~n1221;
  assign Poutreg_new_47_ = n1219 | ~n1222;
  assign n1224 = Poutreg_54_ & n909;
  assign n1225 = Pdata_58_ & n505;
  assign n1226 = Poutreg_46_ & ~Pcount_0_;
  assign n1227 = ~n1225 & ~n1226;
  assign Poutreg_new_46_ = n1224 | ~n1227;
  assign n1229 = Pdata_53_ & ~PD_22_;
  assign n1230 = ~Pdata_53_ & PD_22_;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = Pdata_52_ & ~PD_11_;
  assign n1233 = ~Pdata_52_ & PD_11_;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = Pdata_54_ & ~PD_16_;
  assign n1236 = ~Pdata_54_ & PD_16_;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = Pdata_55_ & ~PD_4_;
  assign n1239 = ~Pdata_55_ & PD_4_;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = Pdata_51_ & ~PD_1_;
  assign n1242 = ~Pdata_51_ & PD_1_;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = n1240 & n1243;
  assign n1245 = ~n1237 & n1244;
  assign n1246 = n1240 & ~n1243;
  assign n1247 = Pdata_56_ & ~PD_19_;
  assign n1248 = ~Pdata_56_ & PD_19_;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = n1237 & n1249;
  assign n1251 = n1246 & n1250;
  assign n1252 = ~n1245 & ~n1251;
  assign n1253 = ~n1234 & ~n1252;
  assign n1254 = n1234 & n1249;
  assign n1255 = n1237 & n1243;
  assign n1256 = n1240 & n1255;
  assign n1257 = n1254 & n1256;
  assign n1258 = n1234 & ~n1249;
  assign n1259 = ~n1237 & ~n1243;
  assign n1260 = ~n1255 & ~n1259;
  assign n1261 = n1258 & n1260;
  assign n1262 = ~n1257 & ~n1261;
  assign n1263 = ~n1253 & n1262;
  assign n1264 = ~n1231 & ~n1263;
  assign n1265 = ~n1240 & n1259;
  assign n1266 = ~n1234 & ~n1249;
  assign n1267 = ~n1231 & n1266;
  assign n1268 = n1265 & n1267;
  assign n1269 = n1231 & n1266;
  assign n1270 = n1245 & n1269;
  assign n1271 = ~n1268 & ~n1270;
  assign n1272 = ~n1234 & n1249;
  assign n1273 = ~n1231 & n1272;
  assign n1274 = ~n1240 & ~n1243;
  assign n1275 = n1237 & n1274;
  assign n1276 = n1273 & n1275;
  assign n1277 = ~n1240 & n1255;
  assign n1278 = n1231 & n1272;
  assign n1279 = n1277 & n1278;
  assign n1280 = ~n1276 & ~n1279;
  assign n1281 = n1271 & n1280;
  assign n1282 = ~n1240 & n1243;
  assign n1283 = ~n1246 & ~n1282;
  assign n1284 = ~n1237 & ~n1283;
  assign n1285 = n1273 & n1284;
  assign n1286 = n1267 & n1277;
  assign n1287 = n1237 & n1246;
  assign n1288 = n1269 & n1287;
  assign n1289 = ~n1286 & ~n1288;
  assign n1290 = ~n1285 & n1289;
  assign n1291 = n1281 & n1290;
  assign n1292 = ~n1264 & n1291;
  assign n1293 = ~n1237 & ~n1249;
  assign n1294 = ~n1250 & ~n1293;
  assign n1295 = n1234 & n1294;
  assign n1296 = n1274 & n1295;
  assign n1297 = n1245 & n1249;
  assign n1298 = ~n1234 & n1297;
  assign n1299 = ~n1296 & ~n1298;
  assign n1300 = n1273 & n1277;
  assign n1301 = n1278 & n1287;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = n1231 & n1254;
  assign n1304 = n1284 & n1303;
  assign n1305 = n1231 & n1258;
  assign n1306 = n1277 & n1305;
  assign n1307 = ~n1237 & n1240;
  assign n1308 = ~n1243 & n1307;
  assign n1309 = ~n1231 & n1258;
  assign n1310 = n1308 & n1309;
  assign n1311 = ~n1306 & ~n1310;
  assign n1312 = ~n1304 & n1311;
  assign n1313 = n1265 & n1269;
  assign n1314 = n1256 & n1309;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = n1312 & n1315;
  assign n1317 = n1302 & n1316;
  assign n1318 = ~n1277 & ~n1308;
  assign n1319 = n1269 & ~n1318;
  assign n1320 = n1237 & n1254;
  assign n1321 = ~n1283 & n1320;
  assign n1322 = n1231 & n1321;
  assign n1323 = ~n1319 & ~n1322;
  assign n1324 = n1317 & n1323;
  assign n1325 = n1299 & n1324;
  assign n1326 = n1292 & n1325;
  assign n1327 = Pdata_18_ & ~n1326;
  assign n1328 = ~Pdata_18_ & n1326;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = n505 & n1329;
  assign n1331 = Poutreg_53_ & n909;
  assign n1332 = Poutreg_45_ & ~Pcount_0_;
  assign n1333 = ~n1331 & ~n1332;
  assign Poutreg_new_45_ = n1330 | ~n1333;
  assign n1335 = Poutreg_52_ & n909;
  assign n1336 = Poutreg_44_ & ~Pcount_0_;
  assign n1337 = Pdata_50_ & n505;
  assign n1338 = ~n1336 & ~n1337;
  assign Poutreg_new_44_ = n1335 | ~n1338;
  assign n1340 = ~n1275 & ~n1284;
  assign n1341 = n1305 & ~n1340;
  assign n1342 = n1234 & n1265;
  assign n1343 = ~n1321 & ~n1342;
  assign n1344 = ~n1231 & ~n1343;
  assign n1345 = ~n1240 & n1260;
  assign n1346 = n1269 & n1345;
  assign n1347 = n1275 & n1303;
  assign n1348 = n1256 & n1273;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1346 & n1349;
  assign n1351 = ~n1344 & n1350;
  assign n1352 = ~n1341 & n1351;
  assign n1353 = n1265 & n1272;
  assign n1354 = n1254 & n1307;
  assign n1355 = n1243 & n1354;
  assign n1356 = ~n1353 & ~n1355;
  assign n1357 = n1231 & ~n1293;
  assign n1358 = n1244 & n1357;
  assign n1359 = ~n1250 & n1358;
  assign n1360 = n1260 & n1267;
  assign n1361 = n1240 & n1360;
  assign n1362 = ~n1359 & ~n1361;
  assign n1363 = n1356 & n1362;
  assign n1364 = n1317 & n1363;
  assign n1365 = n1290 & n1364;
  assign n1366 = n1352 & n1365;
  assign n1367 = Pdata_10_ & ~n1366;
  assign n1368 = ~Pdata_10_ & n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = n505 & n1369;
  assign n1371 = Poutreg_51_ & n909;
  assign n1372 = Poutreg_43_ & ~Pcount_0_;
  assign n1373 = ~n1371 & ~n1372;
  assign Poutreg_new_43_ = n1370 | ~n1373;
  assign n1375 = Poutreg_50_ & n909;
  assign n1376 = Poutreg_42_ & ~Pcount_0_;
  assign n1377 = Pdata_42_ & n505;
  assign n1378 = ~n1376 & ~n1377;
  assign Poutreg_new_42_ = n1375 | ~n1378;
  assign n1380 = ~n515 & n537;
  assign n1381 = ~n539 & n1380;
  assign n1382 = ~n530 & ~n1381;
  assign n1383 = ~n515 & n528;
  assign n1384 = ~n579 & n1383;
  assign n1385 = ~n573 & ~n1384;
  assign n1386 = n518 & ~n1385;
  assign n1387 = n542 & n557;
  assign n1388 = ~n553 & n1387;
  assign n1389 = n555 & n578;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = ~n1386 & n1390;
  assign n1392 = n1382 & n1391;
  assign n1393 = n542 & n555;
  assign n1394 = n553 & n1393;
  assign n1395 = n557 & n562;
  assign n1396 = n528 & n561;
  assign n1397 = ~n527 & ~n1396;
  assign n1398 = n548 & ~n1397;
  assign n1399 = ~n1395 & ~n1398;
  assign n1400 = ~n1394 & n1399;
  assign n1401 = ~n524 & ~n546;
  assign n1402 = n512 & n1401;
  assign n1403 = ~n591 & ~n1402;
  assign n1404 = n515 & ~n1403;
  assign n1405 = n1400 & ~n1404;
  assign n1406 = n1392 & n1405;
  assign n1407 = n566 & n1406;
  assign n1408 = ~Pdata_2_ & ~n1407;
  assign n1409 = Pdata_2_ & n1407;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = n505 & ~n1410;
  assign n1412 = Poutreg_49_ & n909;
  assign n1413 = Poutreg_41_ & ~Pcount_0_;
  assign n1414 = ~n1412 & ~n1413;
  assign Poutreg_new_41_ = n1411 | ~n1414;
  assign n1416 = Poutreg_48_ & n909;
  assign n1417 = Poutreg_40_ & ~Pcount_0_;
  assign n1418 = Pdata_34_ & n505;
  assign n1419 = ~n1417 & ~n1418;
  assign Poutreg_new_40_ = n1416 | ~n1419;
  assign n1421 = n1008 & n1075;
  assign n1422 = n924 & n942;
  assign n1423 = ~n1069 & ~n1422;
  assign n1424 = ~n935 & ~n1423;
  assign n1425 = n924 & ~n938;
  assign n1426 = ~n944 & ~n1425;
  assign n1427 = n932 & ~n953;
  assign n1428 = ~n1085 & ~n1427;
  assign n1429 = ~n1426 & ~n1428;
  assign n1430 = ~n1424 & ~n1429;
  assign n1431 = ~n921 & ~n1430;
  assign n1432 = n1071 & ~n1422;
  assign n1433 = n953 & ~n1432;
  assign n1434 = n921 & n1426;
  assign n1435 = n965 & n1434;
  assign n1436 = ~n1433 & ~n1435;
  assign n1437 = ~n1431 & n1436;
  assign n1438 = n973 & n1437;
  assign n1439 = n1421 & n1438;
  assign n1440 = Pdata_27_ & ~n1439;
  assign n1441 = ~Pdata_27_ & n1439;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = n505 & n1442;
  assign n1444 = Poutreg_47_ & n909;
  assign n1445 = Poutreg_39_ & ~Pcount_0_;
  assign n1446 = ~n1444 & ~n1445;
  assign Poutreg_new_39_ = n1443 | ~n1446;
  assign n1448 = Poutreg_46_ & n909;
  assign n1449 = Pdata_59_ & n505;
  assign n1450 = Poutreg_38_ & ~Pcount_0_;
  assign n1451 = ~n1449 & ~n1450;
  assign Poutreg_new_38_ = n1448 | ~n1451;
  assign n1453 = ~n800 & ~n825;
  assign n1454 = ~n779 & ~n1453;
  assign n1455 = ~n802 & ~n808;
  assign n1456 = ~n776 & ~n1455;
  assign n1457 = ~n849 & n1456;
  assign n1458 = ~n858 & ~n1457;
  assign n1459 = ~n772 & ~n1458;
  assign n1460 = ~n1454 & ~n1459;
  assign n1461 = n782 & ~n1460;
  assign n1462 = ~n876 & ~n885;
  assign n1463 = n832 & ~n1462;
  assign n1464 = n785 & n1037;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = n813 & n851;
  assign n1467 = ~n818 & ~n881;
  assign n1468 = ~n1466 & n1467;
  assign n1469 = n1465 & n1468;
  assign n1470 = n1044 & n1469;
  assign n1471 = n829 & n1470;
  assign n1472 = ~n1461 & n1471;
  assign n1473 = Pdata_19_ & ~n1472;
  assign n1474 = ~Pdata_19_ & n1472;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n505 & n1475;
  assign n1477 = Poutreg_45_ & n909;
  assign n1478 = Poutreg_37_ & ~Pcount_0_;
  assign n1479 = ~n1477 & ~n1478;
  assign Poutreg_new_37_ = n1476 | ~n1479;
  assign n1481 = Poutreg_44_ & n909;
  assign n1482 = Pdata_51_ & n505;
  assign n1483 = Poutreg_36_ & ~Pcount_0_;
  assign n1484 = ~n1482 & ~n1483;
  assign Poutreg_new_36_ = n1481 | ~n1484;
  assign n1486 = Pdata_56_ & ~PD_20_;
  assign n1487 = ~Pdata_56_ & PD_20_;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = Pdata_58_ & ~PD_27_;
  assign n1490 = ~Pdata_58_ & PD_27_;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = n1488 & n1491;
  assign n1493 = Pdata_57_ & ~PD_10_;
  assign n1494 = ~Pdata_57_ & PD_10_;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = Pdata_60_ & ~PD_24_;
  assign n1497 = ~Pdata_60_ & PD_24_;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = n1495 & ~n1498;
  assign n1500 = ~n1495 & n1498;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = Pdata_55_ & ~PD_15_;
  assign n1503 = ~Pdata_55_ & PD_15_;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = Pdata_59_ & ~PD_5_;
  assign n1506 = ~Pdata_59_ & PD_5_;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = n1504 & ~n1507;
  assign n1509 = ~n1504 & n1507;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = n1501 & n1510;
  assign n1512 = n1492 & n1511;
  assign n1513 = n1495 & n1498;
  assign n1514 = ~n1488 & ~n1491;
  assign n1515 = n1509 & n1514;
  assign n1516 = n1513 & n1515;
  assign n1517 = n1504 & n1507;
  assign n1518 = ~n1488 & n1500;
  assign n1519 = n1517 & n1518;
  assign n1520 = ~n1516 & ~n1519;
  assign n1521 = n1495 & n1504;
  assign n1522 = n1514 & n1521;
  assign n1523 = ~n1498 & n1522;
  assign n1524 = n1492 & n1509;
  assign n1525 = ~n1501 & n1524;
  assign n1526 = ~n1523 & ~n1525;
  assign n1527 = n1520 & n1526;
  assign n1528 = ~n1512 & n1527;
  assign n1529 = n1488 & ~n1491;
  assign n1530 = n1509 & n1529;
  assign n1531 = n1500 & n1530;
  assign n1532 = n1521 & n1529;
  assign n1533 = ~n1498 & n1532;
  assign n1534 = n1498 & n1522;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = ~n1507 & ~n1535;
  assign n1537 = ~n1504 & ~n1507;
  assign n1538 = ~n1495 & ~n1498;
  assign n1539 = n1529 & n1538;
  assign n1540 = n1537 & n1539;
  assign n1541 = ~n1536 & ~n1540;
  assign n1542 = ~n1531 & n1541;
  assign n1543 = ~n1488 & n1491;
  assign n1544 = n1513 & n1537;
  assign n1545 = n1543 & n1544;
  assign n1546 = n1538 & n1543;
  assign n1547 = n1508 & n1546;
  assign n1548 = ~n1545 & ~n1547;
  assign n1549 = n1499 & n1537;
  assign n1550 = n1514 & n1549;
  assign n1551 = n1492 & n1517;
  assign n1552 = n1500 & n1551;
  assign n1553 = ~n1550 & ~n1552;
  assign n1554 = n1548 & n1553;
  assign n1555 = ~n1491 & n1538;
  assign n1556 = ~n1488 & n1555;
  assign n1557 = n1498 & n1543;
  assign n1558 = n1521 & n1557;
  assign n1559 = ~n1556 & ~n1558;
  assign n1560 = ~n1501 & n1543;
  assign n1561 = ~n1504 & n1560;
  assign n1562 = n1559 & ~n1561;
  assign n1563 = ~n1507 & ~n1562;
  assign n1564 = n1554 & ~n1563;
  assign n1565 = n1500 & n1508;
  assign n1566 = ~n1544 & ~n1565;
  assign n1567 = n1529 & ~n1566;
  assign n1568 = ~n1530 & ~n1551;
  assign n1569 = n1499 & ~n1568;
  assign n1570 = ~n1567 & ~n1569;
  assign n1571 = n1500 & n1537;
  assign n1572 = n1508 & n1513;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = n1529 & ~n1573;
  assign n1575 = n1499 & n1543;
  assign n1576 = n1517 & n1575;
  assign n1577 = n1509 & n1546;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = ~n1574 & n1578;
  assign n1580 = n1570 & n1579;
  assign n1581 = n1564 & n1580;
  assign n1582 = n1542 & n1581;
  assign n1583 = n1528 & n1582;
  assign n1584 = Pdata_11_ & ~n1583;
  assign n1585 = ~Pdata_11_ & n1583;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = n505 & n1586;
  assign n1588 = Poutreg_43_ & n909;
  assign n1589 = Poutreg_35_ & ~Pcount_0_;
  assign n1590 = ~n1588 & ~n1589;
  assign Poutreg_new_35_ = n1587 | ~n1590;
  assign n1592 = Poutreg_42_ & n909;
  assign n1593 = Pdata_43_ & n505;
  assign n1594 = Poutreg_34_ & ~Pcount_0_;
  assign n1595 = ~n1593 & ~n1594;
  assign Poutreg_new_34_ = n1592 | ~n1595;
  assign n1597 = n1283 & ~n1293;
  assign n1598 = n1231 & ~n1274;
  assign n1599 = ~n1283 & ~n1294;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = ~n1597 & n1600;
  assign n1602 = ~n1358 & ~n1601;
  assign n1603 = n1234 & ~n1602;
  assign n1604 = n1231 & n1353;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = n1267 & n1284;
  assign n1607 = ~n1231 & n1246;
  assign n1608 = ~n1282 & n1320;
  assign n1609 = ~n1607 & n1608;
  assign n1610 = ~n1606 & ~n1609;
  assign n1611 = n1312 & n1610;
  assign n1612 = n1291 & n1611;
  assign n1613 = n1350 & n1612;
  assign n1614 = n1605 & n1613;
  assign n1615 = ~Pdata_3_ & ~n1614;
  assign n1616 = Pdata_3_ & n1614;
  assign n1617 = ~n1615 & ~n1616;
  assign n1618 = n505 & ~n1617;
  assign n1619 = Poutreg_41_ & n909;
  assign n1620 = Poutreg_33_ & ~Pcount_0_;
  assign n1621 = ~n1619 & ~n1620;
  assign Poutreg_new_33_ = n1618 | ~n1621;
  assign n1623 = Poutreg_40_ & n909;
  assign n1624 = Poutreg_32_ & ~Pcount_0_;
  assign n1625 = Pdata_35_ & n505;
  assign n1626 = ~n1624 & ~n1625;
  assign Poutreg_new_32_ = n1623 | ~n1626;
  assign n1628 = n1267 & n1287;
  assign n1629 = n1256 & n1269;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1281 & n1350;
  assign n1632 = n1630 & n1631;
  assign n1633 = ~n1240 & n1258;
  assign n1634 = ~n1259 & n1633;
  assign n1635 = ~n1297 & ~n1634;
  assign n1636 = ~n1353 & n1635;
  assign n1637 = ~n1354 & n1636;
  assign n1638 = ~n1231 & ~n1637;
  assign n1639 = n1240 & n1261;
  assign n1640 = n1272 & ~n1283;
  assign n1641 = ~n1342 & ~n1640;
  assign n1642 = ~n1257 & n1641;
  assign n1643 = ~n1639 & n1642;
  assign n1644 = n1231 & ~n1643;
  assign n1645 = ~n1638 & ~n1644;
  assign n1646 = n1317 & n1645;
  assign n1647 = n1632 & n1646;
  assign n1648 = Pdata_28_ & ~n1647;
  assign n1649 = ~Pdata_28_ & n1647;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = n505 & n1650;
  assign n1652 = Poutreg_39_ & n909;
  assign n1653 = Poutreg_31_ & ~Pcount_0_;
  assign n1654 = ~n1652 & ~n1653;
  assign Poutreg_new_31_ = n1651 | ~n1654;
  assign n1656 = Poutreg_38_ & n909;
  assign n1657 = Poutreg_30_ & ~Pcount_0_;
  assign n1658 = Pdata_60_ & n505;
  assign n1659 = ~n1657 & ~n1658;
  assign Poutreg_new_30_ = n1656 | ~n1659;
  assign n1661 = n1170 & n1175;
  assign n1662 = ~n1134 & ~n1144;
  assign n1663 = ~n1111 & n1133;
  assign n1664 = n1662 & n1663;
  assign n1665 = ~n1661 & ~n1664;
  assign n1666 = ~n1123 & ~n1665;
  assign n1667 = n1133 & n1183;
  assign n1668 = ~n1142 & ~n1667;
  assign n1669 = ~n1662 & ~n1668;
  assign n1670 = ~n1114 & n1132;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1666 & n1671;
  assign n1673 = n1167 & n1170;
  assign n1674 = n1123 & n1673;
  assign n1675 = n1126 & n1189;
  assign n1676 = ~n1123 & n1675;
  assign n1677 = ~n1674 & ~n1676;
  assign n1678 = n1168 & n1204;
  assign n1679 = n1178 & n1183;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n1677 & n1680;
  assign n1682 = n1171 & n1205;
  assign n1683 = n1166 & n1662;
  assign n1684 = ~n1184 & n1683;
  assign n1685 = ~n1682 & ~n1684;
  assign n1686 = n1119 & n1127;
  assign n1687 = n1108 & n1686;
  assign n1688 = n1685 & ~n1687;
  assign n1689 = n1201 & n1688;
  assign n1690 = n1192 & n1689;
  assign n1691 = n1681 & n1690;
  assign n1692 = n1672 & n1691;
  assign n1693 = Pdata_20_ & ~n1692;
  assign n1694 = ~Pdata_20_ & n1692;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = n505 & n1695;
  assign n1697 = Poutreg_37_ & n909;
  assign n1698 = Poutreg_29_ & ~Pcount_0_;
  assign n1699 = ~n1697 & ~n1698;
  assign Poutreg_new_29_ = n1696 | ~n1699;
  assign n1701 = Poutreg_36_ & n909;
  assign n1702 = Poutreg_28_ & ~Pcount_0_;
  assign n1703 = Pdata_52_ & n505;
  assign n1704 = ~n1702 & ~n1703;
  assign Poutreg_new_28_ = n1701 | ~n1704;
  assign n1706 = n954 & n1076;
  assign n1707 = n942 & n953;
  assign n1708 = ~n954 & n1707;
  assign n1709 = ~n1706 & ~n1708;
  assign n1710 = ~n962 & ~n1422;
  assign n1711 = ~n932 & n935;
  assign n1712 = n1082 & n1711;
  assign n1713 = n1710 & ~n1712;
  assign n1714 = ~n921 & n938;
  assign n1715 = ~n1713 & n1714;
  assign n1716 = n1709 & ~n1715;
  assign n1717 = n962 & n964;
  assign n1718 = ~n935 & ~n1079;
  assign n1719 = n925 & n1718;
  assign n1720 = ~n1717 & ~n1719;
  assign n1721 = ~n1084 & ~n1720;
  assign n1722 = ~n1063 & n1425;
  assign n1723 = n959 & ~n1722;
  assign n1724 = ~n1721 & n1723;
  assign n1725 = n1716 & n1724;
  assign n1726 = n1421 & n1725;
  assign n1727 = Pdata_12_ & ~n1726;
  assign n1728 = ~Pdata_12_ & n1726;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n505 & n1729;
  assign n1731 = Poutreg_35_ & n909;
  assign n1732 = Poutreg_27_ & ~Pcount_0_;
  assign n1733 = ~n1731 & ~n1732;
  assign Poutreg_new_27_ = n1730 | ~n1733;
  assign n1735 = Poutreg_34_ & n909;
  assign n1736 = Poutreg_26_ & ~Pcount_0_;
  assign n1737 = Pdata_44_ & n505;
  assign n1738 = ~n1736 & ~n1737;
  assign Poutreg_new_26_ = n1735 | ~n1738;
  assign n1740 = n1135 & n1141;
  assign n1741 = ~n1140 & ~n1740;
  assign n1742 = n1123 & ~n1741;
  assign n1743 = n1120 & ~n1126;
  assign n1744 = n1126 & n1161;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = ~n1742 & n1745;
  assign n1747 = n1212 & n1681;
  assign n1748 = n1114 & n1148;
  assign n1749 = ~n1143 & ~n1748;
  assign n1750 = n1193 & ~n1749;
  assign n1751 = n1156 & n1202;
  assign n1752 = ~n1686 & ~n1751;
  assign n1753 = n1131 & n1139;
  assign n1754 = ~n1664 & ~n1753;
  assign n1755 = n1752 & n1754;
  assign n1756 = ~n1750 & n1755;
  assign n1757 = n1191 & n1756;
  assign n1758 = n1747 & n1757;
  assign n1759 = n1746 & n1758;
  assign n1760 = Pdata_4_ & ~n1759;
  assign n1761 = ~Pdata_4_ & n1759;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n505 & n1762;
  assign n1764 = Poutreg_33_ & n909;
  assign n1765 = Poutreg_25_ & ~Pcount_0_;
  assign n1766 = ~n1764 & ~n1765;
  assign Poutreg_new_25_ = n1763 | ~n1766;
  assign n1768 = Poutreg_32_ & n909;
  assign n1769 = Pdata_36_ & n505;
  assign n1770 = Poutreg_24_ & ~Pcount_0_;
  assign n1771 = ~n1769 & ~n1770;
  assign Poutreg_new_24_ = n1768 | ~n1771;
  assign n1773 = Pdata_40_ & ~PC_18_;
  assign n1774 = ~Pdata_40_ & PC_18_;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = Pdata_41_ & ~PC_11_;
  assign n1777 = ~Pdata_41_ & PC_11_;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1775 & n1778;
  assign n1780 = Pdata_39_ & ~PC_22_;
  assign n1781 = ~Pdata_39_ & PC_22_;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = Pdata_43_ & ~PC_25_;
  assign n1784 = ~Pdata_43_ & PC_25_;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = ~n1782 & ~n1785;
  assign n1787 = Pdata_44_ & ~PC_7_;
  assign n1788 = ~Pdata_44_ & PC_7_;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = Pdata_42_ & ~PC_3_;
  assign n1791 = ~Pdata_42_ & PC_3_;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1789 & n1792;
  assign n1794 = n1786 & n1793;
  assign n1795 = n1779 & n1794;
  assign n1796 = n1775 & ~n1782;
  assign n1797 = n1789 & n1792;
  assign n1798 = ~n1785 & n1797;
  assign n1799 = n1796 & n1798;
  assign n1800 = n1789 & ~n1792;
  assign n1801 = n1782 & n1785;
  assign n1802 = n1775 & n1801;
  assign n1803 = n1800 & n1802;
  assign n1804 = ~n1799 & ~n1803;
  assign n1805 = ~n1778 & ~n1804;
  assign n1806 = ~n1789 & ~n1792;
  assign n1807 = ~n1775 & ~n1778;
  assign n1808 = n1806 & n1807;
  assign n1809 = n1801 & n1808;
  assign n1810 = ~n1805 & ~n1809;
  assign n1811 = ~n1795 & n1810;
  assign n1812 = n1782 & ~n1785;
  assign n1813 = n1775 & n1812;
  assign n1814 = n1778 & n1813;
  assign n1815 = ~n1778 & n1785;
  assign n1816 = ~n1775 & ~n1782;
  assign n1817 = n1815 & n1816;
  assign n1818 = ~n1814 & ~n1817;
  assign n1819 = n1800 & ~n1818;
  assign n1820 = ~n1786 & ~n1801;
  assign n1821 = n1779 & n1806;
  assign n1822 = n1820 & n1821;
  assign n1823 = ~n1819 & ~n1822;
  assign n1824 = n1782 & ~n1807;
  assign n1825 = n1785 & ~n1824;
  assign n1826 = ~n1779 & ~n1782;
  assign n1827 = n1797 & ~n1826;
  assign n1828 = n1825 & n1827;
  assign n1829 = n1793 & n1807;
  assign n1830 = n1820 & n1829;
  assign n1831 = ~n1828 & ~n1830;
  assign n1832 = n1823 & n1831;
  assign n1833 = n1775 & ~n1778;
  assign n1834 = n1806 & n1833;
  assign n1835 = n1800 & n1807;
  assign n1836 = ~n1834 & ~n1835;
  assign n1837 = n1786 & ~n1836;
  assign n1838 = n1778 & n1800;
  assign n1839 = ~n1775 & ~n1785;
  assign n1840 = n1838 & n1839;
  assign n1841 = n1782 & n1840;
  assign n1842 = n1793 & n1814;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = ~n1837 & n1843;
  assign n1845 = n1778 & ~n1785;
  assign n1846 = ~n1815 & ~n1845;
  assign n1847 = ~n1775 & ~n1846;
  assign n1848 = n1806 & n1847;
  assign n1849 = n1798 & n1807;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1782 & ~n1850;
  assign n1852 = n1844 & ~n1851;
  assign n1853 = n1826 & ~n1833;
  assign n1854 = n1825 & ~n1853;
  assign n1855 = n1800 & n1854;
  assign n1856 = n1785 & n1793;
  assign n1857 = n1779 & n1782;
  assign n1858 = ~n1833 & ~n1857;
  assign n1859 = n1856 & ~n1858;
  assign n1860 = n1797 & n1802;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = ~n1793 & ~n1800;
  assign n1863 = n1782 & n1833;
  assign n1864 = n1862 & n1863;
  assign n1865 = n1792 & n1845;
  assign n1866 = n1796 & n1865;
  assign n1867 = ~n1864 & ~n1866;
  assign n1868 = n1861 & n1867;
  assign n1869 = ~n1855 & n1868;
  assign n1870 = n1852 & n1869;
  assign n1871 = n1832 & n1870;
  assign n1872 = n1811 & n1871;
  assign n1873 = Pdata_29_ & ~n1872;
  assign n1874 = ~Pdata_29_ & n1872;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = n505 & n1875;
  assign n1877 = Poutreg_31_ & n909;
  assign n1878 = Poutreg_23_ & ~Pcount_0_;
  assign n1879 = ~n1877 & ~n1878;
  assign Poutreg_new_23_ = n1876 | ~n1879;
  assign n1881 = Poutreg_30_ & n909;
  assign n1882 = Poutreg_22_ & ~Pcount_0_;
  assign n1883 = Pdata_61_ & n505;
  assign n1884 = ~n1882 & ~n1883;
  assign Poutreg_new_22_ = n1881 | ~n1884;
  assign n1886 = n1507 & n1533;
  assign n1887 = n1513 & n1530;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = ~n1549 & ~n1572;
  assign n1890 = n1492 & ~n1889;
  assign n1891 = n1554 & ~n1890;
  assign n1892 = n1888 & n1891;
  assign n1893 = n1542 & n1892;
  assign n1894 = n1504 & n1560;
  assign n1895 = ~n1555 & ~n1894;
  assign n1896 = ~n1510 & ~n1895;
  assign n1897 = ~n1488 & n1495;
  assign n1898 = ~n1491 & n1504;
  assign n1899 = n1897 & ~n1898;
  assign n1900 = ~n1532 & ~n1899;
  assign n1901 = n1498 & n1507;
  assign n1902 = ~n1900 & n1901;
  assign n1903 = n1499 & n1524;
  assign n1904 = ~n1902 & ~n1903;
  assign n1905 = ~n1896 & n1904;
  assign n1906 = ~n1491 & n1518;
  assign n1907 = ~n1546 & ~n1906;
  assign n1908 = n1510 & ~n1907;
  assign n1909 = n1492 & n1571;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1905 & n1910;
  assign n1912 = n1579 & n1911;
  assign n1913 = n1893 & n1912;
  assign n1914 = Pdata_21_ & ~n1913;
  assign n1915 = ~Pdata_21_ & n1913;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n505 & n1916;
  assign n1918 = Poutreg_29_ & n909;
  assign n1919 = Poutreg_21_ & ~Pcount_0_;
  assign n1920 = ~n1918 & ~n1919;
  assign Poutreg_new_21_ = n1917 | ~n1920;
  assign n1922 = Poutreg_28_ & n909;
  assign n1923 = Poutreg_20_ & ~Pcount_0_;
  assign n1924 = Pdata_53_ & n505;
  assign n1925 = ~n1923 & ~n1924;
  assign Poutreg_new_20_ = n1922 | ~n1925;
  assign n1927 = n518 & ~n528;
  assign n1928 = n511 & ~n524;
  assign n1929 = ~n557 & ~n1928;
  assign n1930 = ~n1927 & ~n1929;
  assign n1931 = n518 & n1929;
  assign n1932 = n508 & ~n1931;
  assign n1933 = ~n1930 & n1932;
  assign n1934 = n548 & n1401;
  assign n1935 = ~n573 & ~n1934;
  assign n1936 = ~n1933 & n1935;
  assign n1937 = ~n544 & n1936;
  assign n1938 = n515 & ~n1937;
  assign n1939 = ~n518 & ~n537;
  assign n1940 = n579 & ~n1927;
  assign n1941 = ~n518 & n567;
  assign n1942 = n1940 & ~n1941;
  assign n1943 = ~n1939 & n1942;
  assign n1944 = ~n589 & ~n1943;
  assign n1945 = ~n515 & ~n1944;
  assign n1946 = n594 & n1400;
  assign n1947 = ~n1945 & n1946;
  assign n1948 = n561 & n1393;
  assign n1949 = n565 & ~n1948;
  assign n1950 = n1947 & n1949;
  assign n1951 = ~n1938 & n1950;
  assign n1952 = Pdata_13_ & ~n1951;
  assign n1953 = ~Pdata_13_ & n1951;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = n505 & n1954;
  assign n1956 = Poutreg_27_ & n909;
  assign n1957 = Poutreg_19_ & ~Pcount_0_;
  assign n1958 = ~n1956 & ~n1957;
  assign Poutreg_new_19_ = n1955 | ~n1958;
  assign n1960 = Poutreg_26_ & n909;
  assign n1961 = Pdata_45_ & n505;
  assign n1962 = Poutreg_18_ & ~Pcount_0_;
  assign n1963 = ~n1961 & ~n1962;
  assign Poutreg_new_18_ = n1960 | ~n1963;
  assign n1965 = n1797 & n1817;
  assign n1966 = n1793 & n1802;
  assign n1967 = n1785 & n1862;
  assign n1968 = n1796 & n1967;
  assign n1969 = ~n1966 & ~n1968;
  assign n1970 = n1778 & ~n1969;
  assign n1971 = n1798 & n1857;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = n1811 & n1972;
  assign n1974 = n1844 & n1973;
  assign n1975 = ~n1965 & n1974;
  assign n1976 = n1796 & n1856;
  assign n1977 = ~n1775 & n1862;
  assign n1978 = ~n1820 & n1977;
  assign n1979 = ~n1976 & ~n1978;
  assign n1980 = n1806 & n1813;
  assign n1981 = n1778 & ~n1980;
  assign n1982 = n1979 & n1981;
  assign n1983 = n1789 & n1813;
  assign n1984 = ~n1966 & ~n1983;
  assign n1985 = ~n1794 & n1984;
  assign n1986 = ~n1778 & n1985;
  assign n1987 = ~n1982 & ~n1986;
  assign n1988 = n1778 & n1802;
  assign n1989 = n1796 & ~n1846;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = n1800 & ~n1990;
  assign n1992 = n1808 & n1812;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n1987 & n1993;
  assign n1995 = n1831 & n1994;
  assign n1996 = n1975 & n1995;
  assign n1997 = Pdata_5_ & ~n1996;
  assign n1998 = ~Pdata_5_ & n1996;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = n505 & n1999;
  assign n2001 = Poutreg_25_ & n909;
  assign n2002 = Poutreg_17_ & ~Pcount_0_;
  assign n2003 = ~n2001 & ~n2002;
  assign Poutreg_new_17_ = n2000 | ~n2003;
  assign n2005 = Poutreg_24_ & n909;
  assign n2006 = Poutreg_16_ & ~Pcount_0_;
  assign n2007 = Pdata_37_ & n505;
  assign n2008 = ~n2006 & ~n2007;
  assign Poutreg_new_16_ = n2005 | ~n2008;
  assign n2010 = ~n614 & n653;
  assign n2011 = ~n695 & ~n697;
  assign n2012 = ~n2010 & n2011;
  assign n2013 = n657 & ~n2012;
  assign n2014 = ~n653 & ~n694;
  assign n2015 = n654 & n2014;
  assign n2016 = ~n633 & ~n2015;
  assign n2017 = ~n630 & n706;
  assign n2018 = n753 & ~n2017;
  assign n2019 = n2016 & n2018;
  assign n2020 = ~n2013 & n2019;
  assign n2021 = n676 & n2020;
  assign n2022 = Pdata_30_ & ~n2021;
  assign n2023 = ~Pdata_30_ & n2021;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = n505 & n2024;
  assign n2026 = Poutreg_23_ & n909;
  assign n2027 = Poutreg_15_ & ~Pcount_0_;
  assign n2028 = ~n2026 & ~n2027;
  assign Poutreg_new_15_ = n2025 | ~n2028;
  assign n2030 = Poutreg_22_ & n909;
  assign n2031 = Poutreg_14_ & ~Pcount_0_;
  assign n2032 = Pdata_62_ & n505;
  assign n2033 = ~n2031 & ~n2032;
  assign Poutreg_new_14_ = n2030 | ~n2033;
  assign n2035 = n617 & ~n630;
  assign n2036 = ~n699 & ~n2035;
  assign n2037 = ~n624 & n659;
  assign n2038 = n684 & n2035;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~n2036 & ~n2039;
  assign n2041 = ~n632 & ~n734;
  assign n2042 = n624 & n734;
  assign n2043 = ~n728 & ~n2042;
  assign n2044 = ~n2041 & ~n2043;
  assign n2045 = n664 & ~n2044;
  assign n2046 = ~n2040 & n2045;
  assign n2047 = n614 & n730;
  assign n2048 = ~n747 & ~n2047;
  assign n2049 = n712 & ~n2048;
  assign n2050 = n675 & ~n2049;
  assign n2051 = n754 & n2050;
  assign n2052 = n2046 & n2051;
  assign n2053 = Pdata_22_ & ~n2052;
  assign n2054 = ~Pdata_22_ & n2052;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = n505 & n2055;
  assign n2057 = Poutreg_21_ & n909;
  assign n2058 = Poutreg_13_ & ~Pcount_0_;
  assign n2059 = ~n2057 & ~n2058;
  assign Poutreg_new_13_ = n2056 | ~n2059;
  assign n2061 = Poutreg_20_ & n909;
  assign n2062 = Poutreg_12_ & ~Pcount_0_;
  assign n2063 = Pdata_54_ & n505;
  assign n2064 = ~n2062 & ~n2063;
  assign Poutreg_new_12_ = n2061 | ~n2064;
  assign n2066 = n1108 & ~n1126;
  assign n2067 = ~n1148 & ~n2066;
  assign n2068 = n1175 & ~n2067;
  assign n2069 = ~n1172 & ~n2068;
  assign n2070 = ~n1120 & n2069;
  assign n2071 = ~n1123 & ~n2070;
  assign n2072 = n1117 & n1663;
  assign n2073 = ~n1185 & ~n2072;
  assign n2074 = n1130 & n1166;
  assign n2075 = n1146 & ~n2074;
  assign n2076 = n2073 & n2075;
  assign n2077 = n1123 & ~n2076;
  assign n2078 = ~n1119 & ~n2072;
  assign n2079 = n1126 & ~n2078;
  assign n2080 = ~n2077 & ~n2079;
  assign n2081 = n1181 & n1747;
  assign n2082 = n2080 & n2081;
  assign n2083 = ~n2071 & n2082;
  assign n2084 = Pdata_14_ & ~n2083;
  assign n2085 = ~Pdata_14_ & n2083;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n505 & n2086;
  assign n2088 = Poutreg_19_ & n909;
  assign n2089 = Poutreg_11_ & ~Pcount_0_;
  assign n2090 = ~n2088 & ~n2089;
  assign Poutreg_new_11_ = n2087 | ~n2090;
  assign n2092 = Poutreg_18_ & n909;
  assign n2093 = Poutreg_10_ & ~Pcount_0_;
  assign n2094 = Pdata_46_ & n505;
  assign n2095 = ~n2093 & ~n2094;
  assign Poutreg_new_10_ = n2092 | ~n2095;
  assign n2097 = n1504 & n1906;
  assign n2098 = ~n1575 & ~n2097;
  assign n2099 = ~n1517 & ~n2098;
  assign n2100 = n1513 & n1524;
  assign n2101 = n1517 & n1539;
  assign n2102 = ~n1495 & n1515;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~n2100 & n2103;
  assign n2105 = n1570 & n2104;
  assign n2106 = n1488 & ~n1498;
  assign n2107 = ~n1495 & n2106;
  assign n2108 = ~n1510 & n2107;
  assign n2109 = ~n1571 & ~n2108;
  assign n2110 = n1491 & ~n2109;
  assign n2111 = n1504 & n1557;
  assign n2112 = ~n1522 & ~n2111;
  assign n2113 = n1507 & ~n2112;
  assign n2114 = ~n2110 & ~n2113;
  assign n2115 = n2105 & n2114;
  assign n2116 = ~n2099 & n2115;
  assign n2117 = n1893 & n2116;
  assign n2118 = Pdata_6_ & ~n2117;
  assign n2119 = ~Pdata_6_ & n2117;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = n505 & n2120;
  assign n2122 = Poutreg_17_ & n909;
  assign n2123 = Poutreg_9_ & ~Pcount_0_;
  assign n2124 = ~n2122 & ~n2123;
  assign Poutreg_new_9_ = n2121 | ~n2124;
  assign n2126 = Poutreg_16_ & n909;
  assign n2127 = Pdata_38_ & n505;
  assign n2128 = Poutreg_8_ & ~Pcount_0_;
  assign n2129 = ~n2127 & ~n2128;
  assign Poutreg_new_8_ = n2126 | ~n2129;
  assign n2131 = ~n1491 & n1495;
  assign n2132 = ~n1504 & ~n2131;
  assign n2133 = ~n1521 & n2106;
  assign n2134 = ~n2132 & n2133;
  assign n2135 = ~n1523 & ~n2134;
  assign n2136 = ~n2111 & n2135;
  assign n2137 = ~n1507 & ~n2136;
  assign n2138 = n1517 & n1529;
  assign n2139 = ~n1515 & ~n1524;
  assign n2140 = ~n2138 & n2139;
  assign n2141 = n1500 & ~n2140;
  assign n2142 = ~n2137 & ~n2141;
  assign n2143 = n1495 & n1543;
  assign n2144 = ~n1539 & ~n2143;
  assign n2145 = n1509 & ~n2144;
  assign n2146 = n1511 & n1514;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = n1580 & n2147;
  assign n2149 = n1892 & n2148;
  assign n2150 = n2142 & n2149;
  assign n2151 = ~Pdata_31_ & ~n2150;
  assign n2152 = Pdata_31_ & n2150;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = n505 & ~n2153;
  assign n2155 = Poutreg_15_ & n909;
  assign n2156 = Poutreg_7_ & ~Pcount_0_;
  assign n2157 = ~n2155 & ~n2156;
  assign Poutreg_new_7_ = n2154 | ~n2157;
  assign n2159 = Poutreg_14_ & n909;
  assign n2160 = Poutreg_6_ & ~Pcount_0_;
  assign n2161 = Pdata_63_ & n505;
  assign n2162 = ~n2160 & ~n2161;
  assign Poutreg_new_6_ = n2159 | ~n2162;
  assign n2164 = ~n1786 & ~n1847;
  assign n2165 = n1793 & ~n2164;
  assign n2166 = ~n1816 & n2165;
  assign n2167 = n1789 & n1988;
  assign n2168 = n1812 & n1835;
  assign n2169 = ~n1980 & ~n2168;
  assign n2170 = ~n2167 & n2169;
  assign n2171 = ~n1778 & n1839;
  assign n2172 = n1775 & n1815;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = ~n1782 & n1862;
  assign n2175 = ~n2173 & n2174;
  assign n2176 = ~n1820 & n1838;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = n2170 & n2177;
  assign n2179 = ~n2166 & n2178;
  assign n2180 = n1832 & n2179;
  assign n2181 = n1973 & n2180;
  assign n2182 = Pdata_23_ & ~n2181;
  assign n2183 = ~Pdata_23_ & n2181;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = n505 & n2184;
  assign n2186 = Poutreg_13_ & n909;
  assign n2187 = Poutreg_5_ & ~Pcount_0_;
  assign n2188 = ~n2186 & ~n2187;
  assign Poutreg_new_5_ = n2185 | ~n2188;
  assign n2190 = Poutreg_12_ & n909;
  assign n2191 = Pdata_55_ & n505;
  assign n2192 = Poutreg_4_ & ~Pcount_0_;
  assign n2193 = ~n2191 & ~n2192;
  assign Poutreg_new_4_ = n2190 | ~n2193;
  assign n2195 = ~n1789 & n2171;
  assign n2196 = ~n1840 & ~n2195;
  assign n2197 = ~n1782 & ~n2196;
  assign n2198 = n1785 & n1838;
  assign n2199 = ~n1798 & ~n2198;
  assign n2200 = n1796 & ~n2199;
  assign n2201 = ~n2197 & ~n2200;
  assign n2202 = n1793 & n1854;
  assign n2203 = n1782 & n1849;
  assign n2204 = n1785 & n1857;
  assign n2205 = ~n1792 & n2204;
  assign n2206 = ~n2203 & ~n2205;
  assign n2207 = ~n2202 & n2206;
  assign n2208 = ~n1785 & ~n1862;
  assign n2209 = ~n1967 & ~n2208;
  assign n2210 = n1863 & ~n2209;
  assign n2211 = n1823 & ~n2210;
  assign n2212 = n2207 & n2211;
  assign n2213 = n1975 & n2212;
  assign n2214 = n2201 & n2213;
  assign n2215 = Pdata_15_ & ~n2214;
  assign n2216 = ~Pdata_15_ & n2214;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n505 & n2217;
  assign n2219 = Poutreg_11_ & n909;
  assign n2220 = Poutreg_3_ & ~Pcount_0_;
  assign n2221 = ~n2219 & ~n2220;
  assign Poutreg_new_3_ = n2218 | ~n2221;
  assign n2223 = Poutreg_10_ & n909;
  assign n2224 = Poutreg_2_ & ~Pcount_0_;
  assign n2225 = Pdata_47_ & n505;
  assign n2226 = ~n2224 & ~n2225;
  assign Poutreg_new_2_ = n2223 | ~n2226;
  assign n2228 = ~n526 & ~n547;
  assign n2229 = n1380 & ~n2228;
  assign n2230 = ~n518 & ~n567;
  assign n2231 = n580 & n2230;
  assign n2232 = n515 & n555;
  assign n2233 = ~n1383 & ~n2232;
  assign n2234 = n542 & n2233;
  assign n2235 = ~n508 & ~n529;
  assign n2236 = n512 & ~n557;
  assign n2237 = ~n1939 & ~n2236;
  assign n2238 = ~n2235 & n2237;
  assign n2239 = ~n2234 & n2238;
  assign n2240 = n562 & n567;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = ~n2231 & n2241;
  assign n2243 = ~n2229 & n2242;
  assign n2244 = n552 & n2243;
  assign n2245 = n1946 & n2244;
  assign n2246 = Pdata_7_ & ~n2245;
  assign n2247 = ~Pdata_7_ & n2245;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = n505 & n2248;
  assign n2250 = Poutreg_9_ & n909;
  assign n2251 = Poutreg_1_ & ~Pcount_0_;
  assign n2252 = ~n2250 & ~n2251;
  assign Poutreg_new_1_ = n2249 | ~n2252;
  assign n2254 = Poutreg_8_ & n909;
  assign n2255 = Poutreg_0_ & ~Pcount_0_;
  assign n2256 = Pdata_39_ & n505;
  assign n2257 = ~n2255 & ~n2256;
  assign Poutreg_new_0_ = n2254 | ~n2257;
  assign n2259 = Pinreg_55_ & ~Pcount_0_;
  assign n2260 = Pinreg_47_ & n909;
  assign Pinreg_new_55_ = n2259 | n2260;
  assign n2262 = Pinreg_54_ & ~Pcount_0_;
  assign n2263 = Pinreg_46_ & n909;
  assign Pinreg_new_54_ = n2262 | n2263;
  assign n2265 = Pinreg_53_ & ~Pcount_0_;
  assign n2266 = Pinreg_45_ & n909;
  assign Pinreg_new_53_ = n2265 | n2266;
  assign n2268 = Pinreg_52_ & ~Pcount_0_;
  assign n2269 = Pinreg_44_ & n909;
  assign Pinreg_new_52_ = n2268 | n2269;
  assign n2271 = Pinreg_51_ & ~Pcount_0_;
  assign n2272 = Pinreg_43_ & n909;
  assign Pinreg_new_51_ = n2271 | n2272;
  assign n2274 = Pinreg_50_ & ~Pcount_0_;
  assign n2275 = Pinreg_42_ & n909;
  assign Pinreg_new_50_ = n2274 | n2275;
  assign n2277 = Pinreg_49_ & ~Pcount_0_;
  assign n2278 = Pinreg_41_ & n909;
  assign Pinreg_new_49_ = n2277 | n2278;
  assign n2280 = Pinreg_48_ & ~Pcount_0_;
  assign n2281 = Pinreg_40_ & n909;
  assign Pinreg_new_48_ = n2280 | n2281;
  assign n2283 = Pinreg_47_ & ~Pcount_0_;
  assign n2284 = Pinreg_39_ & n909;
  assign Pinreg_new_47_ = n2283 | n2284;
  assign n2286 = Pinreg_46_ & ~Pcount_0_;
  assign n2287 = Pinreg_38_ & n909;
  assign Pinreg_new_46_ = n2286 | n2287;
  assign n2289 = Pinreg_45_ & ~Pcount_0_;
  assign n2290 = Pinreg_37_ & n909;
  assign Pinreg_new_45_ = n2289 | n2290;
  assign n2292 = Pinreg_44_ & ~Pcount_0_;
  assign n2293 = Pinreg_36_ & n909;
  assign Pinreg_new_44_ = n2292 | n2293;
  assign n2295 = Pinreg_43_ & ~Pcount_0_;
  assign n2296 = Pinreg_35_ & n909;
  assign Pinreg_new_43_ = n2295 | n2296;
  assign n2298 = Pinreg_42_ & ~Pcount_0_;
  assign n2299 = Pinreg_34_ & n909;
  assign Pinreg_new_42_ = n2298 | n2299;
  assign n2301 = Pinreg_41_ & ~Pcount_0_;
  assign n2302 = Pinreg_33_ & n909;
  assign Pinreg_new_41_ = n2301 | n2302;
  assign n2304 = Pinreg_40_ & ~Pcount_0_;
  assign n2305 = Pinreg_32_ & n909;
  assign Pinreg_new_40_ = n2304 | n2305;
  assign n2307 = Pinreg_39_ & ~Pcount_0_;
  assign n2308 = Pinreg_31_ & n909;
  assign Pinreg_new_39_ = n2307 | n2308;
  assign n2310 = Pinreg_38_ & ~Pcount_0_;
  assign n2311 = Pinreg_30_ & n909;
  assign Pinreg_new_38_ = n2310 | n2311;
  assign n2313 = Pinreg_37_ & ~Pcount_0_;
  assign n2314 = Pinreg_29_ & n909;
  assign Pinreg_new_37_ = n2313 | n2314;
  assign n2316 = Pinreg_36_ & ~Pcount_0_;
  assign n2317 = Pinreg_28_ & n909;
  assign Pinreg_new_36_ = n2316 | n2317;
  assign n2319 = Pinreg_35_ & ~Pcount_0_;
  assign n2320 = Pinreg_27_ & n909;
  assign Pinreg_new_35_ = n2319 | n2320;
  assign n2322 = Pinreg_34_ & ~Pcount_0_;
  assign n2323 = Pinreg_26_ & n909;
  assign Pinreg_new_34_ = n2322 | n2323;
  assign n2325 = Pinreg_33_ & ~Pcount_0_;
  assign n2326 = Pinreg_25_ & n909;
  assign Pinreg_new_33_ = n2325 | n2326;
  assign n2328 = Pinreg_32_ & ~Pcount_0_;
  assign n2329 = Pinreg_24_ & n909;
  assign Pinreg_new_32_ = n2328 | n2329;
  assign n2331 = Pinreg_31_ & ~Pcount_0_;
  assign n2332 = Pinreg_23_ & n909;
  assign Pinreg_new_31_ = n2331 | n2332;
  assign n2334 = Pinreg_30_ & ~Pcount_0_;
  assign n2335 = Pinreg_22_ & n909;
  assign Pinreg_new_30_ = n2334 | n2335;
  assign n2337 = Pinreg_29_ & ~Pcount_0_;
  assign n2338 = Pinreg_21_ & n909;
  assign Pinreg_new_29_ = n2337 | n2338;
  assign n2340 = Pinreg_28_ & ~Pcount_0_;
  assign n2341 = Pinreg_20_ & n909;
  assign Pinreg_new_28_ = n2340 | n2341;
  assign n2343 = Pinreg_27_ & ~Pcount_0_;
  assign n2344 = Pinreg_19_ & n909;
  assign Pinreg_new_27_ = n2343 | n2344;
  assign n2346 = Pinreg_26_ & ~Pcount_0_;
  assign n2347 = Pinreg_18_ & n909;
  assign Pinreg_new_26_ = n2346 | n2347;
  assign n2349 = Pinreg_25_ & ~Pcount_0_;
  assign n2350 = Pinreg_17_ & n909;
  assign Pinreg_new_25_ = n2349 | n2350;
  assign n2352 = Pinreg_24_ & ~Pcount_0_;
  assign n2353 = Pinreg_16_ & n909;
  assign Pinreg_new_24_ = n2352 | n2353;
  assign n2355 = Pinreg_23_ & ~Pcount_0_;
  assign n2356 = Pinreg_15_ & n909;
  assign Pinreg_new_23_ = n2355 | n2356;
  assign n2358 = Pinreg_22_ & ~Pcount_0_;
  assign n2359 = Pinreg_14_ & n909;
  assign Pinreg_new_22_ = n2358 | n2359;
  assign n2361 = Pinreg_21_ & ~Pcount_0_;
  assign n2362 = Pinreg_13_ & n909;
  assign Pinreg_new_21_ = n2361 | n2362;
  assign n2364 = Pinreg_20_ & ~Pcount_0_;
  assign n2365 = Pinreg_12_ & n909;
  assign Pinreg_new_20_ = n2364 | n2365;
  assign n2367 = Pinreg_19_ & ~Pcount_0_;
  assign n2368 = Pinreg_11_ & n909;
  assign Pinreg_new_19_ = n2367 | n2368;
  assign n2370 = Pinreg_18_ & ~Pcount_0_;
  assign n2371 = Pinreg_10_ & n909;
  assign Pinreg_new_18_ = n2370 | n2371;
  assign n2373 = Pinreg_17_ & ~Pcount_0_;
  assign n2374 = Pinreg_9_ & n909;
  assign Pinreg_new_17_ = n2373 | n2374;
  assign n2376 = Pinreg_16_ & ~Pcount_0_;
  assign n2377 = Pinreg_8_ & n909;
  assign Pinreg_new_16_ = n2376 | n2377;
  assign n2379 = Pinreg_15_ & ~Pcount_0_;
  assign n2380 = Pinreg_7_ & n909;
  assign Pinreg_new_15_ = n2379 | n2380;
  assign n2382 = Pinreg_14_ & ~Pcount_0_;
  assign n2383 = Pinreg_6_ & n909;
  assign Pinreg_new_14_ = n2382 | n2383;
  assign n2385 = Pinreg_13_ & ~Pcount_0_;
  assign n2386 = Pinreg_5_ & n909;
  assign Pinreg_new_13_ = n2385 | n2386;
  assign n2388 = Pinreg_12_ & ~Pcount_0_;
  assign n2389 = Pinreg_4_ & n909;
  assign Pinreg_new_12_ = n2388 | n2389;
  assign n2391 = Pinreg_11_ & ~Pcount_0_;
  assign n2392 = Pinreg_3_ & n909;
  assign Pinreg_new_11_ = n2391 | n2392;
  assign n2394 = Pinreg_10_ & ~Pcount_0_;
  assign n2395 = Pinreg_2_ & n909;
  assign Pinreg_new_10_ = n2394 | n2395;
  assign n2397 = Pinreg_9_ & ~Pcount_0_;
  assign n2398 = Pinreg_1_ & n909;
  assign Pinreg_new_9_ = n2397 | n2398;
  assign n2400 = Pinreg_8_ & ~Pcount_0_;
  assign n2401 = Pinreg_0_ & n909;
  assign Pinreg_new_8_ = n2400 | n2401;
  assign n2403 = Pinreg_7_ & ~Pcount_0_;
  assign n2404 = Pdata_in_7_ & n909;
  assign Pinreg_new_7_ = n2403 | n2404;
  assign n2406 = Pinreg_6_ & ~Pcount_0_;
  assign n2407 = Pdata_in_6_ & n909;
  assign Pinreg_new_6_ = n2406 | n2407;
  assign n2409 = Pinreg_5_ & ~Pcount_0_;
  assign n2410 = Pdata_in_5_ & n909;
  assign Pinreg_new_5_ = n2409 | n2410;
  assign n2412 = Pinreg_4_ & ~Pcount_0_;
  assign n2413 = Pdata_in_4_ & n909;
  assign Pinreg_new_4_ = n2412 | n2413;
  assign n2415 = Pinreg_3_ & ~Pcount_0_;
  assign n2416 = Pdata_in_3_ & n909;
  assign Pinreg_new_3_ = n2415 | n2416;
  assign n2418 = Pinreg_2_ & ~Pcount_0_;
  assign n2419 = Pdata_in_2_ & n909;
  assign Pinreg_new_2_ = n2418 | n2419;
  assign n2421 = Pinreg_1_ & ~Pcount_0_;
  assign n2422 = Pdata_in_1_ & n909;
  assign Pinreg_new_1_ = n2421 | n2422;
  assign n2424 = Pinreg_0_ & ~Pcount_0_;
  assign n2425 = Pdata_in_0_ & n909;
  assign Pinreg_new_0_ = n2424 | n2425;
  assign n2427 = Pencrypt_0_ & n505;
  assign n2428 = Pencrypt_mode_0_ & ~n505;
  assign Pencrypt_mode_new_0_ = n2427 | n2428;
  assign n2430 = ~Pdata_in_6_ & n505;
  assign n2431 = ~n505 & n2153;
  assign Pdata_new_63_ = ~n2430 & ~n2431;
  assign n2433 = ~Pinreg_6_ & n505;
  assign n2434 = ~n505 & ~n2024;
  assign Pdata_new_62_ = ~n2433 & ~n2434;
  assign n2436 = ~Pinreg_14_ & n505;
  assign n2437 = ~n505 & ~n1875;
  assign Pdata_new_61_ = ~n2436 & ~n2437;
  assign n2439 = ~Pinreg_22_ & n505;
  assign n2440 = ~n505 & ~n1650;
  assign Pdata_new_60_ = ~n2439 & ~n2440;
  assign n2442 = ~Pinreg_30_ & n505;
  assign n2443 = ~n505 & ~n1442;
  assign Pdata_new_59_ = ~n2442 & ~n2443;
  assign n2445 = ~Pinreg_38_ & n505;
  assign n2446 = ~n505 & ~n1218;
  assign Pdata_new_58_ = ~n2445 & ~n2446;
  assign n2448 = ~Pinreg_46_ & n505;
  assign n2449 = ~n505 & ~n907;
  assign Pdata_new_57_ = ~n2448 & ~n2449;
  assign n2451 = ~Pinreg_54_ & n505;
  assign n2452 = ~n505 & ~n605;
  assign Pdata_new_56_ = ~n2451 & ~n2452;
  assign n2454 = ~Pdata_in_4_ & n505;
  assign n2455 = ~n505 & ~n2184;
  assign Pdata_new_55_ = ~n2454 & ~n2455;
  assign n2457 = ~Pinreg_4_ & n505;
  assign n2458 = ~n505 & ~n2055;
  assign Pdata_new_54_ = ~n2457 & ~n2458;
  assign n2460 = ~Pinreg_12_ & n505;
  assign n2461 = ~n505 & ~n1916;
  assign Pdata_new_53_ = ~n2460 & ~n2461;
  assign n2463 = ~Pinreg_20_ & n505;
  assign n2464 = ~n505 & ~n1695;
  assign Pdata_new_52_ = ~n2463 & ~n2464;
  assign n2466 = ~Pinreg_28_ & n505;
  assign n2467 = ~n505 & ~n1475;
  assign Pdata_new_51_ = ~n2466 & ~n2467;
  assign n2469 = ~Pinreg_36_ & n505;
  assign n2470 = ~n505 & ~n1329;
  assign Pdata_new_50_ = ~n2469 & ~n2470;
  assign n2472 = ~Pinreg_44_ & n505;
  assign n2473 = ~n505 & ~n1014;
  assign Pdata_new_49_ = ~n2472 & ~n2473;
  assign n2475 = ~Pinreg_52_ & n505;
  assign n2476 = ~n505 & ~n721;
  assign Pdata_new_48_ = ~n2475 & ~n2476;
  assign n2478 = ~Pdata_in_2_ & n505;
  assign n2479 = ~n505 & ~n2217;
  assign Pdata_new_47_ = ~n2478 & ~n2479;
  assign n2481 = ~Pinreg_2_ & n505;
  assign n2482 = ~n505 & ~n2086;
  assign Pdata_new_46_ = ~n2481 & ~n2482;
  assign n2484 = ~Pinreg_10_ & n505;
  assign n2485 = ~n505 & ~n1954;
  assign Pdata_new_45_ = ~n2484 & ~n2485;
  assign n2487 = ~Pinreg_18_ & n505;
  assign n2488 = ~n505 & ~n1729;
  assign Pdata_new_44_ = ~n2487 & ~n2488;
  assign n2490 = ~Pinreg_26_ & n505;
  assign n2491 = ~n505 & ~n1586;
  assign Pdata_new_43_ = ~n2490 & ~n2491;
  assign n2493 = ~Pinreg_34_ & n505;
  assign n2494 = ~n505 & ~n1369;
  assign Pdata_new_42_ = ~n2493 & ~n2494;
  assign n2496 = ~Pinreg_42_ & n505;
  assign n2497 = ~n505 & ~n1049;
  assign Pdata_new_41_ = ~n2496 & ~n2497;
  assign n2499 = ~Pinreg_50_ & n505;
  assign n2500 = ~n505 & ~n760;
  assign Pdata_new_40_ = ~n2499 & ~n2500;
  assign n2502 = ~Pdata_in_0_ & n505;
  assign n2503 = ~n505 & ~n2248;
  assign Pdata_new_39_ = ~n2502 & ~n2503;
  assign n2505 = ~Pinreg_0_ & n505;
  assign n2506 = ~n505 & ~n2120;
  assign Pdata_new_38_ = ~n2505 & ~n2506;
  assign n2508 = Pinreg_8_ & n505;
  assign n2509 = ~n505 & n1999;
  assign Pdata_new_37_ = n2508 | n2509;
  assign n2511 = ~Pinreg_16_ & n505;
  assign n2512 = ~n505 & ~n1762;
  assign Pdata_new_36_ = ~n2511 & ~n2512;
  assign n2514 = ~Pinreg_24_ & n505;
  assign n2515 = ~n505 & n1617;
  assign Pdata_new_35_ = ~n2514 & ~n2515;
  assign n2517 = Pinreg_32_ & n505;
  assign n2518 = ~n505 & ~n1410;
  assign Pdata_new_34_ = n2517 | n2518;
  assign n2520 = ~Pinreg_40_ & n505;
  assign n2521 = ~n505 & n1095;
  assign Pdata_new_33_ = ~n2520 & ~n2521;
  assign n2523 = ~Pinreg_48_ & n505;
  assign n2524 = ~n505 & ~n870;
  assign Pdata_new_32_ = ~n2523 & ~n2524;
  assign n2526 = Pdata_in_7_ & n505;
  assign n2527 = Pdata_63_ & ~n505;
  assign Pdata_new_31_ = n2526 | n2527;
  assign n2529 = Pinreg_7_ & n505;
  assign n2530 = Pdata_62_ & ~n505;
  assign Pdata_new_30_ = n2529 | n2530;
  assign n2532 = Pinreg_15_ & n505;
  assign n2533 = Pdata_61_ & ~n505;
  assign Pdata_new_29_ = n2532 | n2533;
  assign n2535 = Pinreg_23_ & n505;
  assign n2536 = Pdata_60_ & ~n505;
  assign Pdata_new_28_ = n2535 | n2536;
  assign n2538 = Pinreg_31_ & n505;
  assign n2539 = Pdata_59_ & ~n505;
  assign Pdata_new_27_ = n2538 | n2539;
  assign n2541 = Pinreg_39_ & n505;
  assign n2542 = Pdata_58_ & ~n505;
  assign Pdata_new_26_ = n2541 | n2542;
  assign n2544 = Pinreg_47_ & n505;
  assign n2545 = Pdata_57_ & ~n505;
  assign Pdata_new_25_ = n2544 | n2545;
  assign n2547 = Pinreg_55_ & n505;
  assign n2548 = Pdata_56_ & ~n505;
  assign Pdata_new_24_ = n2547 | n2548;
  assign n2550 = Pdata_in_5_ & n505;
  assign n2551 = Pdata_55_ & ~n505;
  assign Pdata_new_23_ = n2550 | n2551;
  assign n2553 = Pinreg_5_ & n505;
  assign n2554 = Pdata_54_ & ~n505;
  assign Pdata_new_22_ = n2553 | n2554;
  assign n2556 = Pinreg_13_ & n505;
  assign n2557 = Pdata_53_ & ~n505;
  assign Pdata_new_21_ = n2556 | n2557;
  assign n2559 = Pinreg_21_ & n505;
  assign n2560 = Pdata_52_ & ~n505;
  assign Pdata_new_20_ = n2559 | n2560;
  assign n2562 = Pinreg_29_ & n505;
  assign n2563 = Pdata_51_ & ~n505;
  assign Pdata_new_19_ = n2562 | n2563;
  assign n2565 = Pinreg_37_ & n505;
  assign n2566 = Pdata_50_ & ~n505;
  assign Pdata_new_18_ = n2565 | n2566;
  assign n2568 = Pinreg_45_ & n505;
  assign n2569 = Pdata_49_ & ~n505;
  assign Pdata_new_17_ = n2568 | n2569;
  assign n2571 = Pinreg_53_ & n505;
  assign n2572 = Pdata_48_ & ~n505;
  assign Pdata_new_16_ = n2571 | n2572;
  assign n2574 = Pdata_in_3_ & n505;
  assign n2575 = Pdata_47_ & ~n505;
  assign Pdata_new_15_ = n2574 | n2575;
  assign n2577 = Pinreg_3_ & n505;
  assign n2578 = Pdata_46_ & ~n505;
  assign Pdata_new_14_ = n2577 | n2578;
  assign n2580 = Pinreg_11_ & n505;
  assign n2581 = Pdata_45_ & ~n505;
  assign Pdata_new_13_ = n2580 | n2581;
  assign n2583 = Pinreg_19_ & n505;
  assign n2584 = Pdata_44_ & ~n505;
  assign Pdata_new_12_ = n2583 | n2584;
  assign n2586 = Pinreg_27_ & n505;
  assign n2587 = Pdata_43_ & ~n505;
  assign Pdata_new_11_ = n2586 | n2587;
  assign n2589 = Pinreg_35_ & n505;
  assign n2590 = Pdata_42_ & ~n505;
  assign Pdata_new_10_ = n2589 | n2590;
  assign n2592 = Pinreg_43_ & n505;
  assign n2593 = Pdata_41_ & ~n505;
  assign Pdata_new_9_ = n2592 | n2593;
  assign n2595 = Pinreg_51_ & n505;
  assign n2596 = Pdata_40_ & ~n505;
  assign Pdata_new_8_ = n2595 | n2596;
  assign n2598 = Pdata_in_1_ & n505;
  assign n2599 = Pdata_39_ & ~n505;
  assign Pdata_new_7_ = n2598 | n2599;
  assign n2601 = Pinreg_1_ & n505;
  assign n2602 = Pdata_38_ & ~n505;
  assign Pdata_new_6_ = n2601 | n2602;
  assign n2604 = Pinreg_9_ & n505;
  assign n2605 = Pdata_37_ & ~n505;
  assign Pdata_new_5_ = n2604 | n2605;
  assign n2607 = Pinreg_17_ & n505;
  assign n2608 = Pdata_36_ & ~n505;
  assign Pdata_new_4_ = n2607 | n2608;
  assign n2610 = Pinreg_25_ & n505;
  assign n2611 = Pdata_35_ & ~n505;
  assign Pdata_new_3_ = n2610 | n2611;
  assign n2613 = Pinreg_33_ & n505;
  assign n2614 = Pdata_34_ & ~n505;
  assign Pdata_new_2_ = n2613 | n2614;
  assign n2616 = Pinreg_41_ & n505;
  assign n2617 = Pdata_33_ & ~n505;
  assign Pdata_new_1_ = n2616 | n2617;
  assign n2619 = Pinreg_49_ & n505;
  assign n2620 = Pdata_32_ & ~n505;
  assign Pdata_new_0_ = n2619 | n2620;
  assign n2622 = ~Pcount_3_ & ~n504;
  assign n2623 = ~Preset_0_ & ~n2622;
  assign Pcount_new_3_ = ~n505 & n2623;
  assign n2625 = ~Pcount_2_ & ~n503;
  assign n2626 = ~Preset_0_ & ~n2625;
  assign Pcount_new_2_ = ~n504 & n2626;
  assign n2628 = Pload_key_0_ & n505;
  assign n2629 = ~Preset_0_ & ~n2628;
  assign n2630 = ~Pcount_1_ & ~Pcount_0_;
  assign n2631 = n2629 & ~n2630;
  assign Pcount_new_1_ = ~n503 & n2631;
  assign Pcount_new_0_ = ~Pcount_0_ & n2629;
  assign n2634 = Pencrypt_mode_0_ & Pencrypt_0_;
  assign n2635 = ~Pencrypt_mode_0_ & ~Pencrypt_0_;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = n505 & n2636;
  assign n2638 = n2629 & n2637;
  assign n2639 = PD_27_ & n2638;
  assign n2640 = n2629 & ~n2637;
  assign n2641 = ~Pencrypt_mode_0_ & n2640;
  assign n2642 = ~Pcount_3_ & ~Pcount_0_;
  assign n2643 = Pcount_2_ & Pcount_1_;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = ~Pcount_2_ & ~Pcount_1_;
  assign n2646 = n2642 & ~n2645;
  assign n2647 = ~n2644 & ~n2646;
  assign n2648 = n2641 & ~n2647;
  assign n2649 = PD_25_ & n2648;
  assign n2650 = ~n2639 & ~n2649;
  assign n2651 = Pencrypt_mode_0_ & n2640;
  assign n2652 = ~n2647 & n2651;
  assign n2653 = PD_1_ & n2652;
  assign n2654 = ~Preset_0_ & n2628;
  assign n2655 = ~Pencrypt_0_ & n2654;
  assign n2656 = Pdata_in_3_ & n2655;
  assign n2657 = Pencrypt_0_ & n2654;
  assign n2658 = Pinreg_54_ & n2657;
  assign n2659 = ~n2656 & ~n2658;
  assign n2660 = ~n2653 & n2659;
  assign n2661 = n2647 & n2651;
  assign n2662 = PD_0_ & n2661;
  assign n2663 = n2641 & n2647;
  assign n2664 = PD_26_ & n2663;
  assign n2665 = ~n2662 & ~n2664;
  assign n2666 = n2660 & n2665;
  assign PD_new_27_ = ~n2650 | ~n2666;
  assign n2668 = PD_24_ & n2648;
  assign n2669 = PD_27_ & n2661;
  assign n2670 = ~n2668 & ~n2669;
  assign n2671 = PD_25_ & n2663;
  assign n2672 = n2670 & ~n2671;
  assign n2673 = PD_26_ & n2638;
  assign n2674 = Pinreg_3_ & n2655;
  assign n2675 = Pdata_in_3_ & n2657;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2673 & n2676;
  assign n2678 = PD_0_ & n2652;
  assign n2679 = n2677 & ~n2678;
  assign PD_new_26_ = ~n2672 | ~n2679;
  assign n2681 = PD_25_ & n2638;
  assign n2682 = PD_27_ & n2652;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = PD_24_ & n2663;
  assign n2685 = Pinreg_11_ & n2655;
  assign n2686 = Pinreg_3_ & n2657;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = ~n2684 & n2687;
  assign n2689 = PD_26_ & n2661;
  assign n2690 = PD_23_ & n2648;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2688 & n2691;
  assign PD_new_25_ = ~n2683 | ~n2692;
  assign n2694 = PD_26_ & n2652;
  assign n2695 = PD_22_ & n2648;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = PD_23_ & n2663;
  assign n2698 = n2696 & ~n2697;
  assign n2699 = Pinreg_19_ & n2655;
  assign n2700 = Pinreg_11_ & n2657;
  assign n2701 = PD_24_ & n2638;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = ~n2699 & n2702;
  assign n2704 = PD_25_ & n2661;
  assign n2705 = n2703 & ~n2704;
  assign PD_new_24_ = ~n2698 | ~n2705;
  assign n2707 = PD_22_ & n2663;
  assign n2708 = PD_24_ & n2661;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = PD_21_ & n2648;
  assign n2711 = n2709 & ~n2710;
  assign n2712 = Pdata_in_4_ & n2655;
  assign n2713 = Pinreg_19_ & n2657;
  assign n2714 = PD_23_ & n2638;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = ~n2712 & n2715;
  assign n2717 = PD_25_ & n2652;
  assign n2718 = n2716 & ~n2717;
  assign PD_new_23_ = ~n2711 | ~n2718;
  assign n2720 = PD_20_ & n2648;
  assign n2721 = PD_24_ & n2652;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = PD_23_ & n2661;
  assign n2724 = n2722 & ~n2723;
  assign n2725 = Pinreg_4_ & n2655;
  assign n2726 = Pdata_in_4_ & n2657;
  assign n2727 = PD_22_ & n2638;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = ~n2725 & n2728;
  assign n2730 = PD_21_ & n2663;
  assign n2731 = n2729 & ~n2730;
  assign PD_new_22_ = ~n2724 | ~n2731;
  assign n2733 = PD_22_ & n2661;
  assign n2734 = PD_20_ & n2663;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = PD_23_ & n2652;
  assign n2737 = n2735 & ~n2736;
  assign n2738 = Pinreg_4_ & n2657;
  assign n2739 = Pinreg_12_ & n2655;
  assign n2740 = PD_21_ & n2638;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = ~n2738 & n2741;
  assign n2743 = PD_19_ & n2648;
  assign n2744 = n2742 & ~n2743;
  assign PD_new_21_ = ~n2737 | ~n2744;
  assign n2746 = PD_18_ & n2648;
  assign n2747 = PD_21_ & n2661;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = PD_22_ & n2652;
  assign n2750 = n2748 & ~n2749;
  assign n2751 = Pinreg_12_ & n2657;
  assign n2752 = PD_20_ & n2638;
  assign n2753 = Pinreg_20_ & n2655;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~n2751 & n2754;
  assign n2756 = PD_19_ & n2663;
  assign n2757 = n2755 & ~n2756;
  assign PD_new_20_ = ~n2750 | ~n2757;
  assign n2759 = PD_17_ & n2648;
  assign n2760 = PD_21_ & n2652;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = PD_20_ & n2661;
  assign n2763 = n2761 & ~n2762;
  assign n2764 = Pinreg_28_ & n2655;
  assign n2765 = PD_19_ & n2638;
  assign n2766 = Pinreg_20_ & n2657;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = ~n2764 & n2767;
  assign n2769 = PD_18_ & n2663;
  assign n2770 = n2768 & ~n2769;
  assign PD_new_19_ = ~n2763 | ~n2770;
  assign n2772 = PD_19_ & n2661;
  assign n2773 = PD_20_ & n2652;
  assign n2774 = Pinreg_36_ & n2655;
  assign n2775 = PD_18_ & n2638;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = ~n2773 & n2776;
  assign n2778 = ~n2772 & n2777;
  assign n2779 = Pinreg_28_ & n2657;
  assign n2780 = PD_17_ & n2663;
  assign n2781 = PD_16_ & n2648;
  assign n2782 = ~n2780 & ~n2781;
  assign n2783 = ~n2779 & n2782;
  assign PD_new_18_ = ~n2778 | ~n2783;
  assign n2785 = Pinreg_44_ & n2655;
  assign n2786 = PD_15_ & n2648;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = PD_18_ & n2661;
  assign n2789 = Pinreg_36_ & n2657;
  assign n2790 = PD_17_ & n2638;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = ~n2788 & n2791;
  assign n2793 = PD_16_ & n2663;
  assign n2794 = PD_19_ & n2652;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = n2792 & n2795;
  assign PD_new_17_ = ~n2787 | ~n2796;
  assign n2798 = PD_15_ & n2663;
  assign n2799 = PD_18_ & n2652;
  assign n2800 = Pinreg_52_ & n2655;
  assign n2801 = Pinreg_44_ & n2657;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = ~n2799 & n2802;
  assign n2804 = ~n2798 & n2803;
  assign n2805 = PD_16_ & n2638;
  assign n2806 = PD_14_ & n2648;
  assign n2807 = PD_17_ & n2661;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = ~n2805 & n2808;
  assign PD_new_16_ = ~n2804 | ~n2809;
  assign n2811 = PD_13_ & n2648;
  assign n2812 = PD_17_ & n2652;
  assign n2813 = ~n2811 & ~n2812;
  assign n2814 = PD_14_ & n2663;
  assign n2815 = n2813 & ~n2814;
  assign n2816 = Pinreg_52_ & n2657;
  assign n2817 = Pdata_in_5_ & n2655;
  assign n2818 = PD_15_ & n2638;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = ~n2816 & n2819;
  assign n2821 = PD_16_ & n2661;
  assign n2822 = n2820 & ~n2821;
  assign PD_new_15_ = ~n2815 | ~n2822;
  assign n2824 = PD_13_ & n2663;
  assign n2825 = PD_15_ & n2661;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = PD_12_ & n2648;
  assign n2828 = n2826 & ~n2827;
  assign n2829 = Pdata_in_5_ & n2657;
  assign n2830 = PD_14_ & n2638;
  assign n2831 = Pinreg_5_ & n2655;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n2829 & n2832;
  assign n2834 = PD_16_ & n2652;
  assign n2835 = n2833 & ~n2834;
  assign PD_new_14_ = ~n2828 | ~n2835;
  assign n2837 = PD_15_ & n2652;
  assign n2838 = PD_11_ & n2648;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = PD_12_ & n2663;
  assign n2841 = n2839 & ~n2840;
  assign n2842 = Pinreg_13_ & n2655;
  assign n2843 = PD_13_ & n2638;
  assign n2844 = Pinreg_5_ & n2657;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = ~n2842 & n2845;
  assign n2847 = PD_14_ & n2661;
  assign n2848 = n2846 & ~n2847;
  assign PD_new_13_ = ~n2841 | ~n2848;
  assign n2850 = PD_11_ & n2663;
  assign n2851 = PD_10_ & n2648;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = PD_14_ & n2652;
  assign n2854 = n2852 & ~n2853;
  assign n2855 = Pinreg_13_ & n2657;
  assign n2856 = Pinreg_21_ & n2655;
  assign n2857 = PD_12_ & n2638;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = ~n2855 & n2858;
  assign n2860 = PD_13_ & n2661;
  assign n2861 = n2859 & ~n2860;
  assign PD_new_12_ = ~n2854 | ~n2861;
  assign n2863 = PD_9_ & n2648;
  assign n2864 = PD_13_ & n2652;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = PD_12_ & n2661;
  assign n2867 = n2865 & ~n2866;
  assign n2868 = Pinreg_21_ & n2657;
  assign n2869 = Pinreg_29_ & n2655;
  assign n2870 = PD_11_ & n2638;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = ~n2868 & n2871;
  assign n2873 = PD_10_ & n2663;
  assign n2874 = n2872 & ~n2873;
  assign PD_new_11_ = ~n2867 | ~n2874;
  assign n2876 = PD_8_ & n2648;
  assign n2877 = PD_11_ & n2661;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = PD_12_ & n2652;
  assign n2880 = n2878 & ~n2879;
  assign n2881 = PD_10_ & n2638;
  assign n2882 = Pinreg_37_ & n2655;
  assign n2883 = Pinreg_29_ & n2657;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~n2881 & n2884;
  assign n2886 = PD_9_ & n2663;
  assign n2887 = n2885 & ~n2886;
  assign PD_new_10_ = ~n2880 | ~n2887;
  assign n2889 = PD_10_ & n2661;
  assign n2890 = PD_11_ & n2652;
  assign n2891 = Pinreg_45_ & n2655;
  assign n2892 = Pinreg_37_ & n2657;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = ~n2890 & n2893;
  assign n2895 = ~n2889 & n2894;
  assign n2896 = PD_9_ & n2638;
  assign n2897 = PD_7_ & n2648;
  assign n2898 = PD_8_ & n2663;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & n2899;
  assign PD_new_9_ = ~n2895 | ~n2900;
  assign n2902 = Pinreg_45_ & n2657;
  assign n2903 = PD_6_ & n2648;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = PD_10_ & n2652;
  assign n2906 = PD_8_ & n2638;
  assign n2907 = Pinreg_53_ & n2655;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = ~n2905 & n2908;
  assign n2910 = PD_7_ & n2663;
  assign n2911 = PD_9_ & n2661;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = n2909 & n2912;
  assign PD_new_8_ = ~n2904 | ~n2913;
  assign n2915 = PD_5_ & n2648;
  assign n2916 = PD_6_ & n2663;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = PD_9_ & n2652;
  assign n2919 = n2917 & ~n2918;
  assign n2920 = PD_7_ & n2638;
  assign n2921 = Pdata_in_6_ & n2655;
  assign n2922 = Pinreg_53_ & n2657;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2920 & n2923;
  assign n2925 = PD_8_ & n2661;
  assign n2926 = n2924 & ~n2925;
  assign PD_new_7_ = ~n2919 | ~n2926;
  assign n2928 = PD_4_ & n2648;
  assign n2929 = PD_7_ & n2661;
  assign n2930 = ~n2928 & ~n2929;
  assign n2931 = PD_5_ & n2663;
  assign n2932 = n2930 & ~n2931;
  assign n2933 = Pinreg_6_ & n2655;
  assign n2934 = Pdata_in_6_ & n2657;
  assign n2935 = PD_6_ & n2638;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = ~n2933 & n2936;
  assign n2938 = PD_8_ & n2652;
  assign n2939 = n2937 & ~n2938;
  assign PD_new_6_ = ~n2932 | ~n2939;
  assign n2941 = PD_6_ & n2661;
  assign n2942 = PD_4_ & n2663;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = PD_7_ & n2652;
  assign n2945 = n2943 & ~n2944;
  assign n2946 = Pinreg_6_ & n2657;
  assign n2947 = Pinreg_14_ & n2655;
  assign n2948 = PD_5_ & n2638;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = ~n2946 & n2949;
  assign n2951 = PD_3_ & n2648;
  assign n2952 = n2950 & ~n2951;
  assign PD_new_5_ = ~n2945 | ~n2952;
  assign n2954 = PD_5_ & n2661;
  assign n2955 = PD_2_ & n2648;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = PD_3_ & n2663;
  assign n2958 = n2956 & ~n2957;
  assign n2959 = Pinreg_14_ & n2657;
  assign n2960 = PD_4_ & n2638;
  assign n2961 = Pinreg_22_ & n2655;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2959 & n2962;
  assign n2964 = PD_6_ & n2652;
  assign n2965 = n2963 & ~n2964;
  assign PD_new_4_ = ~n2958 | ~n2965;
  assign n2967 = PD_4_ & n2661;
  assign n2968 = PD_5_ & n2652;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970 = PD_1_ & n2648;
  assign n2971 = n2969 & ~n2970;
  assign n2972 = Pinreg_22_ & n2657;
  assign n2973 = PD_3_ & n2638;
  assign n2974 = Pinreg_30_ & n2655;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = ~n2972 & n2975;
  assign n2977 = PD_2_ & n2663;
  assign n2978 = n2976 & ~n2977;
  assign PD_new_3_ = ~n2971 | ~n2978;
  assign n2980 = PD_1_ & n2663;
  assign n2981 = PD_0_ & n2648;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = PD_3_ & n2661;
  assign n2984 = n2982 & ~n2983;
  assign n2985 = Pinreg_30_ & n2657;
  assign n2986 = PD_2_ & n2638;
  assign n2987 = Pinreg_38_ & n2655;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = ~n2985 & n2988;
  assign n2990 = PD_4_ & n2652;
  assign n2991 = n2989 & ~n2990;
  assign PD_new_2_ = ~n2984 | ~n2991;
  assign n2993 = PD_2_ & n2661;
  assign n2994 = PD_27_ & n2648;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = PD_3_ & n2652;
  assign n2997 = n2995 & ~n2996;
  assign n2998 = Pinreg_38_ & n2657;
  assign n2999 = PD_1_ & n2638;
  assign n3000 = Pinreg_46_ & n2655;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = ~n2998 & n3001;
  assign n3003 = PD_0_ & n2663;
  assign n3004 = n3002 & ~n3003;
  assign PD_new_1_ = ~n2997 | ~n3004;
  assign n3006 = PD_26_ & n2648;
  assign n3007 = PD_2_ & n2652;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = PD_27_ & n2663;
  assign n3010 = n3008 & ~n3009;
  assign n3011 = Pinreg_54_ & n2655;
  assign n3012 = Pinreg_46_ & n2657;
  assign n3013 = PD_0_ & n2638;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = ~n3011 & n3014;
  assign n3016 = PD_1_ & n2661;
  assign n3017 = n3015 & ~n3016;
  assign PD_new_0_ = ~n3010 | ~n3017;
  assign n3019 = PC_1_ & n2652;
  assign n3020 = PC_25_ & n2648;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = PC_0_ & n2661;
  assign n3023 = n3021 & ~n3022;
  assign n3024 = Pinreg_27_ & n2655;
  assign n3025 = Pinreg_48_ & n2657;
  assign n3026 = PC_27_ & n2638;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = ~n3024 & n3027;
  assign n3029 = PC_26_ & n2663;
  assign n3030 = n3028 & ~n3029;
  assign PC_new_27_ = ~n3023 | ~n3030;
  assign n3032 = PC_26_ & n2638;
  assign n3033 = PC_0_ & n2652;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = PC_27_ & n2661;
  assign n3036 = Pinreg_35_ & n2655;
  assign n3037 = Pinreg_27_ & n2657;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = ~n3035 & n3038;
  assign n3040 = PC_24_ & n2648;
  assign n3041 = PC_25_ & n2663;
  assign n3042 = ~n3040 & ~n3041;
  assign n3043 = n3039 & n3042;
  assign PC_new_26_ = ~n3034 | ~n3043;
  assign n3045 = Pinreg_43_ & n2655;
  assign n3046 = PC_23_ & n2648;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = PC_27_ & n2652;
  assign n3049 = Pinreg_35_ & n2657;
  assign n3050 = PC_25_ & n2638;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = ~n3048 & n3051;
  assign n3053 = PC_26_ & n2661;
  assign n3054 = PC_24_ & n2663;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = n3052 & n3055;
  assign PC_new_25_ = ~n3047 | ~n3056;
  assign n3058 = PC_23_ & n2663;
  assign n3059 = PC_25_ & n2661;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = PC_26_ & n2652;
  assign n3062 = n3060 & ~n3061;
  assign n3063 = Pinreg_51_ & n2655;
  assign n3064 = PC_24_ & n2638;
  assign n3065 = Pinreg_43_ & n2657;
  assign n3066 = ~n3064 & ~n3065;
  assign n3067 = ~n3063 & n3066;
  assign n3068 = PC_22_ & n2648;
  assign n3069 = n3067 & ~n3068;
  assign PC_new_24_ = ~n3062 | ~n3069;
  assign n3071 = PC_22_ & n2663;
  assign n3072 = PC_24_ & n2661;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = PC_25_ & n2652;
  assign n3075 = n3073 & ~n3074;
  assign n3076 = PC_23_ & n2638;
  assign n3077 = Pdata_in_2_ & n2655;
  assign n3078 = Pinreg_51_ & n2657;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = ~n3076 & n3079;
  assign n3081 = PC_21_ & n2648;
  assign n3082 = n3080 & ~n3081;
  assign PC_new_23_ = ~n3075 | ~n3082;
  assign n3084 = PC_24_ & n2652;
  assign n3085 = PC_21_ & n2663;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = PC_23_ & n2661;
  assign n3088 = n3086 & ~n3087;
  assign n3089 = Pinreg_2_ & n2655;
  assign n3090 = PC_22_ & n2638;
  assign n3091 = Pdata_in_2_ & n2657;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = ~n3089 & n3092;
  assign n3094 = PC_20_ & n2648;
  assign n3095 = n3093 & ~n3094;
  assign PC_new_22_ = ~n3088 | ~n3095;
  assign n3097 = PC_23_ & n2652;
  assign n3098 = PC_19_ & n2648;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = PC_20_ & n2663;
  assign n3101 = n3099 & ~n3100;
  assign n3102 = Pinreg_2_ & n2657;
  assign n3103 = PC_21_ & n2638;
  assign n3104 = Pinreg_10_ & n2655;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = ~n3102 & n3105;
  assign n3107 = PC_22_ & n2661;
  assign n3108 = n3106 & ~n3107;
  assign PC_new_21_ = ~n3101 | ~n3108;
  assign n3110 = PC_18_ & n2648;
  assign n3111 = PC_22_ & n2652;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = PC_21_ & n2661;
  assign n3114 = n3112 & ~n3113;
  assign n3115 = Pinreg_18_ & n2655;
  assign n3116 = Pinreg_10_ & n2657;
  assign n3117 = PC_20_ & n2638;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = ~n3115 & n3118;
  assign n3120 = PC_19_ & n2663;
  assign n3121 = n3119 & ~n3120;
  assign PC_new_20_ = ~n3114 | ~n3121;
  assign n3123 = Pinreg_26_ & n2655;
  assign n3124 = PC_18_ & n2663;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = PC_17_ & n2648;
  assign n3127 = PC_19_ & n2638;
  assign n3128 = Pinreg_18_ & n2657;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = ~n3126 & n3129;
  assign n3131 = PC_20_ & n2661;
  assign n3132 = PC_21_ & n2652;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n3130 & n3133;
  assign PC_new_19_ = ~n3125 | ~n3134;
  assign n3136 = PC_17_ & n2663;
  assign n3137 = PC_16_ & n2648;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = PC_19_ & n2661;
  assign n3140 = n3138 & ~n3139;
  assign n3141 = PC_18_ & n2638;
  assign n3142 = Pinreg_34_ & n2655;
  assign n3143 = Pinreg_26_ & n2657;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3141 & n3144;
  assign n3146 = PC_20_ & n2652;
  assign n3147 = n3145 & ~n3146;
  assign PC_new_18_ = ~n3140 | ~n3147;
  assign n3149 = PC_18_ & n2661;
  assign n3150 = PC_16_ & n2663;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = PC_19_ & n2652;
  assign n3153 = n3151 & ~n3152;
  assign n3154 = Pinreg_34_ & n2657;
  assign n3155 = PC_17_ & n2638;
  assign n3156 = Pinreg_42_ & n2655;
  assign n3157 = ~n3155 & ~n3156;
  assign n3158 = ~n3154 & n3157;
  assign n3159 = PC_15_ & n2648;
  assign n3160 = n3158 & ~n3159;
  assign PC_new_17_ = ~n3153 | ~n3160;
  assign n3162 = PC_16_ & n2638;
  assign n3163 = PC_18_ & n2652;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = PC_14_ & n2648;
  assign n3166 = Pinreg_42_ & n2657;
  assign n3167 = Pinreg_50_ & n2655;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = ~n3165 & n3168;
  assign n3170 = PC_15_ & n2663;
  assign n3171 = PC_17_ & n2661;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = n3169 & n3172;
  assign PC_new_16_ = ~n3164 | ~n3173;
  assign n3175 = PC_16_ & n2661;
  assign n3176 = PC_14_ & n2663;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = PC_17_ & n2652;
  assign n3179 = n3177 & ~n3178;
  assign n3180 = PC_15_ & n2638;
  assign n3181 = Pdata_in_1_ & n2655;
  assign n3182 = Pinreg_50_ & n2657;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = ~n3180 & n3183;
  assign n3185 = PC_13_ & n2648;
  assign n3186 = n3184 & ~n3185;
  assign PC_new_15_ = ~n3179 | ~n3186;
  assign n3188 = PC_16_ & n2652;
  assign n3189 = PC_12_ & n2648;
  assign n3190 = ~n3188 & ~n3189;
  assign n3191 = PC_13_ & n2663;
  assign n3192 = n3190 & ~n3191;
  assign n3193 = Pinreg_1_ & n2655;
  assign n3194 = Pdata_in_1_ & n2657;
  assign n3195 = PC_14_ & n2638;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = ~n3193 & n3196;
  assign n3198 = PC_15_ & n2661;
  assign n3199 = n3197 & ~n3198;
  assign PC_new_14_ = ~n3192 | ~n3199;
  assign n3201 = PC_12_ & n2663;
  assign n3202 = PC_11_ & n2648;
  assign n3203 = ~n3201 & ~n3202;
  assign n3204 = PC_14_ & n2661;
  assign n3205 = n3203 & ~n3204;
  assign n3206 = Pinreg_9_ & n2655;
  assign n3207 = Pinreg_1_ & n2657;
  assign n3208 = PC_13_ & n2638;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~n3206 & n3209;
  assign n3211 = PC_15_ & n2652;
  assign n3212 = n3210 & ~n3211;
  assign PC_new_13_ = ~n3205 | ~n3212;
  assign n3214 = PC_10_ & n2648;
  assign n3215 = PC_13_ & n2661;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = PC_14_ & n2652;
  assign n3218 = n3216 & ~n3217;
  assign n3219 = Pinreg_17_ & n2655;
  assign n3220 = PC_12_ & n2638;
  assign n3221 = Pinreg_9_ & n2657;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~n3219 & n3222;
  assign n3224 = PC_11_ & n2663;
  assign n3225 = n3223 & ~n3224;
  assign PC_new_12_ = ~n3218 | ~n3225;
  assign n3227 = Pinreg_25_ & n2655;
  assign n3228 = PC_9_ & n2648;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = PC_12_ & n2661;
  assign n3231 = Pinreg_17_ & n2657;
  assign n3232 = PC_11_ & n2638;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = ~n3230 & n3233;
  assign n3235 = PC_10_ & n2663;
  assign n3236 = PC_13_ & n2652;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = n3234 & n3237;
  assign PC_new_11_ = ~n3229 | ~n3238;
  assign n3240 = PC_8_ & n2648;
  assign n3241 = PC_9_ & n2663;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = PC_12_ & n2652;
  assign n3244 = n3242 & ~n3243;
  assign n3245 = Pinreg_25_ & n2657;
  assign n3246 = PC_10_ & n2638;
  assign n3247 = Pinreg_33_ & n2655;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = ~n3245 & n3248;
  assign n3250 = PC_11_ & n2661;
  assign n3251 = n3249 & ~n3250;
  assign PC_new_10_ = ~n3244 | ~n3251;
  assign n3253 = PC_11_ & n2652;
  assign n3254 = PC_8_ & n2663;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = PC_7_ & n2648;
  assign n3257 = n3255 & ~n3256;
  assign n3258 = PC_9_ & n2638;
  assign n3259 = Pinreg_41_ & n2655;
  assign n3260 = Pinreg_33_ & n2657;
  assign n3261 = ~n3259 & ~n3260;
  assign n3262 = ~n3258 & n3261;
  assign n3263 = PC_10_ & n2661;
  assign n3264 = n3262 & ~n3263;
  assign PC_new_9_ = ~n3257 | ~n3264;
  assign n3266 = PC_7_ & n2663;
  assign n3267 = PC_8_ & n2638;
  assign n3268 = PC_6_ & n2648;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = ~n3266 & n3269;
  assign n3271 = Pinreg_49_ & n2655;
  assign n3272 = Pinreg_41_ & n2657;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = PC_10_ & n2652;
  assign n3275 = PC_9_ & n2661;
  assign n3276 = ~n3274 & ~n3275;
  assign n3277 = n3273 & n3276;
  assign PC_new_8_ = ~n3270 | ~n3277;
  assign n3279 = PC_6_ & n2663;
  assign n3280 = PC_9_ & n2652;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = PC_8_ & n2661;
  assign n3283 = n3281 & ~n3282;
  assign n3284 = PC_7_ & n2638;
  assign n3285 = Pinreg_49_ & n2657;
  assign n3286 = Pdata_in_0_ & n2655;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n3284 & n3287;
  assign n3289 = PC_5_ & n2648;
  assign n3290 = n3288 & ~n3289;
  assign PC_new_7_ = ~n3283 | ~n3290;
  assign n3292 = PC_7_ & n2661;
  assign n3293 = PC_8_ & n2652;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = PC_4_ & n2648;
  assign n3296 = n3294 & ~n3295;
  assign n3297 = PC_6_ & n2638;
  assign n3298 = Pdata_in_0_ & n2657;
  assign n3299 = Pinreg_0_ & n2655;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = ~n3297 & n3300;
  assign n3302 = PC_5_ & n2663;
  assign n3303 = n3301 & ~n3302;
  assign PC_new_6_ = ~n3296 | ~n3303;
  assign n3305 = Pinreg_8_ & n2655;
  assign n3306 = PC_4_ & n2663;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = PC_7_ & n2652;
  assign n3309 = PC_5_ & n2638;
  assign n3310 = Pinreg_0_ & n2657;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = ~n3308 & n3311;
  assign n3313 = PC_6_ & n2661;
  assign n3314 = PC_3_ & n2648;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = n3312 & n3315;
  assign PC_new_5_ = ~n3307 | ~n3316;
  assign n3318 = PC_5_ & n2661;
  assign n3319 = PC_6_ & n2652;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = PC_2_ & n2648;
  assign n3322 = n3320 & ~n3321;
  assign n3323 = Pinreg_8_ & n2657;
  assign n3324 = PC_4_ & n2638;
  assign n3325 = Pinreg_16_ & n2655;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = ~n3323 & n3326;
  assign n3328 = PC_3_ & n2663;
  assign n3329 = n3327 & ~n3328;
  assign PC_new_4_ = ~n3322 | ~n3329;
  assign n3331 = PC_1_ & n2648;
  assign n3332 = PC_5_ & n2652;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = PC_4_ & n2661;
  assign n3335 = n3333 & ~n3334;
  assign n3336 = Pinreg_16_ & n2657;
  assign n3337 = PC_3_ & n2638;
  assign n3338 = Pinreg_24_ & n2655;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = ~n3336 & n3339;
  assign n3341 = PC_2_ & n2663;
  assign n3342 = n3340 & ~n3341;
  assign PC_new_3_ = ~n3335 | ~n3342;
  assign n3344 = Pinreg_32_ & n2655;
  assign n3345 = PC_3_ & n2661;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = PC_0_ & n2648;
  assign n3348 = PC_2_ & n2638;
  assign n3349 = Pinreg_24_ & n2657;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = ~n3347 & n3350;
  assign n3352 = PC_4_ & n2652;
  assign n3353 = PC_1_ & n2663;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = n3351 & n3354;
  assign PC_new_2_ = ~n3346 | ~n3355;
  assign n3357 = PC_2_ & n2661;
  assign n3358 = PC_0_ & n2663;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = PC_3_ & n2652;
  assign n3361 = n3359 & ~n3360;
  assign n3362 = PC_1_ & n2638;
  assign n3363 = Pinreg_40_ & n2655;
  assign n3364 = Pinreg_32_ & n2657;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = ~n3362 & n3365;
  assign n3367 = PC_27_ & n2648;
  assign n3368 = n3366 & ~n3367;
  assign PC_new_1_ = ~n3361 | ~n3368;
  assign n3370 = PC_1_ & n2661;
  assign n3371 = PC_26_ & n2648;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = PC_27_ & n2663;
  assign n3374 = n3372 & ~n3373;
  assign n3375 = PC_0_ & n2638;
  assign n3376 = Pinreg_40_ & n2657;
  assign n3377 = Pinreg_48_ & n2655;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3375 & n3378;
  assign n3380 = PC_2_ & n2652;
  assign n3381 = n3379 & ~n3380;
  assign PC_new_0_ = ~n3374 | ~n3381;
endmodule


