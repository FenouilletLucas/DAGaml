// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:37 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_;
  wire n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n996, n997,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1919, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2432, n2433, n2434, n2436, n2437, n2439, n2440, n2441, n2442,
    n2444, n2445, n2446, n2447, n2448, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2463, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2495, n2496, n2498, n2499, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2580, n2581, n2582,
    n2584, n2585, n2586, n2587, n2588, n2590, n2591, n2592, n2593, n2594,
    n2595, n2597, n2598, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3257, n3258, n3260, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3328;
  assign n63 = i_0_ & ~i_1_;
  assign n64 = ~i_3_ & ~i_4_;
  assign n65 = i_5_ & n64;
  assign n66 = ~i_10_ & ~i_11_;
  assign n67 = ~i_9_ & n66;
  assign n68 = ~i_15_ & n67;
  assign n69 = ~i_12_ & ~i_13_;
  assign n70 = ~i_14_ & n69;
  assign n71 = n68 & n70;
  assign n72 = i_1_ & ~i_2_;
  assign n73 = i_0_ & n72;
  assign n74 = n71 & n73;
  assign n75 = n65 & n74;
  assign n76 = ~i_6_ & ~i_8_;
  assign n77 = ~i_7_ & n76;
  assign n78 = n75 & n77;
  assign o_0_ = n63 | n78;
  assign o_2_ = n75 & n76;
  assign n81 = i_7_ & o_2_;
  assign n82 = i_0_ & i_2_;
  assign n83 = ~i_2_ & ~n63;
  assign n84 = ~n82 & ~n83;
  assign o_1_ = n81 | n84;
  assign n86 = ~i_5_ & n64;
  assign n87 = ~i_0_ & n72;
  assign n88 = n86 & n87;
  assign n89 = ~i_7_ & ~i_8_;
  assign n90 = n88 & n89;
  assign n91 = ~i_12_ & i_13_;
  assign n92 = i_9_ & n66;
  assign n93 = ~i_15_ & n92;
  assign n94 = ~i_14_ & n93;
  assign n95 = n91 & n94;
  assign n96 = n90 & n95;
  assign n97 = i_14_ & n69;
  assign n98 = i_10_ & ~i_11_;
  assign n99 = i_9_ & n98;
  assign n100 = ~i_15_ & n99;
  assign n101 = n97 & n100;
  assign n102 = i_15_ & n99;
  assign n103 = n70 & n102;
  assign n104 = i_13_ & ~i_14_;
  assign n105 = ~i_12_ & n104;
  assign n106 = n100 & n105;
  assign n107 = ~n103 & ~n106;
  assign n108 = ~n101 & n107;
  assign n109 = n90 & ~n108;
  assign n110 = ~n96 & ~n109;
  assign n111 = ~i_6_ & ~n110;
  assign n112 = ~i_6_ & i_7_;
  assign n113 = i_14_ & n93;
  assign n114 = n69 & n113;
  assign n115 = ~i_9_ & n98;
  assign n116 = i_15_ & n115;
  assign n117 = n70 & n116;
  assign n118 = ~i_15_ & n115;
  assign n119 = n97 & n118;
  assign n120 = ~n117 & ~n119;
  assign n121 = i_15_ & n92;
  assign n122 = n70 & n121;
  assign n123 = n105 & n118;
  assign n124 = ~n122 & ~n123;
  assign n125 = n120 & n124;
  assign n126 = ~n114 & n125;
  assign n127 = n76 & ~n126;
  assign n128 = ~n112 & ~n127;
  assign n129 = n88 & ~n128;
  assign n130 = n70 & n118;
  assign n131 = n69 & n94;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~n71 & n132;
  assign n134 = ~i_6_ & ~i_7_;
  assign n135 = i_8_ & n134;
  assign n136 = n88 & n135;
  assign n137 = ~n133 & n136;
  assign n138 = ~n129 & ~n137;
  assign n139 = ~n111 & n138;
  assign n140 = i_6_ & ~n110;
  assign n141 = i_6_ & ~i_7_;
  assign n142 = i_8_ & n141;
  assign n143 = n88 & n142;
  assign n144 = ~n133 & n143;
  assign n145 = i_6_ & n114;
  assign n146 = n90 & n145;
  assign n147 = ~n144 & ~n146;
  assign n148 = ~n140 & n147;
  assign n149 = i_6_ & i_7_;
  assign n150 = ~i_8_ & n141;
  assign n151 = ~n125 & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = n88 & ~n152;
  assign n154 = ~i_3_ & n63;
  assign n155 = ~i_4_ & n154;
  assign n156 = ~n153 & ~n155;
  assign n157 = n148 & n156;
  assign o_3_ = ~n139 | ~n157;
  assign n159 = ~i_3_ & i_4_;
  assign n160 = ~i_5_ & n159;
  assign n161 = n87 & n160;
  assign n162 = n89 & ~n108;
  assign n163 = n161 & n162;
  assign n164 = i_6_ & n163;
  assign n165 = i_5_ & n159;
  assign n166 = n63 & n165;
  assign n167 = ~n95 & n126;
  assign n168 = n150 & ~n167;
  assign n169 = ~n149 & ~n168;
  assign n170 = n161 & ~n169;
  assign n171 = ~n166 & ~n170;
  assign n172 = n142 & n161;
  assign n173 = ~n132 & n172;
  assign n174 = n171 & ~n173;
  assign n175 = ~n164 & n174;
  assign n176 = n135 & n161;
  assign n177 = ~n132 & n176;
  assign n178 = n77 & n161;
  assign n179 = ~n167 & n178;
  assign n180 = n87 & n112;
  assign n181 = ~n63 & ~n180;
  assign n182 = n160 & ~n181;
  assign n183 = ~n179 & ~n182;
  assign n184 = ~n108 & n178;
  assign n185 = n183 & ~n184;
  assign n186 = ~n177 & n185;
  assign o_4_ = ~n175 | ~n186;
  assign n188 = i_10_ & i_11_;
  assign n189 = i_9_ & n188;
  assign n190 = ~i_15_ & n189;
  assign n191 = i_12_ & ~i_13_;
  assign n192 = ~i_14_ & n191;
  assign n193 = n190 & n192;
  assign n194 = ~i_0_ & ~i_1_;
  assign n195 = ~i_2_ & n194;
  assign n196 = n160 & n195;
  assign n197 = n141 & n196;
  assign n198 = i_8_ & n197;
  assign n199 = n65 & n195;
  assign n200 = n141 & n199;
  assign n201 = i_8_ & n200;
  assign n202 = n165 & n195;
  assign n203 = i_7_ & n202;
  assign n204 = ~i_6_ & i_8_;
  assign n205 = n203 & n204;
  assign n206 = ~n201 & ~n205;
  assign n207 = ~n198 & n206;
  assign n208 = n193 & ~n207;
  assign n209 = i_8_ & n203;
  assign n210 = ~i_10_ & i_11_;
  assign n211 = i_9_ & n210;
  assign n212 = ~i_15_ & n211;
  assign n213 = i_14_ & n212;
  assign n214 = n69 & n213;
  assign n215 = n209 & n214;
  assign n216 = ~i_8_ & n149;
  assign n217 = n65 & n216;
  assign n218 = n195 & n217;
  assign n219 = n68 & n192;
  assign n220 = n218 & n219;
  assign n221 = n134 & n199;
  assign n222 = n101 & n221;
  assign n223 = ~n220 & ~n222;
  assign n224 = ~n215 & n223;
  assign n225 = n97 & n190;
  assign n226 = n76 & n203;
  assign n227 = ~n221 & ~n226;
  assign n228 = n225 & ~n227;
  assign n229 = n224 & ~n228;
  assign n230 = ~n208 & n229;
  assign n231 = n76 & n199;
  assign n232 = ~i_7_ & n231;
  assign n233 = ~i_9_ & n210;
  assign n234 = ~i_15_ & n233;
  assign n235 = n97 & n234;
  assign n236 = n232 & n235;
  assign n237 = n141 & n202;
  assign n238 = ~i_8_ & n237;
  assign n239 = i_12_ & ~i_14_;
  assign n240 = n99 & n239;
  assign n241 = ~i_13_ & n240;
  assign n242 = ~i_15_ & n241;
  assign n243 = n238 & n242;
  assign n244 = n192 & n234;
  assign n245 = ~n119 & ~n244;
  assign n246 = n198 & ~n245;
  assign n247 = ~i_9_ & n188;
  assign n248 = ~i_15_ & n247;
  assign n249 = n97 & n248;
  assign n250 = n205 & n249;
  assign n251 = ~n246 & ~n250;
  assign n252 = ~n243 & n251;
  assign n253 = ~n236 & n252;
  assign n254 = n230 & n253;
  assign n255 = i_6_ & n203;
  assign n256 = i_8_ & n255;
  assign n257 = ~n114 & ~n119;
  assign n258 = ~n249 & n257;
  assign n259 = n256 & ~n258;
  assign n260 = n226 & n249;
  assign n261 = ~i_8_ & n197;
  assign n262 = n242 & n261;
  assign n263 = ~n260 & ~n262;
  assign n264 = ~n259 & n263;
  assign n265 = n254 & n264;
  assign n266 = n94 & n191;
  assign n267 = i_7_ & n231;
  assign n268 = n196 & n216;
  assign n269 = ~n218 & ~n268;
  assign n270 = ~n267 & n269;
  assign n271 = ~n261 & n270;
  assign n272 = n266 & ~n271;
  assign n273 = n192 & n211;
  assign n274 = ~i_15_ & n273;
  assign n275 = ~n242 & ~n274;
  assign n276 = ~n266 & n275;
  assign n277 = n198 & ~n276;
  assign n278 = ~n193 & ~n214;
  assign n279 = ~n274 & n278;
  assign n280 = ~n244 & n279;
  assign n281 = n261 & ~n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = n192 & n248;
  assign n284 = i_8_ & n221;
  assign n285 = ~i_6_ & n196;
  assign n286 = i_8_ & n285;
  assign n287 = ~i_7_ & n286;
  assign n288 = ~n284 & ~n287;
  assign n289 = ~n226 & n288;
  assign n290 = n283 & ~n289;
  assign n291 = n282 & ~n290;
  assign n292 = ~n272 & n291;
  assign n293 = ~n101 & ~n235;
  assign n294 = n256 & ~n293;
  assign n295 = ~i_8_ & n255;
  assign n296 = n118 & n192;
  assign n297 = ~n235 & ~n244;
  assign n298 = ~n296 & n297;
  assign n299 = n257 & n298;
  assign n300 = ~n101 & ~n225;
  assign n301 = ~n214 & n300;
  assign n302 = n299 & n301;
  assign n303 = n295 & ~n302;
  assign n304 = ~n294 & ~n303;
  assign n305 = ~n114 & ~n266;
  assign n306 = ~n100 & ~n190;
  assign n307 = n192 & ~n306;
  assign n308 = ~n274 & ~n307;
  assign n309 = ~i_8_ & n308;
  assign n310 = n305 & n309;
  assign n311 = ~n274 & n305;
  assign n312 = n298 & n311;
  assign n313 = i_8_ & n312;
  assign n314 = ~n310 & ~n313;
  assign n315 = n200 & n314;
  assign n316 = ~n114 & n298;
  assign n317 = n267 & ~n316;
  assign n318 = ~i_8_ & n200;
  assign n319 = ~n197 & ~n318;
  assign n320 = n296 & ~n319;
  assign n321 = ~n317 & ~n320;
  assign n322 = ~n315 & n321;
  assign n323 = n304 & n322;
  assign n324 = n292 & n323;
  assign n325 = n265 & n324;
  assign n326 = n68 & n97;
  assign n327 = i_8_ & n149;
  assign n328 = n196 & n327;
  assign n329 = ~n198 & ~n255;
  assign n330 = ~n328 & n329;
  assign n331 = n326 & ~n330;
  assign n332 = ~n198 & ~n200;
  assign n333 = n214 & ~n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~n226 & ~n238;
  assign n336 = n101 & ~n335;
  assign n337 = n114 & n197;
  assign n338 = ~n336 & ~n337;
  assign n339 = n119 & n284;
  assign n340 = n244 & n318;
  assign n341 = ~n339 & ~n340;
  assign n342 = n338 & n341;
  assign n343 = n334 & n342;
  assign n344 = i_7_ & n285;
  assign n345 = i_8_ & n344;
  assign n346 = n207 & ~n345;
  assign n347 = n201 & n242;
  assign n348 = n300 & ~n347;
  assign n349 = ~n346 & ~n348;
  assign n350 = n249 & ~n288;
  assign n351 = ~n274 & ~n296;
  assign n352 = ~n283 & n351;
  assign n353 = n256 & ~n352;
  assign n354 = ~n249 & ~n266;
  assign n355 = n295 & ~n354;
  assign n356 = ~n353 & ~n355;
  assign n357 = ~n350 & n356;
  assign n358 = ~n349 & n357;
  assign n359 = n343 & n358;
  assign n360 = n226 & ~n278;
  assign n361 = ~i_6_ & n203;
  assign n362 = ~n219 & ~n242;
  assign n363 = n312 & n362;
  assign n364 = ~n119 & n363;
  assign n365 = n361 & ~n364;
  assign n366 = ~n360 & ~n365;
  assign n367 = n326 & n361;
  assign n368 = n366 & ~n367;
  assign n369 = ~n206 & n283;
  assign n370 = n149 & n199;
  assign n371 = i_8_ & n370;
  assign n372 = ~n198 & n288;
  assign n373 = n199 & n204;
  assign n374 = i_7_ & n373;
  assign n375 = ~n328 & ~n374;
  assign n376 = n372 & n375;
  assign n377 = ~n371 & n376;
  assign n378 = ~n249 & ~n283;
  assign n379 = n198 & ~n378;
  assign n380 = n326 & n373;
  assign n381 = ~n219 & ~n380;
  assign n382 = ~n379 & n381;
  assign n383 = ~n377 & ~n382;
  assign n384 = ~n369 & ~n383;
  assign n385 = n368 & n384;
  assign n386 = n359 & n385;
  assign n387 = n325 & n386;
  assign n388 = i_12_ & i_13_;
  assign n389 = i_14_ & n388;
  assign n390 = n190 & n389;
  assign n391 = ~n200 & ~n261;
  assign n392 = ~n344 & n391;
  assign n393 = n390 & ~n392;
  assign n394 = n213 & n388;
  assign n395 = n248 & n389;
  assign n396 = ~n394 & ~n395;
  assign n397 = n205 & ~n396;
  assign n398 = n234 & n389;
  assign n399 = i_7_ & ~i_8_;
  assign n400 = n285 & n399;
  assign n401 = ~n318 & ~n400;
  assign n402 = n398 & ~n401;
  assign n403 = n113 & n388;
  assign n404 = ~n398 & ~n403;
  assign n405 = n267 & ~n404;
  assign n406 = ~n402 & ~n405;
  assign n407 = ~n397 & n406;
  assign n408 = ~n393 & n407;
  assign n409 = i_14_ & n191;
  assign n410 = i_15_ & n233;
  assign n411 = n409 & n410;
  assign n412 = ~n398 & ~n411;
  assign n413 = n102 & n409;
  assign n414 = n412 & ~n413;
  assign n415 = n100 & n389;
  assign n416 = ~n394 & ~n415;
  assign n417 = i_15_ & n211;
  assign n418 = i_14_ & n417;
  assign n419 = n191 & n418;
  assign n420 = n118 & n389;
  assign n421 = ~n419 & ~n420;
  assign n422 = n416 & n421;
  assign n423 = n414 & n422;
  assign n424 = n232 & ~n423;
  assign n425 = i_8_ & n237;
  assign n426 = ~n411 & ~n413;
  assign n427 = ~n415 & n426;
  assign n428 = n425 & ~n427;
  assign n429 = i_15_ & n189;
  assign n430 = n409 & n429;
  assign n431 = n318 & n430;
  assign n432 = ~n428 & ~n431;
  assign n433 = ~n424 & n432;
  assign n434 = n408 & n433;
  assign n435 = n116 & n409;
  assign n436 = ~n420 & ~n435;
  assign n437 = n396 & n436;
  assign n438 = ~n390 & ~n415;
  assign n439 = n437 & n438;
  assign n440 = n284 & ~n439;
  assign n441 = ~n394 & ~n419;
  assign n442 = n201 & ~n441;
  assign n443 = i_15_ & n247;
  assign n444 = i_14_ & n443;
  assign n445 = n191 & n444;
  assign n446 = ~n430 & ~n445;
  assign n447 = n261 & ~n446;
  assign n448 = ~n442 & ~n447;
  assign n449 = ~n226 & ~n286;
  assign n450 = n395 & ~n449;
  assign n451 = ~n226 & ~n232;
  assign n452 = ~n390 & ~n430;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n450 & ~n453;
  assign n455 = n448 & n454;
  assign n456 = ~n440 & n455;
  assign n457 = n237 & n419;
  assign n458 = n121 & n409;
  assign n459 = ~n268 & ~n370;
  assign n460 = n458 & ~n459;
  assign n461 = ~n457 & ~n460;
  assign n462 = n68 & n389;
  assign n463 = n295 & n462;
  assign n464 = i_15_ & n67;
  assign n465 = n409 & n464;
  assign n466 = n370 & n465;
  assign n467 = ~n463 & ~n466;
  assign n468 = n461 & n467;
  assign n469 = n456 & n468;
  assign n470 = n434 & n469;
  assign n471 = ~n403 & ~n458;
  assign n472 = i_8_ & ~n436;
  assign n473 = n471 & ~n472;
  assign n474 = ~n413 & n473;
  assign n475 = n200 & ~n474;
  assign n476 = n201 & n398;
  assign n477 = n318 & ~n441;
  assign n478 = n201 & n430;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n476 & n479;
  assign n481 = ~n475 & n480;
  assign n482 = n396 & ~n403;
  assign n483 = ~n420 & n482;
  assign n484 = n256 & ~n483;
  assign n485 = n481 & ~n484;
  assign n486 = n256 & n398;
  assign n487 = ~n390 & n412;
  assign n488 = n436 & n487;
  assign n489 = n482 & n488;
  assign n490 = n295 & ~n489;
  assign n491 = n255 & n415;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n486 & n492;
  assign n494 = n485 & n493;
  assign n495 = n470 & n494;
  assign n496 = ~i_8_ & n285;
  assign n497 = ~i_7_ & n496;
  assign n498 = n451 & ~n497;
  assign n499 = ~n318 & n498;
  assign n500 = ~n435 & ~n445;
  assign n501 = ~n499 & ~n500;
  assign n502 = ~n411 & ~n430;
  assign n503 = n436 & n502;
  assign n504 = ~n419 & ~n458;
  assign n505 = ~n462 & ~n465;
  assign n506 = n504 & n505;
  assign n507 = n503 & n506;
  assign n508 = n198 & ~n507;
  assign n509 = n261 & n415;
  assign n510 = ~n508 & ~n509;
  assign n511 = n412 & ~n435;
  assign n512 = n441 & ~n458;
  assign n513 = n511 & n512;
  assign n514 = n261 & ~n513;
  assign n515 = n197 & n413;
  assign n516 = ~n514 & ~n515;
  assign n517 = n510 & n516;
  assign n518 = ~n501 & n517;
  assign n519 = ~i_7_ & n285;
  assign n520 = ~n238 & ~n519;
  assign n521 = ~n284 & n520;
  assign n522 = ~n200 & n521;
  assign n523 = n238 & n398;
  assign n524 = ~n411 & ~n523;
  assign n525 = ~n522 & ~n524;
  assign n526 = ~n200 & ~n345;
  assign n527 = n415 & ~n526;
  assign n528 = n328 & n462;
  assign n529 = ~n527 & ~n528;
  assign n530 = n232 & n395;
  assign n531 = ~n394 & ~n445;
  assign n532 = n400 & ~n531;
  assign n533 = n197 & n403;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n530 & n534;
  assign n536 = ~n345 & ~n497;
  assign n537 = n430 & ~n536;
  assign n538 = ~n344 & n449;
  assign n539 = n465 & ~n538;
  assign n540 = ~n537 & ~n539;
  assign n541 = n535 & n540;
  assign n542 = n529 & n541;
  assign n543 = ~n525 & n542;
  assign n544 = n518 & n543;
  assign n545 = n287 & n445;
  assign n546 = ~n445 & n505;
  assign n547 = n284 & ~n546;
  assign n548 = n328 & n465;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~n256 & ~n374;
  assign n551 = n462 & ~n550;
  assign n552 = ~n198 & ~n201;
  assign n553 = ~n395 & ~n445;
  assign n554 = ~n552 & ~n553;
  assign n555 = n205 & n445;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n551 & n556;
  assign n558 = n549 & n557;
  assign n559 = n201 & n465;
  assign n560 = n558 & ~n559;
  assign n561 = ~n545 & n560;
  assign n562 = n414 & ~n462;
  assign n563 = n421 & n562;
  assign n564 = n471 & n563;
  assign n565 = n361 & ~n564;
  assign n566 = ~n430 & ~n465;
  assign n567 = ~n435 & n566;
  assign n568 = n205 & ~n567;
  assign n569 = n226 & ~n416;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n565 & n570;
  assign n572 = n561 & n571;
  assign n573 = n544 & n572;
  assign n574 = n495 & n573;
  assign n575 = n118 & n409;
  assign n576 = ~n198 & ~n284;
  assign n577 = n89 & n196;
  assign n578 = ~n318 & ~n577;
  assign n579 = ~n232 & n578;
  assign n580 = ~n295 & n579;
  assign n581 = ~n267 & ~n400;
  assign n582 = ~n361 & n581;
  assign n583 = n580 & n582;
  assign n584 = n576 & n583;
  assign n585 = n575 & ~n584;
  assign n586 = n234 & n409;
  assign n587 = ~n256 & ~n284;
  assign n588 = ~n201 & n587;
  assign n589 = n583 & n588;
  assign n590 = n586 & ~n589;
  assign n591 = ~n585 & ~n590;
  assign n592 = n288 & ~n496;
  assign n593 = ~n232 & ~n345;
  assign n594 = n592 & n593;
  assign n595 = ~n256 & n594;
  assign n596 = ~n273 & ~n296;
  assign n597 = ~n594 & ~n596;
  assign n598 = ~n266 & ~n597;
  assign n599 = ~n595 & ~n598;
  assign n600 = n121 & n192;
  assign n601 = ~n197 & n594;
  assign n602 = ~n371 & n601;
  assign n603 = n600 & ~n602;
  assign n604 = ~n599 & ~n603;
  assign n605 = n591 & n604;
  assign n606 = n574 & n605;
  assign n607 = n387 & n606;
  assign n608 = i_14_ & n91;
  assign n609 = n115 & n608;
  assign n610 = ~i_15_ & n609;
  assign n611 = ~n119 & ~n610;
  assign n612 = ~n420 & n611;
  assign n613 = n113 & ~n191;
  assign n614 = n612 & ~n613;
  assign n615 = ~n191 & n213;
  assign n616 = n614 & ~n615;
  assign n617 = i_14_ & n234;
  assign n618 = ~n191 & n617;
  assign n619 = n616 & ~n618;
  assign n620 = n497 & ~n619;
  assign n621 = n287 & n586;
  assign n622 = n100 & n608;
  assign n623 = ~n101 & ~n622;
  assign n624 = ~n415 & n623;
  assign n625 = n100 & n409;
  assign n626 = n624 & ~n625;
  assign n627 = n497 & ~n626;
  assign n628 = n287 & ~n624;
  assign n629 = i_14_ & n190;
  assign n630 = ~n191 & n629;
  assign n631 = n287 & n630;
  assign n632 = ~n628 & ~n631;
  assign n633 = ~n627 & n632;
  assign n634 = ~n621 & n633;
  assign n635 = ~n620 & n634;
  assign n636 = n191 & n213;
  assign n637 = ~n201 & ~n261;
  assign n638 = n636 & ~n637;
  assign n639 = ~n221 & ~n638;
  assign n640 = ~i_13_ & n213;
  assign n641 = ~n613 & ~n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = n635 & ~n642;
  assign n644 = ~n268 & ~n371;
  assign n645 = n613 & ~n644;
  assign n646 = n266 & n371;
  assign n647 = n237 & n394;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n645 & n648;
  assign n650 = i_14_ & n68;
  assign n651 = ~n191 & n650;
  assign n652 = ~n113 & ~n651;
  assign n653 = n218 & ~n652;
  assign n654 = n649 & ~n653;
  assign n655 = n86 & n195;
  assign n656 = ~n134 & n655;
  assign n657 = ~n149 & n656;
  assign n658 = n98 & n657;
  assign n659 = n267 & ~n612;
  assign n660 = ~n658 & ~n659;
  assign n661 = n191 & ~n306;
  assign n662 = ~n274 & ~n413;
  assign n663 = ~n661 & n662;
  assign n664 = n295 & ~n663;
  assign n665 = i_8_ & n575;
  assign n666 = ~n625 & ~n665;
  assign n667 = n237 & ~n666;
  assign n668 = ~n664 & ~n667;
  assign n669 = n660 & n668;
  assign n670 = n654 & n669;
  assign n671 = ~n267 & n594;
  assign n672 = n458 & ~n671;
  assign n673 = n256 & ~n426;
  assign n674 = n446 & n504;
  assign n675 = ~n219 & n674;
  assign n676 = n255 & ~n675;
  assign n677 = ~n673 & ~n676;
  assign n678 = ~n672 & n677;
  assign n679 = n670 & n678;
  assign n680 = n643 & n679;
  assign n681 = n248 & n409;
  assign n682 = ~n198 & n587;
  assign n683 = n681 & ~n682;
  assign n684 = n371 & n650;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n575 & ~n636;
  assign n687 = ~n651 & n686;
  assign n688 = n619 & n687;
  assign n689 = n287 & ~n688;
  assign n690 = n685 & ~n689;
  assign n691 = n113 & n191;
  assign n692 = n295 & n691;
  assign n693 = n256 & n630;
  assign n694 = n295 & n681;
  assign n695 = ~n693 & ~n694;
  assign n696 = n190 & n409;
  assign n697 = ~n636 & ~n696;
  assign n698 = n256 & ~n697;
  assign n699 = n695 & ~n698;
  assign n700 = ~n692 & n699;
  assign n701 = n232 & n610;
  assign n702 = n238 & n575;
  assign n703 = ~n701 & ~n702;
  assign n704 = n438 & ~n691;
  assign n705 = n205 & ~n704;
  assign n706 = ~n205 & ~n318;
  assign n707 = n625 & ~n706;
  assign n708 = ~n705 & ~n707;
  assign n709 = n703 & n708;
  assign n710 = n700 & n709;
  assign n711 = ~n197 & ~n201;
  assign n712 = n451 & n711;
  assign n713 = ~n256 & ~n287;
  assign n714 = ~n345 & n713;
  assign n715 = n712 & n714;
  assign n716 = n625 & ~n715;
  assign n717 = ~n295 & ~n496;
  assign n718 = ~n198 & ~n361;
  assign n719 = n717 & n718;
  assign n720 = ~n318 & n719;
  assign n721 = n636 & ~n720;
  assign n722 = ~n201 & ~n256;
  assign n723 = n575 & ~n722;
  assign n724 = n438 & ~n617;
  assign n725 = ~n394 & n724;
  assign n726 = n198 & ~n725;
  assign n727 = ~n723 & ~n726;
  assign n728 = ~n721 & n727;
  assign n729 = ~n716 & n728;
  assign n730 = n710 & n729;
  assign n731 = n690 & n730;
  assign n732 = n680 & n731;
  assign n733 = n68 & n409;
  assign n734 = ~n201 & ~n345;
  assign n735 = ~n261 & ~n318;
  assign n736 = ~n496 & n735;
  assign n737 = ~n232 & n736;
  assign n738 = n734 & n737;
  assign n739 = n372 & n738;
  assign n740 = ~n203 & n739;
  assign n741 = ~n218 & n375;
  assign n742 = n740 & n741;
  assign n743 = n733 & ~n742;
  assign n744 = n691 & ~n739;
  assign n745 = ~n244 & ~n307;
  assign n746 = ~n595 & ~n745;
  assign n747 = ~n744 & ~n746;
  assign n748 = ~n743 & n747;
  assign n749 = n614 & n626;
  assign n750 = n400 & ~n749;
  assign n751 = n616 & n686;
  assign n752 = ~n617 & n751;
  assign n753 = n345 & ~n752;
  assign n754 = ~n750 & ~n753;
  assign n755 = n592 & n735;
  assign n756 = n346 & n755;
  assign n757 = n451 & n756;
  assign n758 = n696 & ~n757;
  assign n759 = n248 & n608;
  assign n760 = ~n249 & ~n759;
  assign n761 = ~n734 & ~n760;
  assign n762 = ~n497 & ~n761;
  assign n763 = ~n395 & n760;
  assign n764 = ~n630 & n763;
  assign n765 = ~n762 & ~n764;
  assign n766 = ~n261 & n401;
  assign n767 = ~i_12_ & n617;
  assign n768 = n763 & ~n767;
  assign n769 = ~n766 & ~n768;
  assign n770 = ~n765 & ~n769;
  assign n771 = ~n413 & ~n419;
  assign n772 = ~n430 & n771;
  assign n773 = ~n618 & ~n625;
  assign n774 = n772 & n773;
  assign n775 = n284 & ~n774;
  assign n776 = n219 & ~n738;
  assign n777 = ~n775 & ~n776;
  assign n778 = n770 & n777;
  assign n779 = ~n758 & n778;
  assign n780 = n754 & n779;
  assign n781 = n748 & n780;
  assign n782 = n732 & n781;
  assign n783 = i_15_ & n273;
  assign n784 = ~n610 & ~n783;
  assign n785 = n190 & n608;
  assign n786 = i_15_ & n241;
  assign n787 = n192 & n429;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~n785 & n788;
  assign n790 = ~n622 & n789;
  assign n791 = n211 & n608;
  assign n792 = ~i_15_ & n791;
  assign n793 = i_12_ & n443;
  assign n794 = ~i_14_ & n793;
  assign n795 = ~i_13_ & n794;
  assign n796 = ~n792 & ~n795;
  assign n797 = n91 & n113;
  assign n798 = n116 & n239;
  assign n799 = ~i_13_ & n798;
  assign n800 = ~n797 & ~n799;
  assign n801 = n796 & n800;
  assign n802 = n790 & n801;
  assign n803 = n784 & n802;
  assign n804 = n295 & ~n803;
  assign n805 = ~i_14_ & n410;
  assign n806 = n191 & n805;
  assign n807 = n234 & n608;
  assign n808 = ~n806 & ~n807;
  assign n809 = n255 & ~n808;
  assign n810 = n68 & n608;
  assign n811 = ~n786 & ~n810;
  assign n812 = ~n622 & n811;
  assign n813 = n256 & ~n812;
  assign n814 = ~n809 & ~n813;
  assign n815 = ~n804 & n814;
  assign n816 = ~n759 & ~n795;
  assign n817 = ~n785 & n816;
  assign n818 = n226 & ~n817;
  assign n819 = n610 & ~n682;
  assign n820 = n198 & n759;
  assign n821 = n192 & n464;
  assign n822 = ~n810 & ~n821;
  assign n823 = n373 & ~n822;
  assign n824 = ~n820 & ~n823;
  assign n825 = n201 & n795;
  assign n826 = n328 & n821;
  assign n827 = ~n825 & ~n826;
  assign n828 = n824 & n827;
  assign n829 = n256 & ~n801;
  assign n830 = n828 & ~n829;
  assign n831 = ~n819 & n830;
  assign n832 = ~n818 & n831;
  assign n833 = n815 & n832;
  assign n834 = ~n600 & ~n797;
  assign n835 = n808 & n834;
  assign n836 = n267 & ~n835;
  assign n837 = ~n209 & n711;
  assign n838 = n783 & ~n837;
  assign n839 = ~n836 & ~n838;
  assign n840 = n232 & ~n808;
  assign n841 = n295 & n810;
  assign n842 = ~n706 & n795;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n840 & n843;
  assign n845 = n201 & n799;
  assign n846 = n318 & n783;
  assign n847 = ~n845 & ~n846;
  assign n848 = n201 & ~n808;
  assign n849 = n200 & ~n834;
  assign n850 = ~n848 & ~n849;
  assign n851 = n847 & n850;
  assign n852 = n844 & n851;
  assign n853 = n839 & n852;
  assign n854 = n255 & n600;
  assign n855 = n790 & ~n792;
  assign n856 = n221 & ~n855;
  assign n857 = ~n209 & ~n284;
  assign n858 = n759 & ~n857;
  assign n859 = n261 & n792;
  assign n860 = ~n787 & ~n792;
  assign n861 = n205 & ~n860;
  assign n862 = ~n859 & ~n861;
  assign n863 = ~n858 & n862;
  assign n864 = ~n856 & n863;
  assign n865 = ~n854 & n864;
  assign n866 = n853 & n865;
  assign n867 = n833 & n866;
  assign n868 = n205 & n821;
  assign n869 = ~n610 & n811;
  assign n870 = ~n799 & n869;
  assign n871 = n835 & n870;
  assign n872 = n361 & ~n871;
  assign n873 = ~n783 & ~n792;
  assign n874 = n226 & ~n873;
  assign n875 = n226 & n787;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n872 & n876;
  assign n878 = ~n868 & n877;
  assign n879 = n226 & n821;
  assign n880 = n878 & ~n879;
  assign n881 = n718 & n734;
  assign n882 = n205 & n785;
  assign n883 = ~n622 & ~n882;
  assign n884 = ~n881 & ~n883;
  assign n885 = ~n198 & n734;
  assign n886 = ~n789 & ~n885;
  assign n887 = n425 & n622;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n329 & n821;
  assign n890 = ~n269 & n600;
  assign n891 = ~n198 & ~n318;
  assign n892 = n799 & ~n891;
  assign n893 = ~n890 & ~n892;
  assign n894 = ~n198 & ~n328;
  assign n895 = n810 & ~n894;
  assign n896 = n893 & ~n895;
  assign n897 = ~n889 & n896;
  assign n898 = ~n200 & ~n400;
  assign n899 = ~n198 & n898;
  assign n900 = n792 & ~n899;
  assign n901 = ~n287 & ~n295;
  assign n902 = n759 & ~n901;
  assign n903 = ~n900 & ~n902;
  assign n904 = n197 & n797;
  assign n905 = n238 & n786;
  assign n906 = ~n904 & ~n905;
  assign n907 = n903 & n906;
  assign n908 = n897 & n907;
  assign n909 = n888 & n908;
  assign n910 = ~n884 & n909;
  assign n911 = n880 & n910;
  assign n912 = n867 & n911;
  assign n913 = ~n201 & ~n286;
  assign n914 = n737 & n913;
  assign n915 = ~n370 & n914;
  assign n916 = n821 & ~n915;
  assign n917 = ~n119 & n760;
  assign n918 = n232 & ~n917;
  assign n919 = n612 & ~n799;
  assign n920 = ~n296 & ~n435;
  assign n921 = n919 & n920;
  assign n922 = n237 & ~n921;
  assign n923 = ~n413 & ~n415;
  assign n924 = n238 & ~n923;
  assign n925 = n238 & n622;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n922 & n926;
  assign n928 = ~n287 & ~n400;
  assign n929 = n430 & ~n928;
  assign n930 = ~n267 & ~n344;
  assign n931 = n411 & ~n930;
  assign n932 = ~n929 & ~n931;
  assign n933 = n927 & n932;
  assign n934 = ~n918 & n933;
  assign n935 = ~n916 & n934;
  assign n936 = ~n361 & n914;
  assign n937 = n681 & ~n936;
  assign n938 = ~n255 & n579;
  assign n939 = ~n374 & n938;
  assign n940 = n465 & ~n939;
  assign n941 = ~n519 & n766;
  assign n942 = ~n623 & ~n735;
  assign n943 = n214 & n400;
  assign n944 = n788 & ~n943;
  assign n945 = ~n942 & n944;
  assign n946 = ~n941 & ~n945;
  assign n947 = ~n940 & ~n946;
  assign n948 = ~n937 & n947;
  assign n949 = n935 & n948;
  assign n950 = ~n256 & ~n267;
  assign n951 = n644 & n950;
  assign n952 = ~n226 & n951;
  assign n953 = n691 & ~n952;
  assign n954 = n256 & n787;
  assign n955 = ~n953 & ~n954;
  assign n956 = n651 & ~n738;
  assign n957 = n285 & ~n771;
  assign n958 = ~i_12_ & n629;
  assign n959 = ~n766 & n958;
  assign n960 = ~n957 & ~n959;
  assign n961 = ~n956 & n960;
  assign n962 = n955 & n961;
  assign n963 = ~n671 & n799;
  assign n964 = ~n344 & n580;
  assign n965 = n283 & ~n964;
  assign n966 = ~n963 & ~n965;
  assign n967 = n962 & n966;
  assign n968 = n345 & n445;
  assign n969 = ~n101 & ~n241;
  assign n970 = n425 & ~n969;
  assign n971 = ~n968 & ~n970;
  assign n972 = n713 & n930;
  assign n973 = n435 & ~n972;
  assign n974 = ~n149 & n196;
  assign n975 = ~n284 & ~n318;
  assign n976 = ~n974 & n975;
  assign n977 = n806 & ~n976;
  assign n978 = ~n973 & ~n977;
  assign n979 = ~i_8_ & n420;
  assign n980 = n611 & ~n979;
  assign n981 = n200 & ~n980;
  assign n982 = n398 & n425;
  assign n983 = ~n981 & ~n982;
  assign n984 = n261 & ~n919;
  assign n985 = n983 & ~n984;
  assign n986 = n978 & n985;
  assign n987 = n971 & n986;
  assign n988 = ~n601 & n795;
  assign n989 = n987 & ~n988;
  assign n990 = n967 & n989;
  assign n991 = n949 & n990;
  assign n992 = n912 & n991;
  assign n993 = n782 & n992;
  assign n994 = n607 & n993;
  assign o_5_ = ~n175 | ~n994;
  assign n996 = n63 & n65;
  assign n997 = ~n153 & ~n996;
  assign o_6_ = ~n148 | ~n997;
  assign n999 = i_13_ & n798;
  assign n1000 = i_14_ & ~n388;
  assign n1001 = n116 & n1000;
  assign n1002 = n410 & n1000;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~n999 & n1003;
  assign n1005 = n267 & ~n1004;
  assign n1006 = n398 & ~n536;
  assign n1007 = n97 & n102;
  assign n1008 = ~n451 & n1007;
  assign n1009 = n389 & n429;
  assign n1010 = n295 & n1009;
  assign n1011 = ~n1008 & ~n1010;
  assign n1012 = ~n1006 & n1011;
  assign n1013 = ~n1005 & n1012;
  assign n1014 = n97 & n121;
  assign n1015 = ~n200 & ~n232;
  assign n1016 = ~n577 & n1015;
  assign n1017 = n372 & n1016;
  assign n1018 = n1014 & ~n1017;
  assign n1019 = i_14_ & n121;
  assign n1020 = ~n388 & n1019;
  assign n1021 = ~n950 & n1020;
  assign n1022 = n395 & ~n736;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n1018 & n1023;
  assign n1025 = n388 & n418;
  assign n1026 = n1003 & ~n1025;
  assign n1027 = ~n388 & n444;
  assign n1028 = i_14_ & n429;
  assign n1029 = n464 & n1000;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~n1027 & n1030;
  assign n1032 = n1026 & n1031;
  assign n1033 = n256 & ~n1032;
  assign n1034 = ~n388 & n418;
  assign n1035 = n429 & n1000;
  assign n1036 = ~n444 & ~n1035;
  assign n1037 = ~n1020 & n1036;
  assign n1038 = ~n1034 & n1037;
  assign n1039 = n295 & ~n1038;
  assign n1040 = n102 & n1000;
  assign n1041 = n255 & n1040;
  assign n1042 = ~n1039 & ~n1041;
  assign n1043 = ~n1033 & n1042;
  assign n1044 = n388 & n805;
  assign n1045 = ~n976 & n1044;
  assign n1046 = n1043 & ~n1045;
  assign n1047 = n1024 & n1046;
  assign n1048 = n97 & n410;
  assign n1049 = ~n398 & ~n1044;
  assign n1050 = ~n1048 & n1049;
  assign n1051 = n425 & ~n1050;
  assign n1052 = n198 & n1009;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = n256 & n1034;
  assign n1055 = n287 & n1034;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n1053 & n1056;
  assign n1058 = n1047 & n1057;
  assign n1059 = n1013 & n1058;
  assign n1060 = n459 & n594;
  assign n1061 = n403 & ~n1060;
  assign n1062 = ~i_14_ & n388;
  assign n1063 = n247 & n1062;
  assign n1064 = ~i_15_ & n1063;
  assign n1065 = n226 & n1064;
  assign n1066 = ~n459 & n1014;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~i_15_ & n1062;
  assign n1069 = n361 & n1068;
  assign n1070 = ~i_8_ & n247;
  assign n1071 = n1069 & ~n1070;
  assign n1072 = n1067 & ~n1071;
  assign n1073 = n68 & n1062;
  assign n1074 = n374 & n1073;
  assign n1075 = n238 & n1048;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = n1072 & n1076;
  assign n1078 = ~n328 & ~n370;
  assign n1079 = n97 & n464;
  assign n1080 = ~n1073 & ~n1079;
  assign n1081 = ~n1078 & ~n1080;
  assign n1082 = n92 & n1062;
  assign n1083 = ~i_15_ & n1082;
  assign n1084 = ~n267 & ~n1083;
  assign n1085 = n233 & n1068;
  assign n1086 = n118 & n1062;
  assign n1087 = ~n1083 & ~n1086;
  assign n1088 = ~n1085 & n1087;
  assign n1089 = ~n1084 & ~n1088;
  assign n1090 = ~n270 & n1089;
  assign n1091 = n237 & n1068;
  assign n1092 = n210 & n1091;
  assign n1093 = ~n1090 & ~n1092;
  assign n1094 = ~n1081 & n1093;
  assign n1095 = n1077 & n1094;
  assign n1096 = n97 & n417;
  assign n1097 = ~n394 & ~n1096;
  assign n1098 = n388 & n417;
  assign n1099 = n1097 & ~n1098;
  assign n1100 = n237 & ~n1099;
  assign n1101 = ~n69 & n1020;
  assign n1102 = n438 & ~n1101;
  assign n1103 = n519 & ~n1102;
  assign n1104 = ~n1100 & ~n1103;
  assign n1105 = n1095 & n1104;
  assign n1106 = ~n1061 & n1105;
  assign n1107 = n102 & n389;
  assign n1108 = n1088 & ~n1107;
  assign n1109 = i_9_ & n1068;
  assign n1110 = ~n66 & n1109;
  assign n1111 = ~n1064 & ~n1110;
  assign n1112 = ~n1073 & n1111;
  assign n1113 = n1108 & n1112;
  assign n1114 = n255 & ~n1113;
  assign n1115 = ~n237 & ~n267;
  assign n1116 = ~n345 & n1115;
  assign n1117 = n420 & ~n1116;
  assign n1118 = ~n1114 & ~n1117;
  assign n1119 = n464 & n1062;
  assign n1120 = ~n462 & ~n1119;
  assign n1121 = ~n915 & ~n1120;
  assign n1122 = n102 & n1062;
  assign n1123 = n429 & n1062;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = ~n420 & n1124;
  assign n1126 = ~n941 & ~n1125;
  assign n1127 = n97 & n429;
  assign n1128 = ~n498 & n1127;
  assign n1129 = ~n1126 & ~n1128;
  assign n1130 = ~n1121 & n1129;
  assign n1131 = n1118 & n1130;
  assign n1132 = n1106 & n1131;
  assign n1133 = ~n267 & n740;
  assign n1134 = n121 & n389;
  assign n1135 = ~i_14_ & n1098;
  assign n1136 = ~n999 & ~n1135;
  assign n1137 = n388 & n443;
  assign n1138 = n1113 & ~n1137;
  assign n1139 = n1136 & n1138;
  assign n1140 = ~n739 & ~n1139;
  assign n1141 = n389 & n410;
  assign n1142 = n116 & n389;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n1140 & n1143;
  assign n1145 = ~n1134 & n1144;
  assign n1146 = ~n1133 & ~n1145;
  assign n1147 = n1132 & ~n1146;
  assign n1148 = n1059 & n1147;
  assign n1149 = ~n1044 & ~n1122;
  assign n1150 = n256 & ~n1149;
  assign n1151 = i_15_ & n1063;
  assign n1152 = n1124 & ~n1151;
  assign n1153 = i_15_ & n609;
  assign n1154 = n410 & n608;
  assign n1155 = ~n1044 & ~n1154;
  assign n1156 = ~n1153 & n1155;
  assign n1157 = n1136 & n1156;
  assign n1158 = n1152 & n1157;
  assign n1159 = n295 & ~n1158;
  assign n1160 = ~n1150 & ~n1159;
  assign n1161 = ~n375 & n1119;
  assign n1162 = n91 & n444;
  assign n1163 = ~n284 & n552;
  assign n1164 = n1162 & ~n1163;
  assign n1165 = ~n1161 & ~n1164;
  assign n1166 = n464 & n608;
  assign n1167 = ~n894 & n1166;
  assign n1168 = ~n1119 & ~n1166;
  assign n1169 = n284 & ~n1168;
  assign n1170 = ~n1167 & ~n1169;
  assign n1171 = n1165 & n1170;
  assign n1172 = n121 & n608;
  assign n1173 = ~n1154 & ~n1172;
  assign n1174 = ~n1153 & n1173;
  assign n1175 = n102 & n608;
  assign n1176 = i_15_ & n791;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = n1174 & n1177;
  assign n1179 = n261 & ~n1178;
  assign n1180 = n232 & n1175;
  assign n1181 = ~n459 & n1172;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~n1179 & n1182;
  assign n1184 = n1171 & n1183;
  assign n1185 = n425 & n1154;
  assign n1186 = n91 & n1028;
  assign n1187 = ~n1176 & ~n1186;
  assign n1188 = n1155 & n1187;
  assign n1189 = n200 & n1186;
  assign n1190 = ~n232 & ~n1189;
  assign n1191 = ~n1188 & ~n1190;
  assign n1192 = ~n198 & ~n1153;
  assign n1193 = ~n576 & ~n1174;
  assign n1194 = ~n1192 & n1193;
  assign n1195 = i_15_ & n1082;
  assign n1196 = n255 & n1195;
  assign n1197 = ~n1194 & ~n1196;
  assign n1198 = ~n1191 & n1197;
  assign n1199 = ~n1185 & n1198;
  assign n1200 = n1184 & n1199;
  assign n1201 = n1160 & n1200;
  assign n1202 = ~n1135 & ~n1151;
  assign n1203 = n209 & ~n1202;
  assign n1204 = n221 & ~n1124;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n1044 & ~n1195;
  assign n1207 = n267 & ~n1206;
  assign n1208 = ~n1162 & ~n1186;
  assign n1209 = n261 & ~n1208;
  assign n1210 = n370 & n1166;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1207 & n1211;
  assign n1213 = n1205 & n1212;
  assign n1214 = n201 & ~n1156;
  assign n1215 = n201 & n1166;
  assign n1216 = ~n1172 & ~n1175;
  assign n1217 = ~n1195 & n1216;
  assign n1218 = n200 & ~n1217;
  assign n1219 = n318 & n1176;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~n1215 & n1220;
  assign n1222 = ~n1214 & n1221;
  assign n1223 = ~n1162 & ~n1176;
  assign n1224 = n205 & ~n1223;
  assign n1225 = n256 & n999;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~n201 & ~n237;
  assign n1228 = n1176 & ~n1227;
  assign n1229 = ~n1123 & ~n1186;
  assign n1230 = ~n1151 & n1229;
  assign n1231 = n226 & ~n1230;
  assign n1232 = ~n1228 & ~n1231;
  assign n1233 = n1226 & n1232;
  assign n1234 = n1222 & n1233;
  assign n1235 = n1213 & n1234;
  assign n1236 = n1201 & n1235;
  assign n1237 = ~n881 & n1122;
  assign n1238 = ~n538 & n1166;
  assign n1239 = n520 & n975;
  assign n1240 = n1154 & ~n1239;
  assign n1241 = ~n1238 & ~n1240;
  assign n1242 = ~n1237 & n1241;
  assign n1243 = n499 & n928;
  assign n1244 = n1162 & ~n1243;
  assign n1245 = ~n536 & n1186;
  assign n1246 = ~n329 & n1119;
  assign n1247 = ~n269 & n1195;
  assign n1248 = n238 & n1044;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~n1246 & n1249;
  assign n1251 = ~n1245 & n1250;
  assign n1252 = ~n1244 & n1251;
  assign n1253 = n1242 & n1252;
  assign n1254 = ~n1153 & n1168;
  assign n1255 = n205 & ~n1254;
  assign n1256 = n1155 & ~n1195;
  assign n1257 = ~n999 & n1256;
  assign n1258 = n361 & ~n1257;
  assign n1259 = ~n1135 & n1177;
  assign n1260 = n226 & ~n1259;
  assign n1261 = ~n1258 & ~n1260;
  assign n1262 = ~n1255 & n1261;
  assign n1263 = ~i_8_ & n1119;
  assign n1264 = ~n1172 & ~n1263;
  assign n1265 = n361 & ~n1264;
  assign n1266 = n1262 & ~n1265;
  assign n1267 = ~n499 & n1153;
  assign n1268 = ~n346 & n1123;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = n1266 & n1269;
  assign n1271 = n1253 & n1270;
  assign n1272 = n1236 & n1271;
  assign n1273 = ~n374 & n740;
  assign n1274 = n1078 & n1273;
  assign n1275 = n389 & n464;
  assign n1276 = ~n1274 & n1275;
  assign n1277 = ~n201 & n580;
  assign n1278 = n1048 & ~n1277;
  assign n1279 = ~n1025 & ~n1278;
  assign n1280 = ~n198 & n1277;
  assign n1281 = ~n400 & n1280;
  assign n1282 = ~n1279 & ~n1281;
  assign n1283 = ~n295 & n739;
  assign n1284 = n1079 & ~n1283;
  assign n1285 = ~n602 & n1195;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1282 & n1286;
  assign n1288 = ~n1276 & n1287;
  assign n1289 = n1272 & n1288;
  assign n1290 = ~n390 & ~n1186;
  assign n1291 = ~n1127 & n1290;
  assign n1292 = ~n415 & ~n1175;
  assign n1293 = ~n1007 & n1292;
  assign n1294 = n1291 & n1293;
  assign n1295 = i_8_ & ~n1294;
  assign n1296 = n97 & n116;
  assign n1297 = ~n1014 & ~n1048;
  assign n1298 = ~n1296 & n1297;
  assign n1299 = ~n1295 & n1298;
  assign n1300 = n69 & n444;
  assign n1301 = n388 & n444;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~n1009 & ~n1079;
  assign n1304 = ~n1096 & ~n1107;
  assign n1305 = n1303 & n1304;
  assign n1306 = n1302 & n1305;
  assign n1307 = n1299 & n1306;
  assign n1308 = ~n1025 & n1307;
  assign n1309 = n361 & ~n1308;
  assign n1310 = ~n1035 & ~n1040;
  assign n1311 = ~n1025 & n1310;
  assign n1312 = ~n1001 & n1311;
  assign n1313 = n287 & ~n1312;
  assign n1314 = ~n1034 & ~n1040;
  assign n1315 = n497 & ~n1314;
  assign n1316 = ~n1313 & ~n1315;
  assign n1317 = ~n390 & ~n1123;
  assign n1318 = n256 & ~n1317;
  assign n1319 = n232 & n1096;
  assign n1320 = n371 & n1083;
  assign n1321 = ~n924 & ~n1320;
  assign n1322 = ~n1319 & n1321;
  assign n1323 = ~n459 & n1134;
  assign n1324 = n1322 & ~n1323;
  assign n1325 = ~n1040 & ~n1127;
  assign n1326 = n345 & ~n1325;
  assign n1327 = ~n1007 & ~n1096;
  assign n1328 = ~n1127 & n1327;
  assign n1329 = ~n391 & ~n1328;
  assign n1330 = ~n435 & ~n1141;
  assign n1331 = n237 & ~n1330;
  assign n1332 = n284 & n1034;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1329 & n1333;
  assign n1335 = ~n1326 & n1334;
  assign n1336 = n1324 & n1335;
  assign n1337 = ~n1318 & n1336;
  assign n1338 = n1316 & n1337;
  assign n1339 = ~n1309 & n1338;
  assign n1340 = ~i_8_ & ~n1314;
  assign n1341 = i_8_ & n418;
  assign n1342 = n1003 & ~n1341;
  assign n1343 = ~n1340 & n1342;
  assign n1344 = ~n1020 & n1343;
  assign n1345 = n344 & ~n1344;
  assign n1346 = n284 & ~n1311;
  assign n1347 = n221 & n1101;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1345 & n1348;
  assign n1350 = n1097 & ~n1176;
  assign n1351 = n1294 & n1350;
  assign n1352 = n198 & ~n1351;
  assign n1353 = ~n286 & ~n519;
  assign n1354 = n394 & ~n1353;
  assign n1355 = n210 & n657;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = ~n415 & ~n1035;
  assign n1358 = n400 & ~n1357;
  assign n1359 = n1356 & ~n1358;
  assign n1360 = ~n1352 & n1359;
  assign n1361 = n1349 & n1360;
  assign n1362 = n580 & n1163;
  assign n1363 = n1296 & ~n1362;
  assign n1364 = ~n1048 & ~n1300;
  assign n1365 = ~n398 & n1364;
  assign n1366 = ~n372 & ~n1365;
  assign n1367 = n345 & n1027;
  assign n1368 = n256 & n1301;
  assign n1369 = n374 & n1029;
  assign n1370 = n201 & n1300;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1368 & n1371;
  assign n1373 = ~n1367 & n1372;
  assign n1374 = ~n1366 & n1373;
  assign n1375 = ~n1363 & n1374;
  assign n1376 = ~n465 & ~n1166;
  assign n1377 = ~n580 & ~n1376;
  assign n1378 = ~n737 & n1300;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = ~n284 & n914;
  assign n1381 = n1009 & ~n1380;
  assign n1382 = n1379 & ~n1381;
  assign n1383 = n1375 & n1382;
  assign n1384 = n1361 & n1383;
  assign n1385 = n1339 & n1384;
  assign n1386 = n574 & n1385;
  assign n1387 = n1289 & n1386;
  assign o_7_ = ~n1148 | ~n1387;
  assign o_8_ = i_3_ & n194;
  assign n1390 = n70 & n464;
  assign n1391 = ~n587 & n1390;
  assign n1392 = n68 & n105;
  assign n1393 = ~n375 & n1390;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n377 & ~n1394;
  assign n1396 = n105 & n248;
  assign n1397 = n70 & n443;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = n205 & n1396;
  assign n1400 = n552 & ~n1399;
  assign n1401 = ~n1398 & ~n1400;
  assign n1402 = ~n1395 & ~n1401;
  assign n1403 = ~n1391 & n1402;
  assign n1404 = ~i_14_ & ~n91;
  assign n1405 = n464 & n1404;
  assign n1406 = ~n810 & ~n1405;
  assign n1407 = ~n326 & n1406;
  assign n1408 = n198 & ~n1407;
  assign n1409 = n287 & ~n1376;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = n384 & n1410;
  assign n1412 = n1403 & n1411;
  assign n1413 = n69 & n805;
  assign n1414 = ~n103 & ~n1413;
  assign n1415 = n256 & ~n1414;
  assign n1416 = n105 & n234;
  assign n1417 = ~n1413 & ~n1416;
  assign n1418 = n70 & n429;
  assign n1419 = ~n103 & ~n1418;
  assign n1420 = n70 & n417;
  assign n1421 = n1419 & ~n1420;
  assign n1422 = ~n117 & ~n1397;
  assign n1423 = n1421 & n1422;
  assign n1424 = n1417 & n1423;
  assign n1425 = n295 & ~n1424;
  assign n1426 = ~n1415 & ~n1425;
  assign n1427 = ~n95 & ~n106;
  assign n1428 = n198 & ~n1427;
  assign n1429 = ~i_14_ & n212;
  assign n1430 = n91 & n1429;
  assign n1431 = n197 & n1430;
  assign n1432 = n105 & n190;
  assign n1433 = ~n1416 & ~n1432;
  assign n1434 = n261 & ~n1433;
  assign n1435 = ~n1431 & ~n1434;
  assign n1436 = ~n1428 & n1435;
  assign n1437 = ~n117 & n1419;
  assign n1438 = n232 & ~n1437;
  assign n1439 = n124 & n1417;
  assign n1440 = n231 & n1413;
  assign n1441 = ~n267 & ~n1440;
  assign n1442 = ~n1439 & ~n1441;
  assign n1443 = ~n1438 & ~n1442;
  assign n1444 = n1436 & n1443;
  assign n1445 = n1426 & n1444;
  assign n1446 = ~n205 & n288;
  assign n1447 = n284 & ~n1437;
  assign n1448 = ~n1397 & ~n1447;
  assign n1449 = ~n1446 & ~n1448;
  assign n1450 = n201 & n1432;
  assign n1451 = n122 & n255;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = n106 & n261;
  assign n1454 = n1452 & ~n1453;
  assign n1455 = ~n1449 & n1454;
  assign n1456 = n1445 & n1455;
  assign n1457 = ~n288 & n1396;
  assign n1458 = n218 & n1392;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n221 & n837;
  assign n1461 = n1420 & ~n1460;
  assign n1462 = n226 & ~n1398;
  assign n1463 = ~n1418 & ~n1432;
  assign n1464 = n205 & ~n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1466 = n95 & ~n271;
  assign n1467 = n1465 & ~n1466;
  assign n1468 = ~n1461 & n1467;
  assign n1469 = ~n123 & n1433;
  assign n1470 = n198 & ~n1469;
  assign n1471 = n256 & ~n1422;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = n295 & n1390;
  assign n1474 = n1472 & ~n1473;
  assign n1475 = n1468 & n1474;
  assign n1476 = n1459 & n1475;
  assign n1477 = n1456 & n1476;
  assign n1478 = n1236 & n1477;
  assign n1479 = n325 & n1478;
  assign n1480 = n1412 & n1479;
  assign n1481 = ~n1420 & n1463;
  assign n1482 = ~i_8_ & ~n1481;
  assign n1483 = ~n95 & ~n1430;
  assign n1484 = ~n122 & n1483;
  assign n1485 = n107 & n1484;
  assign n1486 = ~n1482 & n1485;
  assign n1487 = ~n123 & n1417;
  assign n1488 = ~n117 & n1487;
  assign n1489 = ~n1390 & ~n1392;
  assign n1490 = n1488 & n1489;
  assign n1491 = n1486 & n1490;
  assign n1492 = n361 & ~n1491;
  assign n1493 = ~n958 & ~n1123;
  assign n1494 = n205 & ~n1493;
  assign n1495 = ~n1492 & ~n1494;
  assign n1496 = n623 & ~n1122;
  assign n1497 = n361 & ~n1496;
  assign n1498 = n571 & ~n1497;
  assign n1499 = n1495 & n1498;
  assign n1500 = n366 & n1499;
  assign n1501 = ~n123 & ~n1396;
  assign n1502 = n1376 & n1501;
  assign n1503 = ~n283 & n1502;
  assign n1504 = ~n964 & ~n1503;
  assign n1505 = n105 & n116;
  assign n1506 = ~n584 & n1505;
  assign n1507 = n91 & n805;
  assign n1508 = ~n589 & n1507;
  assign n1509 = ~n1506 & ~n1508;
  assign n1510 = ~n1504 & n1509;
  assign n1511 = ~n326 & ~n1390;
  assign n1512 = n1120 & n1511;
  assign n1513 = n822 & n1512;
  assign n1514 = ~n738 & ~n1513;
  assign n1515 = n1510 & ~n1514;
  assign n1516 = n1500 & n1515;
  assign n1517 = n591 & n1516;
  assign n1518 = n867 & n1517;
  assign n1519 = n1480 & n1518;
  assign n1520 = n201 & ~n1488;
  assign n1521 = n200 & ~n1484;
  assign n1522 = ~n1420 & ~n1432;
  assign n1523 = ~n106 & n1522;
  assign n1524 = n318 & ~n1523;
  assign n1525 = ~n1521 & ~n1524;
  assign n1526 = ~n1520 & n1525;
  assign n1527 = n611 & ~n999;
  assign n1528 = n201 & ~n1527;
  assign n1529 = n200 & ~n624;
  assign n1530 = ~n559 & ~n1529;
  assign n1531 = ~n1528 & n1530;
  assign n1532 = ~i_12_ & n213;
  assign n1533 = ~n1135 & ~n1532;
  assign n1534 = n318 & ~n1533;
  assign n1535 = n201 & n411;
  assign n1536 = ~n69 & n1002;
  assign n1537 = ~n244 & ~n1416;
  assign n1538 = ~n1536 & n1537;
  assign n1539 = n318 & ~n1538;
  assign n1540 = ~n1535 & ~n1539;
  assign n1541 = ~n1534 & n1540;
  assign n1542 = ~n435 & ~n1153;
  assign n1543 = n116 & n1404;
  assign n1544 = n1542 & ~n1543;
  assign n1545 = n318 & ~n1544;
  assign n1546 = n106 & n201;
  assign n1547 = ~n347 & ~n1546;
  assign n1548 = ~n1545 & n1547;
  assign n1549 = n1541 & n1548;
  assign n1550 = n1531 & n1549;
  assign n1551 = n1526 & n1550;
  assign n1552 = ~n274 & ~n1430;
  assign n1553 = ~n296 & n1552;
  assign n1554 = ~n595 & ~n1553;
  assign n1555 = ~n787 & ~n1418;
  assign n1556 = ~n885 & ~n1555;
  assign n1557 = n203 & n1172;
  assign n1558 = ~n1536 & n1542;
  assign n1559 = ~n267 & ~n285;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = n102 & n1404;
  assign n1562 = n201 & n1561;
  assign n1563 = ~n1560 & ~n1562;
  assign n1564 = ~n1557 & n1563;
  assign n1565 = ~i_14_ & n464;
  assign n1566 = i_12_ & n1565;
  assign n1567 = ~n326 & ~n1566;
  assign n1568 = n1376 & n1567;
  assign n1569 = n226 & ~n1568;
  assign n1570 = n328 & n651;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = n1564 & n1571;
  assign n1573 = ~n953 & n1572;
  assign n1574 = ~n1556 & n1573;
  assign n1575 = ~n1554 & n1574;
  assign n1576 = n1551 & n1575;
  assign n1577 = n198 & ~n1496;
  assign n1578 = n624 & ~n1561;
  assign n1579 = n345 & ~n1578;
  assign n1580 = ~n887 & ~n970;
  assign n1581 = ~n1579 & n1580;
  assign n1582 = ~n1577 & n1581;
  assign n1583 = n105 & n121;
  assign n1584 = ~n952 & n1583;
  assign n1585 = n1582 & ~n1584;
  assign n1586 = i_8_ & n1536;
  assign n1587 = ~n119 & ~n1586;
  assign n1588 = ~n249 & n1587;
  assign n1589 = n221 & ~n1588;
  assign n1590 = n417 & n1404;
  assign n1591 = ~n615 & ~n1590;
  assign n1592 = n400 & ~n1591;
  assign n1593 = ~n552 & ~n1533;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1589 & n1594;
  assign n1596 = ~n285 & ~n318;
  assign n1597 = ~n69 & n1027;
  assign n1598 = ~n1596 & n1597;
  assign n1599 = n121 & n1404;
  assign n1600 = ~n269 & n1599;
  assign n1601 = ~n1598 & ~n1600;
  assign n1602 = ~n103 & ~n786;
  assign n1603 = ~n1543 & n1602;
  assign n1604 = n198 & ~n1603;
  assign n1605 = n1601 & ~n1604;
  assign n1606 = ~n760 & ~n901;
  assign n1607 = n374 & ~n1376;
  assign n1608 = n197 & n613;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = ~n924 & n1609;
  assign n1611 = ~n1606 & n1610;
  assign n1612 = n1605 & n1611;
  assign n1613 = n1595 & n1612;
  assign n1614 = ~n95 & ~n266;
  assign n1615 = ~n255 & n594;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = n1613 & ~n1616;
  assign n1618 = n1585 & n1617;
  assign n1619 = n495 & n1618;
  assign n1620 = n1576 & n1619;
  assign n1621 = n344 & n1397;
  assign n1622 = n1542 & ~n1597;
  assign n1623 = ~n451 & ~n1622;
  assign n1624 = n209 & n326;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = ~n1621 & n1625;
  assign n1627 = ~n1186 & n1542;
  assign n1628 = n1503 & n1627;
  assign n1629 = n256 & ~n1628;
  assign n1630 = ~n1175 & n1187;
  assign n1631 = n772 & n1630;
  assign n1632 = n285 & ~n1631;
  assign n1633 = ~n1629 & ~n1632;
  assign n1634 = n919 & ~n1536;
  assign n1635 = n238 & ~n1634;
  assign n1636 = n1633 & ~n1635;
  assign n1637 = n1626 & n1636;
  assign n1638 = ~n197 & n898;
  assign n1639 = ~n345 & n1638;
  assign n1640 = ~n1493 & ~n1639;
  assign n1641 = n623 & ~n1135;
  assign n1642 = n261 & ~n1641;
  assign n1643 = ~n1640 & ~n1642;
  assign n1644 = n558 & n1643;
  assign n1645 = n517 & n1644;
  assign n1646 = n1637 & n1645;
  assign n1647 = n105 & n443;
  assign n1648 = ~n681 & ~n1647;
  assign n1649 = ~n936 & ~n1648;
  assign n1650 = ~n395 & ~n1397;
  assign n1651 = ~n1151 & n1650;
  assign n1652 = n816 & n1651;
  assign n1653 = n232 & ~n1652;
  assign n1654 = n425 & ~n919;
  assign n1655 = n920 & n1049;
  assign n1656 = n237 & ~n1655;
  assign n1657 = n123 & ~n288;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1654 & n1658;
  assign n1660 = ~n1653 & n1659;
  assign n1661 = ~n1649 & n1660;
  assign n1662 = n255 & ~n1567;
  assign n1663 = n623 & ~n786;
  assign n1664 = n238 & ~n1663;
  assign n1665 = ~n1662 & ~n1664;
  assign n1666 = ~n612 & ~n735;
  assign n1667 = n1665 & ~n1666;
  assign n1668 = n1262 & n1667;
  assign n1669 = n878 & n1668;
  assign n1670 = n1661 & n1669;
  assign n1671 = n1646 & n1670;
  assign n1672 = n1620 & n1671;
  assign n1673 = n91 & n417;
  assign n1674 = ~i_14_ & n1673;
  assign n1675 = ~n1151 & ~n1674;
  assign n1676 = n200 & ~n1675;
  assign n1677 = n95 & n371;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1543 & ~n1590;
  assign n1680 = n287 & ~n1679;
  assign n1681 = n1678 & ~n1680;
  assign n1682 = ~n576 & ~n1187;
  assign n1683 = n327 & n655;
  assign n1684 = ~i_9_ & n1683;
  assign n1685 = ~n66 & n1684;
  assign n1686 = ~n805 & ~n1647;
  assign n1687 = n198 & ~n1686;
  assign n1688 = ~n1685 & ~n1687;
  assign n1689 = ~n1682 & n1688;
  assign n1690 = ~n91 & n805;
  assign n1691 = ~n288 & n1690;
  assign n1692 = n1689 & ~n1691;
  assign n1693 = n1681 & n1692;
  assign n1694 = n105 & n429;
  assign n1695 = ~n756 & n1694;
  assign n1696 = ~n371 & ~n519;
  assign n1697 = ~n198 & n1696;
  assign n1698 = n1599 & ~n1697;
  assign n1699 = ~n1405 & ~n1583;
  assign n1700 = n218 & ~n1699;
  assign n1701 = n102 & n105;
  assign n1702 = ~n1694 & ~n1701;
  assign n1703 = n226 & ~n1702;
  assign n1704 = ~n1700 & ~n1703;
  assign n1705 = ~n1698 & n1704;
  assign n1706 = n1555 & ~n1561;
  assign n1707 = ~n1690 & n1706;
  assign n1708 = ~n766 & ~n1707;
  assign n1709 = n1705 & ~n1708;
  assign n1710 = ~n1695 & n1709;
  assign n1711 = n1693 & n1710;
  assign n1712 = ~n1674 & ~n1694;
  assign n1713 = n256 & ~n1712;
  assign n1714 = n295 & n1647;
  assign n1715 = n429 & n1404;
  assign n1716 = n256 & n1715;
  assign n1717 = ~n1714 & ~n1716;
  assign n1718 = n295 & n1583;
  assign n1719 = n1717 & ~n1718;
  assign n1720 = ~n1713 & n1719;
  assign n1721 = ~n256 & ~n344;
  assign n1722 = ~n197 & n1015;
  assign n1723 = n1446 & n1722;
  assign n1724 = n1721 & n1723;
  assign n1725 = n1701 & ~n1724;
  assign n1726 = ~n1505 & ~n1674;
  assign n1727 = i_8_ & ~n1726;
  assign n1728 = ~n1561 & ~n1727;
  assign n1729 = n519 & ~n1728;
  assign n1730 = n287 & n1715;
  assign n1731 = n497 & n1701;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1729 & n1732;
  assign n1734 = n1679 & ~n1690;
  assign n1735 = n497 & ~n1734;
  assign n1736 = n287 & n1405;
  assign n1737 = n287 & n1507;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = n1733 & n1739;
  assign n1741 = ~n1725 & n1740;
  assign n1742 = n1720 & n1741;
  assign n1743 = n1711 & n1742;
  assign n1744 = ~n587 & n1647;
  assign n1745 = ~n722 & n1505;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = n371 & n1565;
  assign n1748 = n67 & n1683;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n1746 & n1749;
  assign n1751 = n198 & n1583;
  assign n1752 = ~n1543 & ~n1674;
  assign n1753 = ~n1599 & n1752;
  assign n1754 = n261 & ~n1753;
  assign n1755 = ~n1751 & ~n1754;
  assign n1756 = n255 & ~n1223;
  assign n1757 = n239 & n417;
  assign n1758 = ~n798 & ~n1757;
  assign n1759 = ~n1599 & n1758;
  assign n1760 = n221 & ~n1759;
  assign n1761 = ~n1756 & ~n1760;
  assign n1762 = ~n198 & ~n205;
  assign n1763 = ~n255 & n1762;
  assign n1764 = n1175 & ~n1763;
  assign n1765 = n1761 & ~n1764;
  assign n1766 = n1755 & n1765;
  assign n1767 = n1750 & n1766;
  assign n1768 = n256 & n1154;
  assign n1769 = n318 & n1397;
  assign n1770 = n237 & n1135;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = n232 & n1694;
  assign n1773 = n267 & n1543;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = n1771 & n1774;
  assign n1776 = n91 & n429;
  assign n1777 = n99 & n105;
  assign n1778 = ~n1432 & ~n1777;
  assign n1779 = ~n1430 & n1778;
  assign n1780 = ~n1776 & n1779;
  assign n1781 = n295 & ~n1780;
  assign n1782 = ~n1186 & ~n1583;
  assign n1783 = n205 & ~n1782;
  assign n1784 = ~n1781 & ~n1783;
  assign n1785 = n1775 & n1784;
  assign n1786 = ~n1768 & n1785;
  assign n1787 = n1767 & n1786;
  assign n1788 = n1743 & n1787;
  assign n1789 = n105 & n464;
  assign n1790 = ~n742 & n1789;
  assign n1791 = ~n1380 & n1583;
  assign n1792 = n284 & n1175;
  assign n1793 = ~n1674 & ~n1792;
  assign n1794 = ~n221 & n719;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1791 & ~n1795;
  assign n1797 = ~n1599 & ~n1727;
  assign n1798 = ~n805 & n1679;
  assign n1799 = i_8_ & ~n1798;
  assign n1800 = ~i_8_ & n1543;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = n1797 & n1801;
  assign n1803 = n344 & ~n1802;
  assign n1804 = n443 & n1404;
  assign n1805 = n497 & n1715;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = n577 & ~n1806;
  assign n1808 = ~n1803 & ~n1807;
  assign n1809 = ~n344 & n372;
  assign n1810 = n794 & ~n1809;
  assign n1811 = n1808 & ~n1810;
  assign n1812 = n1796 & n1811;
  assign n1813 = ~n106 & n1433;
  assign n1814 = ~n595 & ~n1813;
  assign n1815 = ~n255 & n738;
  assign n1816 = n1392 & ~n1815;
  assign n1817 = ~n1814 & ~n1816;
  assign n1818 = ~n671 & n1172;
  assign n1819 = n1817 & ~n1818;
  assign n1820 = n1812 & n1819;
  assign n1821 = ~n1790 & n1820;
  assign n1822 = n1788 & n1821;
  assign n1823 = n1672 & n1822;
  assign n1824 = n782 & n1823;
  assign o_9_ = ~n1519 | ~n1824;
  assign n1826 = ~n593 & n1397;
  assign n1827 = n400 & n1420;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = n123 & ~n713;
  assign n1830 = ~n117 & ~n1390;
  assign n1831 = n198 & ~n1830;
  assign n1832 = n318 & n1416;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1546 & n1833;
  assign n1835 = ~n1829 & n1834;
  assign n1836 = n1828 & n1835;
  assign n1837 = ~n885 & ~n1419;
  assign n1838 = ~n1396 & ~n1430;
  assign n1839 = n256 & ~n1838;
  assign n1840 = n95 & n295;
  assign n1841 = n122 & ~n269;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1839 & n1842;
  assign n1844 = ~n1837 & n1843;
  assign n1845 = n1836 & n1844;
  assign n1846 = n1526 & n1845;
  assign n1847 = ~n1492 & n1846;
  assign n1848 = n1477 & n1847;
  assign n1849 = n1403 & n1848;
  assign n1850 = ~n759 & ~n1405;
  assign n1851 = ~n738 & ~n1850;
  assign n1852 = ~n610 & ~n1851;
  assign n1853 = n914 & n1115;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = n285 & ~n1177;
  assign n1856 = ~n1854 & ~n1855;
  assign n1857 = ~n594 & n1430;
  assign n1858 = n237 & n799;
  assign n1859 = n255 & n1172;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = n117 & n318;
  assign n1862 = n1860 & ~n1861;
  assign n1863 = ~n1857 & n1862;
  assign n1864 = ~n256 & n941;
  assign n1865 = n785 & ~n1864;
  assign n1866 = n1135 & ~n1638;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = n1863 & n1867;
  assign n1869 = ~n964 & ~n1501;
  assign n1870 = n807 & ~n976;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n766 & n1123;
  assign n1873 = n1871 & ~n1872;
  assign n1874 = n1868 & n1873;
  assign n1875 = n1856 & n1874;
  assign n1876 = n797 & ~n1060;
  assign n1877 = n95 & ~n595;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n936 & n1647;
  assign n1880 = n810 & ~n915;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n186 & n1881;
  assign n1883 = n1878 & n1882;
  assign n1884 = ~n400 & n713;
  assign n1885 = n1186 & ~n1884;
  assign n1886 = n123 & n284;
  assign n1887 = ~n925 & ~n1886;
  assign n1888 = ~n783 & ~n1397;
  assign n1889 = n400 & ~n1888;
  assign n1890 = n232 & n794;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = n1887 & n1891;
  assign n1893 = ~n1885 & n1892;
  assign n1894 = ~n939 & n1166;
  assign n1895 = ~n972 & n1153;
  assign n1896 = ~n930 & n1154;
  assign n1897 = n345 & n1162;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1895 & n1898;
  assign n1900 = ~n1894 & n1899;
  assign n1901 = n622 & ~n941;
  assign n1902 = ~n332 & n999;
  assign n1903 = ~n786 & ~n1044;
  assign n1904 = n425 & ~n1903;
  assign n1905 = n792 & ~n1353;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = ~n1902 & n1906;
  assign n1908 = ~n1901 & n1907;
  assign n1909 = ~n1584 & n1908;
  assign n1910 = n1900 & n1909;
  assign n1911 = n1893 & n1910;
  assign n1912 = n1509 & n1911;
  assign n1913 = n1883 & n1912;
  assign n1914 = n1875 & n1913;
  assign n1915 = n1849 & n1914;
  assign n1916 = n912 & n1272;
  assign n1917 = n1822 & n1916;
  assign o_10_ = ~n1915 | ~n1917;
  assign n1919 = n63 & n86;
  assign o_11_ = ~n139 | n1919;
  assign n1921 = ~n1300 & n1328;
  assign n1922 = ~n740 & ~n1921;
  assign n1923 = ~n71 & ~n1922;
  assign n1924 = ~n1274 & ~n1923;
  assign n1925 = n1849 & ~n1924;
  assign n1926 = n70 & n190;
  assign n1927 = ~i_8_ & n203;
  assign n1928 = ~n361 & ~n1927;
  assign n1929 = n1722 & n1928;
  assign n1930 = n1926 & ~n1929;
  assign n1931 = n69 & n1429;
  assign n1932 = n579 & n1928;
  assign n1933 = n1931 & ~n1932;
  assign n1934 = ~n1930 & ~n1933;
  assign n1935 = n70 & n100;
  assign n1936 = n198 & n1935;
  assign n1937 = ~n256 & ~n371;
  assign n1938 = ~i_14_ & n190;
  assign n1939 = ~n69 & n1938;
  assign n1940 = n256 & n1939;
  assign n1941 = ~n69 & n94;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = ~n1937 & ~n1942;
  assign n1944 = ~n1936 & ~n1943;
  assign n1945 = n212 & n1062;
  assign n1946 = n99 & n1062;
  assign n1947 = ~i_15_ & n1946;
  assign n1948 = ~n1945 & ~n1947;
  assign n1949 = n200 & ~n1948;
  assign n1950 = n216 & n655;
  assign n1951 = i_9_ & n1950;
  assign n1952 = n201 & n1931;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = ~n1949 & n1953;
  assign n1955 = n1944 & n1954;
  assign n1956 = n1934 & n1955;
  assign n1957 = ~n104 & ~n239;
  assign n1958 = n234 & ~n1957;
  assign n1959 = ~n1931 & ~n1958;
  assign n1960 = ~n1935 & n1959;
  assign n1961 = n287 & ~n1960;
  assign n1962 = n100 & ~n1957;
  assign n1963 = n519 & n1962;
  assign n1964 = ~n69 & n1429;
  assign n1965 = ~n1938 & ~n1964;
  assign n1966 = n497 & ~n1965;
  assign n1967 = ~n1963 & ~n1966;
  assign n1968 = ~n1961 & n1967;
  assign n1969 = n300 & n1437;
  assign n1970 = ~n941 & ~n1969;
  assign n1971 = n206 & n227;
  assign n1972 = n736 & n1971;
  assign n1973 = ~n295 & n1972;
  assign n1974 = n1935 & ~n1973;
  assign n1975 = ~n1970 & ~n1974;
  assign n1976 = n1968 & n1975;
  assign n1977 = n1956 & n1976;
  assign n1978 = ~n1938 & ~n1941;
  assign n1979 = ~i_8_ & ~n1978;
  assign n1980 = ~n1962 & ~n1964;
  assign n1981 = n68 & ~n1957;
  assign n1982 = n1980 & ~n1981;
  assign n1983 = ~n1935 & n1982;
  assign n1984 = i_8_ & ~n1983;
  assign n1985 = n118 & ~n1957;
  assign n1986 = n1959 & ~n1985;
  assign n1987 = ~n1984 & n1986;
  assign n1988 = ~n1979 & n1987;
  assign n1989 = n344 & ~n1988;
  assign n1990 = n214 & ~n594;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = n70 & n248;
  assign n1993 = ~n1945 & ~n1992;
  assign n1994 = ~n225 & n1993;
  assign n1995 = ~n1418 & n1994;
  assign n1996 = n256 & ~n1995;
  assign n1997 = n114 & ~n1060;
  assign n1998 = ~n372 & n1073;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1996 & n1999;
  assign n2001 = ~n400 & n1277;
  assign n2002 = n1981 & ~n2001;
  assign n2003 = n123 & ~n580;
  assign n2004 = ~n296 & ~n1096;
  assign n2005 = n237 & ~n2004;
  assign n2006 = ~n284 & ~n1931;
  assign n2007 = ~n1429 & ~n1962;
  assign n2008 = ~n1958 & n2007;
  assign n2009 = ~n576 & ~n2008;
  assign n2010 = ~n2006 & n2009;
  assign n2011 = ~n2005 & ~n2010;
  assign n2012 = n131 & n371;
  assign n2013 = n256 & n1935;
  assign n2014 = ~n284 & ~n286;
  assign n2015 = ~n1978 & ~n2014;
  assign n2016 = ~n2013 & ~n2015;
  assign n2017 = ~n2012 & n2016;
  assign n2018 = n2011 & n2017;
  assign n2019 = ~n2003 & n2018;
  assign n2020 = ~n2002 & n2019;
  assign n2021 = ~n1088 & ~n1280;
  assign n2022 = n713 & n1163;
  assign n2023 = n1064 & ~n2022;
  assign n2024 = n249 & ~n738;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n2021 & n2025;
  assign n2027 = n2020 & n2026;
  assign n2028 = n2000 & n2027;
  assign n2029 = n1991 & n2028;
  assign n2030 = n1977 & n2029;
  assign n2031 = n1925 & n2030;
  assign n2032 = n1079 & ~n1273;
  assign n2033 = n248 & ~n1957;
  assign n2034 = ~n737 & n2033;
  assign n2035 = n131 & ~n269;
  assign n2036 = ~n235 & ~n1413;
  assign n2037 = ~n976 & ~n2036;
  assign n2038 = n197 & n1110;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~n1939 & n1980;
  assign n2041 = n287 & n1964;
  assign n2042 = ~n232 & ~n2041;
  assign n2043 = ~n2040 & ~n2042;
  assign n2044 = ~n117 & ~n2033;
  assign n2045 = n345 & ~n2044;
  assign n2046 = ~n2043 & ~n2045;
  assign n2047 = n2039 & n2046;
  assign n2048 = ~n2035 & n2047;
  assign n2049 = ~n2034 & n2048;
  assign n2050 = ~n2032 & n2049;
  assign n2051 = n70 & n234;
  assign n2052 = n132 & n1298;
  assign n2053 = ~n2051 & n2052;
  assign n2054 = ~n1133 & ~n2053;
  assign n2055 = ~n915 & ~n1511;
  assign n2056 = ~n713 & n1086;
  assign n2057 = ~n1353 & n1420;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n2055 & n2058;
  assign n2060 = ~n2054 & n2059;
  assign n2061 = n2050 & n2060;
  assign n2062 = ~n1283 & n1992;
  assign n2063 = n122 & ~n602;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = n189 & n1068;
  assign n2066 = n200 & n2065;
  assign n2067 = n400 & ~n1980;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~n2033 & n2040;
  assign n2070 = n295 & ~n2069;
  assign n2071 = ~n1962 & ~n1981;
  assign n2072 = n1959 & n2071;
  assign n2073 = ~n1926 & n2072;
  assign n2074 = n256 & ~n2073;
  assign n2075 = ~n2070 & ~n2074;
  assign n2076 = ~n101 & ~n242;
  assign n2077 = ~n1048 & n2076;
  assign n2078 = n425 & ~n2077;
  assign n2079 = ~n232 & ~n497;
  assign n2080 = ~n1614 & ~n2079;
  assign n2081 = ~n2078 & ~n2080;
  assign n2082 = ~n1537 & ~n2079;
  assign n2083 = ~n736 & n1397;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = n2081 & n2084;
  assign n2086 = n2075 & n2085;
  assign n2087 = n2068 & n2086;
  assign n2088 = n1095 & n2087;
  assign n2089 = n2064 & n2088;
  assign n2090 = ~n237 & n914;
  assign n2091 = n119 & ~n2090;
  assign n2092 = ~n120 & n267;
  assign n2093 = n284 & n1985;
  assign n2094 = n361 & n1992;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n232 & ~n519;
  assign n2097 = n296 & ~n2096;
  assign n2098 = n2095 & ~n2097;
  assign n2099 = ~n2092 & n2098;
  assign n2100 = ~n2091 & n2099;
  assign n2101 = n2089 & n2100;
  assign n2102 = n2061 & n2101;
  assign n2103 = n387 & n2102;
  assign o_12_ = ~n2031 | ~n2103;
  assign n2105 = ~n71 & ~n1275;
  assign n2106 = ~n1789 & n2105;
  assign n2107 = ~n733 & n2106;
  assign n2108 = ~n1134 & n2107;
  assign n2109 = ~n1141 & n2108;
  assign n2110 = ~n131 & n2109;
  assign n2111 = ~n586 & ~n1507;
  assign n2112 = ~n219 & ~n1392;
  assign n2113 = n1080 & n2112;
  assign n2114 = n2111 & n2113;
  assign n2115 = n1513 & n2114;
  assign n2116 = ~n1086 & ~n1296;
  assign n2117 = n2115 & n2116;
  assign n2118 = ~n1048 & ~n1085;
  assign n2119 = n2117 & n2118;
  assign n2120 = n2110 & n2119;
  assign n2121 = n760 & n2120;
  assign n2122 = ~n636 & ~n1674;
  assign n2123 = ~n1025 & n2122;
  assign n2124 = ~n1931 & n2123;
  assign n2125 = ~n123 & n1376;
  assign n2126 = ~n2051 & n2125;
  assign n2127 = n2124 & n2126;
  assign n2128 = n2121 & n2127;
  assign n2129 = n295 & ~n2128;
  assign n2130 = n1043 & n2075;
  assign n2131 = n1426 & n2130;
  assign n2132 = n493 & n1160;
  assign n2133 = n2131 & n2132;
  assign n2134 = ~n1599 & ~n1941;
  assign n2135 = n295 & ~n2134;
  assign n2136 = ~n1054 & ~n2135;
  assign n2137 = ~n1009 & ~n1694;
  assign n2138 = ~n696 & ~n1926;
  assign n2139 = n2137 & n2138;
  assign n2140 = n295 & ~n2139;
  assign n2141 = ~n1301 & n1648;
  assign n2142 = ~n1992 & n2141;
  assign n2143 = ~i_8_ & ~n1992;
  assign n2144 = n255 & ~n2143;
  assign n2145 = ~n2142 & n2144;
  assign n2146 = ~n2140 & ~n2145;
  assign n2147 = ~n625 & ~n1107;
  assign n2148 = ~n1701 & n2147;
  assign n2149 = n256 & ~n2148;
  assign n2150 = n2146 & ~n2149;
  assign n2151 = n2136 & n2150;
  assign n2152 = n304 & n2151;
  assign n2153 = n1720 & n2152;
  assign n2154 = n2133 & n2153;
  assign n2155 = ~n2129 & n2154;
  assign n2156 = ~n249 & n1652;
  assign n2157 = ~n2033 & n2156;
  assign n2158 = n1567 & n2157;
  assign n2159 = ~n1543 & ~n1985;
  assign n2160 = n612 & n2159;
  assign n2161 = n1591 & ~n1964;
  assign n2162 = ~n613 & ~n1599;
  assign n2163 = ~n1020 & n2162;
  assign n2164 = n2161 & n2163;
  assign n2165 = n2160 & n2164;
  assign n2166 = ~n2051 & n2111;
  assign n2167 = ~n691 & ~n1583;
  assign n2168 = ~n94 & ~n1390;
  assign n2169 = n2167 & n2168;
  assign n2170 = n2166 & n2169;
  assign n2171 = ~n462 & n2170;
  assign n2172 = n2165 & n2171;
  assign n2173 = n2158 & n2172;
  assign n2174 = n2109 & n2173;
  assign n2175 = ~n1939 & n2174;
  assign n2176 = n256 & ~n2175;
  assign n2177 = n700 & n815;
  assign n2178 = ~n2176 & n2177;
  assign n2179 = n2155 & n2178;
  assign n2180 = ~n66 & ~n188;
  assign n2181 = n141 & n2180;
  assign n2182 = n655 & n2181;
  assign n2183 = ~n575 & ~n1505;
  assign n2184 = ~n130 & ~n1142;
  assign n2185 = n2183 & n2184;
  assign n2186 = n255 & ~n2185;
  assign n2187 = ~n2013 & ~n2186;
  assign n2188 = ~n1701 & ~n1935;
  assign n2189 = n2147 & n2188;
  assign n2190 = n295 & ~n2189;
  assign n2191 = n2187 & ~n2190;
  assign n2192 = ~n2182 & n2191;
  assign o_13_ = ~n2179 | ~n2192;
  assign n2194 = ~n123 & ~n296;
  assign n2195 = n2124 & n2194;
  assign n2196 = ~n390 & ~n1035;
  assign n2197 = n1493 & n2196;
  assign n2198 = n1555 & n2197;
  assign n2199 = ~n1107 & n2183;
  assign n2200 = n2198 & n2199;
  assign n2201 = ~n1014 & ~n1536;
  assign n2202 = n1537 & n1542;
  assign n2203 = ~n1935 & n2202;
  assign n2204 = ~n1101 & n2203;
  assign n2205 = n2201 & n2204;
  assign n2206 = n2200 & n2205;
  assign n2207 = n2120 & n2206;
  assign n2208 = n2195 & n2207;
  assign n2209 = n497 & ~n2208;
  assign n2210 = n2148 & n2157;
  assign n2211 = ~n1941 & n2210;
  assign n2212 = ~n618 & ~n1690;
  assign n2213 = ~n1002 & n2212;
  assign n2214 = n687 & n2213;
  assign n2215 = n2110 & n2113;
  assign n2216 = n2165 & n2215;
  assign n2217 = n2214 & n2216;
  assign n2218 = n2211 & n2217;
  assign n2219 = n287 & ~n2218;
  assign n2220 = ~n1804 & ~n2033;
  assign n2221 = ~n1027 & n2220;
  assign n2222 = ~i_8_ & n2221;
  assign n2223 = i_8_ & ~n1027;
  assign n2224 = ~n1938 & n2223;
  assign n2225 = ~n2222 & ~n2224;
  assign n2226 = n2142 & ~n2225;
  assign n2227 = n519 & ~n2226;
  assign n2228 = n497 & ~n763;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = n497 & ~n2134;
  assign n2231 = ~n1055 & ~n2230;
  assign n2232 = ~n696 & ~n1694;
  assign n2233 = ~n1009 & n2232;
  assign n2234 = n1376 & n2233;
  assign n2235 = ~n2051 & n2184;
  assign n2236 = n2167 & n2235;
  assign n2237 = n2234 & n2236;
  assign n2238 = n519 & ~n2237;
  assign n2239 = n1968 & ~n2238;
  assign n2240 = n1316 & n2239;
  assign n2241 = n2231 & n2240;
  assign n2242 = n635 & n2241;
  assign n2243 = n2229 & n2242;
  assign n2244 = n1740 & n2243;
  assign n2245 = ~n2219 & n2244;
  assign o_14_ = n2209 | ~n2245;
  assign n2247 = ~n1134 & n2167;
  assign n2248 = n371 & ~n2247;
  assign n2249 = ~n91 & n613;
  assign n2250 = ~n131 & ~n2249;
  assign n2251 = ~n1019 & n2250;
  assign n2252 = ~n797 & n2134;
  assign n2253 = n2167 & n2252;
  assign n2254 = n2251 & n2253;
  assign n2255 = n218 & ~n2254;
  assign n2256 = ~n2248 & ~n2255;
  assign n2257 = ~n1014 & n2167;
  assign n2258 = ~n1101 & ~n1599;
  assign n2259 = n93 & ~n409;
  assign n2260 = ~n1134 & ~n2259;
  assign n2261 = n2258 & n2260;
  assign n2262 = n2257 & n2261;
  assign n2263 = n268 & ~n2262;
  assign n2264 = n2256 & ~n2263;
  assign n2265 = ~n650 & n2106;
  assign n2266 = ~n1405 & n2112;
  assign n2267 = n1080 & n1376;
  assign n2268 = n2266 & n2267;
  assign n2269 = n2265 & n2268;
  assign n2270 = n328 & ~n2269;
  assign n2271 = ~n94 & n2163;
  assign n2272 = i_8_ & ~n2271;
  assign n2273 = n2269 & ~n2272;
  assign n2274 = n370 & ~n2273;
  assign n2275 = ~n2270 & ~n2274;
  assign o_15_ = ~n2264 | ~n2275;
  assign n2277 = ~n1001 & n2160;
  assign n2278 = n2185 & n2277;
  assign n2279 = n267 & ~n2278;
  assign n2280 = ~n91 & n651;
  assign n2281 = ~n810 & ~n1029;
  assign n2282 = n2266 & n2281;
  assign n2283 = ~n2280 & n2282;
  assign n2284 = n374 & ~n2283;
  assign n2285 = ~n2279 & ~n2284;
  assign n2286 = n267 & ~n2262;
  assign n2287 = ~n617 & ~n1507;
  assign n2288 = ~n1002 & n2287;
  assign n2289 = n233 & n239;
  assign n2290 = ~n1141 & ~n2051;
  assign n2291 = ~n2289 & n2290;
  assign n2292 = n1417 & n2291;
  assign n2293 = n2288 & n2292;
  assign n2294 = n267 & ~n2293;
  assign n2295 = ~n1073 & n2107;
  assign n2296 = n374 & ~n2295;
  assign n2297 = ~n2294 & ~n2296;
  assign n2298 = ~n2286 & n2297;
  assign o_16_ = ~n2285 | ~n2298;
  assign n2300 = i_8_ & n1926;
  assign n2301 = n2110 & ~n2300;
  assign n2302 = n2142 & n2236;
  assign n2303 = n2301 & n2302;
  assign n2304 = n1988 & n2303;
  assign n2305 = n1802 & n2304;
  assign n2306 = ~n1029 & n1513;
  assign n2307 = n2211 & n2306;
  assign n2308 = ~n1040 & n2307;
  assign n2309 = i_8_ & ~n2308;
  assign n2310 = n2305 & ~n2309;
  assign n2311 = n344 & ~n2310;
  assign n2312 = ~n1027 & n2157;
  assign n2313 = n400 & ~n2312;
  assign n2314 = n1555 & ~n1939;
  assign n2315 = n2197 & n2314;
  assign n2316 = n345 & ~n2315;
  assign n2317 = ~n1367 & ~n2316;
  assign n2318 = ~n2313 & n2317;
  assign n2319 = n2198 & n2233;
  assign n2320 = n400 & ~n2319;
  assign n2321 = ~n1579 & ~n2320;
  assign n2322 = n345 & ~n2233;
  assign n2323 = ~n1561 & ~n1962;
  assign n2324 = n400 & ~n2323;
  assign n2325 = ~n2322 & ~n2324;
  assign n2326 = ~n1345 & n2325;
  assign n2327 = n2321 & n2326;
  assign n2328 = n1376 & n2212;
  assign n2329 = n2161 & n2328;
  assign n2330 = n2188 & n2199;
  assign n2331 = n2329 & n2330;
  assign n2332 = n2123 & n2331;
  assign n2333 = n2115 & n2332;
  assign n2334 = n400 & ~n2333;
  assign n2335 = n754 & ~n2334;
  assign n2336 = n2327 & n2335;
  assign n2337 = n2318 & n2336;
  assign o_17_ = n2311 | ~n2337;
  assign n2339 = n1291 & n1493;
  assign n2340 = ~n1154 & n1537;
  assign n2341 = n1686 & n2340;
  assign n2342 = ~n617 & n2118;
  assign n2343 = n2341 & n2342;
  assign n2344 = n2339 & n2343;
  assign n2345 = ~n1543 & n2116;
  assign n2346 = ~n1153 & n2345;
  assign n2347 = n2194 & n2346;
  assign n2348 = n611 & n2347;
  assign n2349 = n1602 & ~n1947;
  assign n2350 = n1293 & n1496;
  assign n2351 = n2349 & n2350;
  assign n2352 = n2348 & n2351;
  assign n2353 = ~i_12_ & n1019;
  assign n2354 = ~n1083 & ~n2353;
  assign n2355 = n2162 & n2354;
  assign n2356 = ~n691 & n1407;
  assign n2357 = n2355 & n2356;
  assign n2358 = n2148 & n2357;
  assign n2359 = n2352 & n2358;
  assign n2360 = n2344 & n2359;
  assign n2361 = n2215 & n2360;
  assign n2362 = ~n1992 & n2361;
  assign n2363 = n198 & ~n2362;
  assign n2364 = ~n1025 & ~n1931;
  assign n2365 = n2194 & n2364;
  assign n2366 = ~n613 & ~n1941;
  assign n2367 = ~n1757 & n2137;
  assign n2368 = n2366 & n2367;
  assign n2369 = n2365 & n2368;
  assign n2370 = ~n420 & ~n610;
  assign n2371 = n2257 & n2370;
  assign n2372 = n1376 & ~n1926;
  assign n2373 = n1327 & n2372;
  assign n2374 = n2371 & n2373;
  assign n2375 = n2369 & n2374;
  assign n2376 = n2120 & n2375;
  assign n2377 = ~n767 & ~n1690;
  assign n2378 = ~n1420 & ~n1945;
  assign n2379 = ~n1935 & n2378;
  assign n2380 = n1555 & ~n2065;
  assign n2381 = ~n119 & n2380;
  assign n2382 = n697 & n2381;
  assign n2383 = n2379 & n2382;
  assign n2384 = n2377 & n2383;
  assign n2385 = n2376 & n2384;
  assign n2386 = n261 & ~n2385;
  assign n2387 = ~n2363 & ~n2386;
  assign n2388 = n1493 & n2143;
  assign n2389 = n1648 & n2220;
  assign n2390 = n760 & n2196;
  assign n2391 = n2389 & n2390;
  assign n2392 = n2388 & n2391;
  assign n2393 = i_8_ & ~n681;
  assign n2394 = n378 & n2393;
  assign n2395 = n91 & n248;
  assign n2396 = ~n1064 & ~n2395;
  assign n2397 = ~n1804 & n2396;
  assign n2398 = ~n1694 & n2138;
  assign n2399 = n2314 & n2398;
  assign n2400 = n2397 & n2399;
  assign n2401 = n2394 & n2400;
  assign n2402 = ~n2392 & ~n2401;
  assign n2403 = ~n395 & ~n444;
  assign n2404 = ~n2402 & n2403;
  assign n2405 = n197 & ~n2404;
  assign n2406 = n197 & ~n2185;
  assign n2407 = ~n1936 & ~n2406;
  assign n2408 = ~n1532 & ~n1757;
  assign n2409 = n2378 & n2408;
  assign n2410 = n1350 & n2124;
  assign n2411 = n2409 & n2410;
  assign n2412 = n198 & ~n2411;
  assign n2413 = n623 & n2323;
  assign n2414 = n261 & ~n2413;
  assign n2415 = ~n1052 & ~n2414;
  assign n2416 = ~n2412 & n2415;
  assign n2417 = n517 & n2416;
  assign n2418 = n2407 & n2417;
  assign n2419 = ~n2405 & n2418;
  assign n2420 = n261 & ~n2148;
  assign n2421 = n197 & n2051;
  assign n2422 = n198 & n1166;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~n2420 & n2423;
  assign n2425 = ~n859 & n2424;
  assign n2426 = ~n1179 & n2425;
  assign n2427 = n282 & n2426;
  assign n2428 = n1755 & n2427;
  assign n2429 = n1436 & n2428;
  assign n2430 = n2419 & n2429;
  assign o_18_ = ~n2387 | ~n2430;
  assign n2432 = n74 & n77;
  assign n2433 = i_3_ & i_5_;
  assign n2434 = ~i_4_ & n2433;
  assign o_19_ = n2432 & n2434;
  assign n2436 = i_3_ & i_4_;
  assign n2437 = ~i_5_ & n2436;
  assign o_20_ = n2432 & n2437;
  assign n2439 = ~n172 & ~n176;
  assign n2440 = n130 & ~n2439;
  assign n2441 = n87 & n217;
  assign n2442 = ~n167 & n2441;
  assign o_21_ = n2440 | n2442;
  assign n2444 = n87 & n165;
  assign n2445 = n216 & n2444;
  assign n2446 = ~n167 & n2445;
  assign n2447 = ~n136 & ~n143;
  assign n2448 = n130 & ~n2447;
  assign o_22_ = n2446 | n2448;
  assign n2450 = n171 & n183;
  assign n2451 = ~n129 & ~n146;
  assign n2452 = n156 & ~n2442;
  assign n2453 = n2451 & n2452;
  assign n2454 = n65 & n150;
  assign n2455 = n87 & n2454;
  assign n2456 = n89 & n2444;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2445 & n2457;
  assign n2459 = ~n167 & ~n2458;
  assign n2460 = ~n96 & ~n2459;
  assign n2461 = n2453 & n2460;
  assign o_23_ = ~n2450 | ~n2461;
  assign n2463 = n87 & n2436;
  assign o_24_ = n141 & n2463;
  assign o_25_ = n112 & n2463;
  assign n2466 = n134 & n154;
  assign n2467 = ~n88 & ~n161;
  assign n2468 = n89 & ~n2467;
  assign n2469 = n2457 & ~n2468;
  assign n2470 = ~n2441 & ~n2445;
  assign n2471 = n2469 & n2470;
  assign n2472 = n117 & ~n2471;
  assign n2473 = ~n2466 & ~n2472;
  assign n2474 = n141 & n154;
  assign n2475 = n119 & ~n2471;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n123 & ~n2471;
  assign n2478 = n87 & ~n134;
  assign n2479 = n2437 & n2478;
  assign n2480 = ~n2477 & ~n2479;
  assign n2481 = n2476 & n2480;
  assign o_26_ = ~n2473 | ~n2481;
  assign n2483 = n149 & n154;
  assign n2484 = n114 & ~n2471;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = i_4_ & n2433;
  assign n2487 = n2478 & n2486;
  assign n2488 = n2485 & ~n2487;
  assign n2489 = n112 & n154;
  assign n2490 = n122 & ~n2471;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = n95 & ~n2471;
  assign n2493 = n2491 & ~n2492;
  assign o_27_ = ~n2488 | ~n2493;
  assign n2495 = n103 & ~n2469;
  assign n2496 = n2473 & ~n2495;
  assign o_28_ = ~n2491 | ~n2496;
  assign n2498 = n106 & ~n2469;
  assign n2499 = ~n2477 & ~n2498;
  assign o_29_ = n2492 | ~n2499;
  assign n2501 = n1299 & n2108;
  assign n2502 = n1303 & n2501;
  assign n2503 = n361 & ~n2502;
  assign n2504 = ~n1142 & n2183;
  assign n2505 = n2398 & n2504;
  assign n2506 = n2189 & n2505;
  assign n2507 = ~n91 & n615;
  assign n2508 = ~n1096 & ~n1945;
  assign n2509 = ~n791 & ~n1590;
  assign n2510 = n2508 & n2509;
  assign n2511 = ~n2507 & n2510;
  assign n2512 = n2123 & n2511;
  assign n2513 = n2166 & n2512;
  assign n2514 = n2506 & n2513;
  assign n2515 = ~n131 & n2514;
  assign n2516 = n205 & ~n2515;
  assign n2517 = n2141 & n2232;
  assign n2518 = ~n131 & n2167;
  assign n2519 = n1542 & n2185;
  assign n2520 = n2518 & n2519;
  assign n2521 = n2373 & n2520;
  assign n2522 = n2517 & n2521;
  assign n2523 = n2124 & n2522;
  assign n2524 = n226 & ~n2523;
  assign n2525 = ~n2516 & ~n2524;
  assign n2526 = ~n2503 & n2525;
  assign n2527 = n368 & n880;
  assign n2528 = n1499 & n2527;
  assign n2529 = ~i_12_ & n444;
  assign n2530 = ~n1064 & ~n2529;
  assign n2531 = n2156 & n2530;
  assign n2532 = n205 & ~n2531;
  assign n2533 = ~n430 & n2339;
  assign n2534 = n226 & ~n2533;
  assign n2535 = ~n226 & ~n1399;
  assign n2536 = ~n795 & ~n1063;
  assign n2537 = ~n2395 & n2536;
  assign n2538 = ~n2535 & ~n2537;
  assign n2539 = n226 & n1397;
  assign n2540 = ~n260 & ~n2539;
  assign n2541 = n283 & n361;
  assign n2542 = ~n555 & ~n2541;
  assign n2543 = n2540 & n2542;
  assign n2544 = ~n2538 & n2543;
  assign n2545 = ~n2534 & n2544;
  assign n2546 = ~n2532 & n2545;
  assign n2547 = ~n1141 & ~n1931;
  assign n2548 = n205 & ~n2547;
  assign n2549 = ~n1141 & n2166;
  assign n2550 = n226 & ~n2549;
  assign n2551 = ~n2548 & ~n2550;
  assign n2552 = n2191 & n2551;
  assign n2553 = n1266 & n2552;
  assign n2554 = n361 & ~n2141;
  assign n2555 = i_8_ & n2554;
  assign n2556 = n130 & n205;
  assign n2557 = n226 & ~n2147;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = n226 & ~n2188;
  assign n2560 = ~n2094 & ~n2559;
  assign n2561 = n2558 & n2560;
  assign n2562 = ~n2555 & n2561;
  assign n2563 = i_8_ & i_9_;
  assign n2564 = i_11_ & n2563;
  assign n2565 = n1069 & ~n2564;
  assign n2566 = ~n247 & n2565;
  assign n2567 = n205 & ~n2314;
  assign n2568 = ~n395 & ~n1027;
  assign n2569 = n226 & ~n2568;
  assign n2570 = n205 & ~n2167;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = ~n2567 & n2571;
  assign n2573 = ~n2566 & n2572;
  assign n2574 = n2562 & n2573;
  assign n2575 = n2553 & n2574;
  assign n2576 = n2546 & n2575;
  assign n2577 = n2528 & n2576;
  assign n2578 = n2526 & n2577;
  assign o_34_ = ~n2179 | ~n2578;
  assign n2580 = n101 & ~n2469;
  assign n2581 = n2476 & n2485;
  assign n2582 = ~n2580 & n2581;
  assign o_30_ = o_34_ | ~n2582;
  assign n2584 = i_7_ & ~n2467;
  assign n2585 = n149 & n2463;
  assign n2586 = n134 & n2486;
  assign n2587 = n87 & n2586;
  assign n2588 = ~n2585 & ~n2587;
  assign o_31_ = n2584 | ~n2588;
  assign n2590 = ~o_34_ & ~n2587;
  assign n2591 = n108 & n167;
  assign n2592 = n2456 & ~n2591;
  assign n2593 = ~n2446 & n2450;
  assign n2594 = ~n2592 & n2593;
  assign n2595 = ~n163 & n2594;
  assign o_32_ = ~n2590 | ~n2595;
  assign n2597 = n2455 & ~n2591;
  assign n2598 = n110 & ~n2597;
  assign o_33_ = ~n2453 | ~n2598;
  assign n2600 = ~n240 & ~n1939;
  assign n2601 = ~n622 & ~n1715;
  assign n2602 = ~n958 & n2601;
  assign n2603 = n108 & n2602;
  assign n2604 = n1291 & n2603;
  assign n2605 = n2600 & n2604;
  assign n2606 = ~n415 & n2605;
  assign n2607 = n201 & ~n2606;
  assign n2608 = ~n122 & ~n1082;
  assign n2609 = n834 & n2608;
  assign n2610 = n1614 & ~n1931;
  assign n2611 = n2609 & n2610;
  assign n2612 = n2251 & n2611;
  assign n2613 = n205 & ~n2612;
  assign n2614 = ~n2607 & ~n2613;
  assign n2615 = n1614 & n2355;
  assign n2616 = ~n458 & n2615;
  assign n2617 = ~n552 & ~n2616;
  assign n2618 = n2399 & n2518;
  assign n2619 = n198 & ~n2618;
  assign n2620 = ~n2617 & ~n2619;
  assign n2621 = n2614 & n2620;
  assign n2622 = ~n1035 & n2138;
  assign n2623 = n256 & ~n2622;
  assign n2624 = ~n693 & ~n2623;
  assign n2625 = ~n2570 & n2624;
  assign n2626 = n1944 & n2625;
  assign n2627 = n256 & n1134;
  assign n2628 = ~n1716 & ~n2627;
  assign n2629 = n205 & ~n2399;
  assign n2630 = n2017 & ~n2629;
  assign n2631 = n2628 & n2630;
  assign n2632 = n2626 & n2631;
  assign n2633 = ~n284 & n713;
  assign n2634 = ~n2518 & ~n2633;
  assign n2635 = n345 & ~n2198;
  assign n2636 = ~n256 & n2014;
  assign n2637 = ~n371 & n2636;
  assign n2638 = ~n2163 & ~n2637;
  assign n2639 = ~n2635 & ~n2638;
  assign n2640 = ~n2634 & n2639;
  assign n2641 = n2632 & n2640;
  assign n2642 = n2621 & n2641;
  assign n2643 = ~n413 & ~n1946;
  assign n2644 = ~n103 & n2189;
  assign n2645 = n1663 & n2644;
  assign n2646 = n2643 & n2645;
  assign n2647 = n361 & ~n2646;
  assign n2648 = ~n491 & ~n515;
  assign n2649 = ~n1041 & n2648;
  assign n2650 = ~n2647 & n2649;
  assign n2651 = i_8_ & ~n2650;
  assign n2652 = ~n1040 & n2323;
  assign n2653 = n2188 & n2652;
  assign n2654 = n626 & n2653;
  assign n2655 = n284 & ~n2654;
  assign n2656 = ~n2651 & ~n2655;
  assign n2657 = ~n256 & ~n286;
  assign n2658 = n552 & n2657;
  assign n2659 = ~n2148 & ~n2658;
  assign n2660 = i_8_ & n656;
  assign n2661 = ~n149 & n2660;
  assign n2662 = n99 & n2661;
  assign n2663 = ~n2659 & ~n2662;
  assign n2664 = n198 & ~n2349;
  assign n2665 = n1962 & ~n2657;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = ~n628 & n2666;
  assign n2668 = n2663 & n2667;
  assign n2669 = ~n713 & n1561;
  assign n2670 = ~n1040 & ~n1935;
  assign n2671 = ~n913 & ~n2670;
  assign n2672 = ~n2669 & ~n2671;
  assign n2673 = ~n106 & ~n242;
  assign n2674 = n1293 & n2673;
  assign n2675 = ~n1762 & ~n2674;
  assign n2676 = n256 & ~n623;
  assign n2677 = n284 & n1107;
  assign n2678 = n99 & n409;
  assign n2679 = ~n415 & ~n2678;
  assign n2680 = n425 & ~n2679;
  assign n2681 = ~n2677 & ~n2680;
  assign n2682 = ~n2676 & n2681;
  assign n2683 = ~n2675 & n2682;
  assign n2684 = n2672 & n2683;
  assign n2685 = n1582 & n2684;
  assign n2686 = n2668 & n2685;
  assign n2687 = n2656 & n2686;
  assign n2688 = n201 & ~n2139;
  assign n2689 = n256 & ~n2137;
  assign n2690 = ~n631 & ~n2689;
  assign n2691 = n287 & n1035;
  assign n2692 = ~n390 & ~n1028;
  assign n2693 = n205 & ~n2692;
  assign n2694 = ~n478 & ~n2693;
  assign n2695 = ~n2691 & n2694;
  assign n2696 = n2690 & n2695;
  assign n2697 = ~n2688 & n2696;
  assign n2698 = n284 & ~n2198;
  assign n2699 = ~n1730 & n2233;
  assign n2700 = ~n288 & ~n2699;
  assign n2701 = ~n2698 & ~n2700;
  assign n2702 = ~n1494 & n2701;
  assign n2703 = n2697 & n2702;
  assign n2704 = ~n256 & n913;
  assign n2705 = n1931 & ~n2704;
  assign n2706 = n419 & ~n1762;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = n201 & n1945;
  assign n2709 = ~n207 & ~n1552;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2707 & n2710;
  assign n2712 = ~n1034 & n2161;
  assign n2713 = n345 & ~n2712;
  assign n2714 = ~n284 & ~n2661;
  assign n2715 = n211 & ~n2714;
  assign n2716 = ~n2123 & ~n2657;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = ~n2713 & n2717;
  assign n2719 = n2711 & n2718;
  assign n2720 = n205 & ~n2512;
  assign n2721 = n441 & n2122;
  assign n2722 = ~n104 & ~n409;
  assign n2723 = n417 & n2722;
  assign n2724 = n1533 & ~n2723;
  assign n2725 = n2721 & n2724;
  assign n2726 = n201 & ~n2725;
  assign n2727 = ~n2720 & ~n2726;
  assign n2728 = n2719 & n2727;
  assign n2729 = ~n713 & ~n2161;
  assign n2730 = ~n1098 & ~n1176;
  assign n2731 = n441 & n2508;
  assign n2732 = n2730 & n2731;
  assign n2733 = n425 & ~n2732;
  assign n2734 = ~n2729 & ~n2733;
  assign n2735 = ~n2412 & n2734;
  assign n2736 = n2728 & n2735;
  assign n2737 = n2703 & n2736;
  assign n2738 = n2687 & n2737;
  assign n2739 = n2642 & n2738;
  assign n2740 = n285 & ~n2157;
  assign n2741 = ~n2094 & ~n2740;
  assign n2742 = i_8_ & ~n2741;
  assign n2743 = n247 & n1683;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = i_14_ & n410;
  assign n2746 = n256 & n2745;
  assign n2747 = ~n2322 & ~n2746;
  assign n2748 = ~n848 & n2747;
  assign n2749 = n1049 & n2036;
  assign n2750 = ~n722 & ~n2749;
  assign n2751 = n808 & n2166;
  assign n2752 = n209 & ~n2751;
  assign n2753 = ~n2750 & ~n2752;
  assign n2754 = n1958 & ~n2636;
  assign n2755 = n233 & n2660;
  assign n2756 = ~n288 & ~n2213;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = ~n2754 & n2757;
  assign n2759 = n2753 & n2758;
  assign n2760 = ~n288 & ~n2111;
  assign n2761 = ~n1085 & ~n1141;
  assign n2762 = n237 & ~n2761;
  assign n2763 = i_8_ & n2762;
  assign n2764 = ~n2760 & ~n2763;
  assign n2765 = n345 & ~n2288;
  assign n2766 = n237 & n1586;
  assign n2767 = n345 & n1690;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = ~n2765 & n2768;
  assign n2770 = n2764 & n2769;
  assign n2771 = n1057 & n2770;
  assign n2772 = n2759 & n2771;
  assign n2773 = n2748 & n2772;
  assign n2774 = n412 & n1155;
  assign n2775 = n1417 & n2774;
  assign n2776 = n2118 & n2775;
  assign n2777 = n297 & n2776;
  assign n2778 = n205 & ~n2777;
  assign n2779 = n502 & n2344;
  assign n2780 = n198 & ~n2779;
  assign n2781 = ~n2778 & ~n2780;
  assign n2782 = n201 & ~n2340;
  assign n2783 = n2781 & ~n2782;
  assign n2784 = n2773 & n2783;
  assign n2785 = n2744 & n2784;
  assign n2786 = ~n1063 & n2121;
  assign n2787 = n201 & ~n2786;
  assign n2788 = n345 & n1981;
  assign n2789 = ~n205 & ~n2788;
  assign n2790 = ~n1141 & n1406;
  assign n2791 = n2107 & n2790;
  assign n2792 = n2113 & n2791;
  assign n2793 = ~n2789 & ~n2792;
  assign n2794 = n505 & n2183;
  assign n2795 = n2536 & n2794;
  assign n2796 = n198 & ~n2795;
  assign n2797 = ~n2793 & ~n2796;
  assign n2798 = n561 & n2797;
  assign n2799 = ~n734 & ~n2302;
  assign n2800 = ~n1027 & n2184;
  assign n2801 = ~n1992 & n2281;
  assign n2802 = n2107 & n2801;
  assign n2803 = n2800 & n2802;
  assign n2804 = n256 & ~n2803;
  assign n2805 = ~n2799 & ~n2804;
  assign n2806 = n828 & ~n2532;
  assign n2807 = n2805 & n2806;
  assign n2808 = n2798 & n2807;
  assign n2809 = ~n2787 & n2808;
  assign n2810 = n2785 & n2809;
  assign n2811 = n2739 & n2810;
  assign n2812 = ~n798 & n2183;
  assign n2813 = ~n119 & n2812;
  assign n2814 = n2157 & n2813;
  assign n2815 = n284 & ~n2814;
  assign n2816 = n256 & ~n2158;
  assign n2817 = ~n205 & ~n1215;
  assign n2818 = n1376 & ~n2555;
  assign n2819 = ~n2280 & n2818;
  assign n2820 = ~n2817 & ~n2819;
  assign n2821 = ~n2816 & ~n2820;
  assign n2822 = ~n2815 & n2821;
  assign n2823 = ~n2277 & ~n2657;
  assign n2824 = n2370 & n2504;
  assign n2825 = ~n119 & n920;
  assign n2826 = ~n123 & n2825;
  assign n2827 = n2346 & n2826;
  assign n2828 = n2824 & n2827;
  assign n2829 = n205 & ~n2828;
  assign n2830 = ~n2823 & ~n2829;
  assign n2831 = ~n575 & n921;
  assign n2832 = n425 & ~n2831;
  assign n2833 = n2830 & ~n2832;
  assign n2834 = n436 & n2348;
  assign n2835 = n198 & ~n2834;
  assign n2836 = ~n117 & ~n420;
  assign n2837 = n1542 & n2194;
  assign n2838 = n2836 & n2837;
  assign n2839 = n201 & ~n2838;
  assign n2840 = ~n845 & ~n2839;
  assign n2841 = n69 & n116;
  assign n2842 = ~n609 & ~n1985;
  assign n2843 = n436 & n2842;
  assign n2844 = ~n2841 & n2843;
  assign n2845 = n284 & ~n2844;
  assign n2846 = n115 & n2660;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = n286 & ~n2183;
  assign n2849 = ~n1528 & ~n2848;
  assign n2850 = n2847 & n2849;
  assign n2851 = n2840 & n2850;
  assign n2852 = ~n2835 & n2851;
  assign n2853 = n2833 & n2852;
  assign n2854 = n1302 & ~n1992;
  assign n2855 = n2235 & n2854;
  assign n2856 = n1080 & n2109;
  assign n2857 = n2855 & n2856;
  assign n2858 = ~n372 & ~n2857;
  assign n2859 = n1750 & ~n2858;
  assign n2860 = n2853 & n2859;
  assign n2861 = n2822 & n2860;
  assign n2862 = n2110 & n2306;
  assign n2863 = n345 & ~n2862;
  assign n2864 = n2105 & n2267;
  assign n2865 = n371 & ~n2864;
  assign n2866 = ~n1162 & n1648;
  assign n2867 = ~n651 & n2866;
  assign n2868 = n287 & ~n2867;
  assign n2869 = ~n2865 & ~n2868;
  assign n2870 = ~n2296 & n2869;
  assign n2871 = n1171 & n2870;
  assign n2872 = n256 & n1981;
  assign n2873 = ~n1535 & ~n1736;
  assign n2874 = ~n2872 & n2873;
  assign n2875 = ~n723 & ~n2248;
  assign n2876 = ~n2556 & n2875;
  assign n2877 = n2874 & n2876;
  assign n2878 = n2871 & n2877;
  assign n2879 = ~n2863 & n2878;
  assign n2880 = n1080 & n2265;
  assign n2881 = n328 & ~n2880;
  assign n2882 = n1373 & ~n2881;
  assign n2883 = n685 & n2882;
  assign n2884 = n2879 & n2883;
  assign n2885 = n1412 & n2884;
  assign n2886 = n2861 & n2885;
  assign o_35_ = ~n2811 | ~n2886;
  assign n2888 = n1578 & ~n1947;
  assign n2889 = ~n106 & n2888;
  assign n2890 = n318 & ~n2889;
  assign n2891 = ~n413 & ~n2890;
  assign n2892 = ~n1175 & n2891;
  assign n2893 = ~n735 & ~n2892;
  assign n2894 = ~n627 & ~n1935;
  assign n2895 = ~n509 & n2894;
  assign n2896 = ~n2893 & n2895;
  assign n2897 = ~n578 & ~n2896;
  assign n2898 = ~n335 & ~n923;
  assign n2899 = ~n1731 & ~n2898;
  assign n2900 = n2325 & n2899;
  assign n2901 = ~n1664 & n2900;
  assign n2902 = ~n2420 & n2901;
  assign n2903 = n242 & n318;
  assign n2904 = ~i_8_ & n656;
  assign n2905 = n99 & n2904;
  assign n2906 = n238 & n625;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n243 & n2907;
  assign n2909 = ~n2903 & n2908;
  assign n2910 = n2902 & n2909;
  assign n2911 = ~n625 & ~n1701;
  assign n2912 = n318 & ~n2911;
  assign n2913 = ~n1175 & n1496;
  assign n2914 = n2188 & n2673;
  assign n2915 = n2913 & n2914;
  assign n2916 = n2679 & n2915;
  assign n2917 = n2349 & n2916;
  assign n2918 = n232 & ~n2917;
  assign n2919 = ~n2912 & ~n2918;
  assign n2920 = n624 & n2189;
  assign n2921 = ~n295 & ~n400;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = ~n717 & n1040;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n1107 & ~n2079;
  assign n2926 = ~n295 & ~n497;
  assign n2927 = ~n2323 & ~n2926;
  assign n2928 = ~n2925 & ~n2927;
  assign n2929 = n2924 & n2928;
  assign n2930 = ~n241 & ~n1947;
  assign n2931 = n2188 & n2930;
  assign n2932 = n107 & n2931;
  assign n2933 = n2913 & n2932;
  assign n2934 = n226 & ~n2933;
  assign n2935 = n451 & n735;
  assign n2936 = n1007 & ~n2935;
  assign n2937 = n2415 & ~n2936;
  assign n2938 = ~n2934 & n2937;
  assign n2939 = n2929 & n2938;
  assign n2940 = n198 & ~n2533;
  assign n2941 = n2939 & ~n2940;
  assign n2942 = n2919 & n2941;
  assign n2943 = n2910 & n2942;
  assign n2944 = ~n2897 & n2943;
  assign n2945 = n497 & ~n2161;
  assign n2946 = ~n226 & ~n261;
  assign n2947 = ~n1931 & n2730;
  assign n2948 = n226 & ~n2947;
  assign n2949 = ~n274 & ~n2948;
  assign n2950 = ~n214 & n2949;
  assign n2951 = ~n2946 & ~n2950;
  assign n2952 = ~n717 & n1034;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~n2945 & n2953;
  assign n2955 = ~n226 & n735;
  assign n2956 = ~n273 & n1533;
  assign n2957 = n318 & ~n2956;
  assign n2958 = ~n1430 & n2509;
  assign n2959 = n261 & ~n2958;
  assign n2960 = ~n1219 & ~n2959;
  assign n2961 = n2721 & n2960;
  assign n2962 = ~n2957 & n2961;
  assign n2963 = ~n874 & n2962;
  assign n2964 = ~n2955 & ~n2963;
  assign n2965 = n2954 & ~n2964;
  assign n2966 = ~n226 & ~n318;
  assign n2967 = ~n1926 & n2339;
  assign n2968 = n318 & ~n2967;
  assign n2969 = ~n1432 & n2380;
  assign n2970 = n2232 & n2969;
  assign n2971 = ~n2968 & n2970;
  assign n2972 = ~n2966 & ~n2971;
  assign n2973 = ~n70 & n190;
  assign n2974 = i_12_ & i_14_;
  assign n2975 = ~n105 & ~n2974;
  assign n2976 = n429 & n2975;
  assign n2977 = ~n430 & ~n2976;
  assign n2978 = ~n2973 & n2977;
  assign n2979 = n232 & ~n2978;
  assign n2980 = ~i_13_ & n226;
  assign n2981 = n1938 & n2980;
  assign n2982 = n193 & ~n735;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2979 & n2983;
  assign n2985 = n974 & ~n2233;
  assign n2986 = ~i_8_ & n2985;
  assign n2987 = ~n232 & ~n261;
  assign n2988 = n1926 & ~n2987;
  assign n2989 = ~n1926 & n2196;
  assign n2990 = n496 & ~n2989;
  assign n2991 = n188 & n1951;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n2988 & n2992;
  assign n2994 = ~n2986 & n2993;
  assign n2995 = n2984 & n2994;
  assign n2996 = n261 & ~n2969;
  assign n2997 = ~n451 & n1009;
  assign n2998 = n1493 & n2314;
  assign n2999 = ~n717 & ~n2998;
  assign n3000 = ~n2997 & ~n2999;
  assign n3001 = ~n1772 & n3000;
  assign n3002 = ~n2996 & n3001;
  assign n3003 = n2995 & n3002;
  assign n3004 = ~n2972 & n3003;
  assign n3005 = n2124 & n2161;
  assign n3006 = n400 & ~n3005;
  assign n3007 = ~n580 & ~n2364;
  assign n3008 = ~n1420 & ~n1964;
  assign n3009 = ~n213 & ~n1673;
  assign n3010 = ~n419 & n3009;
  assign n3011 = n3008 & n3010;
  assign n3012 = n232 & ~n3011;
  assign n3013 = n232 & n1757;
  assign n3014 = n211 & n2904;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n3012 & n3015;
  assign n3017 = ~n3007 & n3016;
  assign n3018 = ~n1420 & ~n1430;
  assign n3019 = ~n2966 & ~n3018;
  assign n3020 = ~n2122 & ~n2926;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = n3017 & n3021;
  assign n3023 = ~i_8_ & n1100;
  assign n3024 = n335 & n735;
  assign n3025 = n1945 & ~n3024;
  assign n3026 = n1096 & ~n2935;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = ~n3023 & n3027;
  assign n3029 = n873 & ~n1135;
  assign n3030 = n3008 & n3029;
  assign n3031 = ~n2507 & n3030;
  assign n3032 = n295 & ~n3031;
  assign n3033 = ~n419 & ~n1176;
  assign n3034 = n238 & ~n3033;
  assign n3035 = ~n3032 & ~n3034;
  assign n3036 = n3028 & n3035;
  assign n3037 = n3022 & n3036;
  assign n3038 = ~n3006 & n3037;
  assign n3039 = n3004 & n3038;
  assign n3040 = n2965 & n3039;
  assign n3041 = ~n430 & ~n2353;
  assign n3042 = n1614 & n3041;
  assign n3043 = ~n1009 & ~n1107;
  assign n3044 = ~n458 & n3043;
  assign n3045 = n3042 & n3044;
  assign n3046 = ~n1083 & n3045;
  assign n3047 = n318 & ~n3046;
  assign n3048 = n2139 & ~n2249;
  assign n3049 = ~n390 & n3048;
  assign n3050 = n295 & ~n3049;
  assign n3051 = ~n2366 & ~n2987;
  assign n3052 = n92 & n1950;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = ~n2557 & n3053;
  assign n3055 = ~n3050 & n3054;
  assign n3056 = n496 & n613;
  assign n3057 = n232 & n1599;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = n2136 & n3058;
  assign n3060 = ~n797 & ~n1035;
  assign n3061 = n295 & ~n3060;
  assign n3062 = ~n1020 & ~n3061;
  assign n3063 = n451 & n717;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n2197 & n2258;
  assign n3066 = n261 & ~n3065;
  assign n3067 = ~n3064 & ~n3066;
  assign n3068 = n3059 & n3067;
  assign n3069 = n3055 & n3068;
  assign n3070 = ~n3047 & n3069;
  assign n3071 = ~n2286 & n3070;
  assign n3072 = n226 & n1941;
  assign n3073 = n261 & ~n3042;
  assign n3074 = n1014 & n3073;
  assign n3075 = ~n3072 & ~n3074;
  assign n3076 = ~n2162 & ~n2966;
  assign n3077 = n2231 & ~n3076;
  assign n3078 = n400 & ~n2134;
  assign n3079 = n3077 & ~n3078;
  assign n3080 = n3075 & n3079;
  assign n3081 = n738 & ~n1927;
  assign n3082 = ~n2518 & ~n3081;
  assign n3083 = n3080 & ~n3082;
  assign n3084 = ~n2534 & n3083;
  assign n3085 = n372 & n3081;
  assign n3086 = n1134 & ~n3085;
  assign n3087 = n2264 & ~n3086;
  assign n3088 = n3084 & n3087;
  assign n3089 = n3071 & n3088;
  assign n3090 = n3040 & n3089;
  assign n3091 = n2739 & n3090;
  assign o_36_ = ~n2944 | ~n3091;
  assign n3093 = n2744 & n2853;
  assign n3094 = n201 & ~n2888;
  assign n3095 = n296 & ~n579;
  assign n3096 = n232 & ~n2836;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = ~n3094 & n3097;
  assign n3099 = ~n2003 & n3098;
  assign n3100 = n221 & ~n2813;
  assign n3101 = n2558 & ~n3100;
  assign n3102 = ~n1666 & n3101;
  assign n3103 = ~n149 & n2904;
  assign n3104 = n115 & n3103;
  assign n3105 = n974 & n1800;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = n3102 & n3106;
  assign n3108 = ~n799 & n2836;
  assign n3109 = ~n1001 & ~n1985;
  assign n3110 = n2185 & n3109;
  assign n3111 = n3108 & n3110;
  assign n3112 = n1527 & n3111;
  assign n3113 = n226 & ~n3112;
  assign n3114 = n612 & n2183;
  assign n3115 = n496 & ~n3114;
  assign n3116 = n400 & ~n3109;
  assign n3117 = ~n3115 & ~n3116;
  assign n3118 = ~n3113 & n3117;
  assign n3119 = n1548 & n2187;
  assign n3120 = ~n1542 & ~n2079;
  assign n3121 = n2407 & ~n3120;
  assign n3122 = n3119 & n3121;
  assign n3123 = n261 & ~n1542;
  assign n3124 = n198 & n1647;
  assign n3125 = n703 & ~n3124;
  assign n3126 = ~n3123 & n3125;
  assign n3127 = n3122 & n3126;
  assign n3128 = n3118 & n3127;
  assign n3129 = n200 & ~n2185;
  assign n3130 = n318 & n1107;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = ~n609 & ~n999;
  assign n3133 = n2825 & n3132;
  assign n3134 = n3108 & n3133;
  assign n3135 = n295 & ~n3134;
  assign n3136 = n238 & ~n921;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = n3131 & n3137;
  assign n3139 = n3128 & n3138;
  assign n3140 = n3107 & n3139;
  assign n3141 = n3099 & n3140;
  assign n3142 = n3093 & n3141;
  assign n3143 = i_8_ & n1939;
  assign n3144 = n2312 & ~n3143;
  assign n3145 = n221 & ~n3144;
  assign n3146 = ~n1009 & n2222;
  assign n3147 = ~n193 & ~n1063;
  assign n3148 = n1398 & n3147;
  assign n3149 = n2969 & n3148;
  assign n3150 = n2223 & n2339;
  assign n3151 = n3149 & n3150;
  assign n3152 = ~n283 & n3151;
  assign n3153 = ~n3146 & ~n3152;
  assign n3154 = n763 & n2142;
  assign n3155 = ~n3153 & n3154;
  assign n3156 = n200 & ~n3155;
  assign n3157 = ~n431 & ~n825;
  assign n3158 = ~n3156 & n3157;
  assign n3159 = ~n3145 & n3158;
  assign n3160 = n2229 & n2703;
  assign n3161 = ~n2033 & n2403;
  assign n3162 = ~n793 & n2390;
  assign n3163 = n3161 & n3162;
  assign n3164 = n295 & ~n3163;
  assign n3165 = n2142 & ~n2300;
  assign n3166 = ~n221 & ~n344;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = n295 & n1397;
  assign n3169 = ~n694 & ~n3168;
  assign n3170 = ~n2569 & n3169;
  assign n3171 = ~n3167 & n3170;
  assign n3172 = ~n3164 & n3171;
  assign n3173 = n1717 & n2146;
  assign n3174 = ~n1940 & ~n2554;
  assign n3175 = n2624 & n3174;
  assign n3176 = ~n198 & ~n226;
  assign n3177 = n1992 & ~n3176;
  assign n3178 = ~n2629 & ~n3177;
  assign n3179 = n3175 & n3178;
  assign n3180 = n3173 & n3179;
  assign n3181 = n3172 & n3180;
  assign n3182 = n2546 & n3181;
  assign n3183 = n256 & ~n2312;
  assign n3184 = ~n2405 & ~n3183;
  assign n3185 = n3182 & n3184;
  assign n3186 = n3160 & n3185;
  assign n3187 = n2318 & n3186;
  assign n3188 = n3159 & n3187;
  assign n3189 = ~n594 & ~n2184;
  assign n3190 = ~n1277 & ~n2116;
  assign n3191 = ~n2279 & ~n3190;
  assign n3192 = ~n3189 & n3191;
  assign n3193 = n2687 & n3004;
  assign n3194 = n3192 & n3193;
  assign n3195 = n2944 & n3194;
  assign n3196 = n3188 & n3195;
  assign o_37_ = ~n3142 | ~n3196;
  assign n3198 = ~n1283 & ~n2290;
  assign n3199 = n233 & n3103;
  assign n3200 = ~n1277 & ~n2118;
  assign n3201 = ~n1002 & ~n1958;
  assign n3202 = n400 & ~n3201;
  assign n3203 = n233 & n388;
  assign n3204 = ~n2745 & ~n3203;
  assign n3205 = n238 & ~n3204;
  assign n3206 = ~n3202 & ~n3205;
  assign n3207 = ~n3200 & n3206;
  assign n3208 = ~n3199 & n3207;
  assign n3209 = ~n3198 & n3208;
  assign n3210 = n2736 & n3209;
  assign n3211 = n808 & n2774;
  assign n3212 = n2036 & n3211;
  assign n3213 = n232 & ~n3212;
  assign n3214 = ~n2001 & ~n2111;
  assign n3215 = n226 & ~n2776;
  assign n3216 = n295 & ~n2775;
  assign n3217 = ~n2294 & ~n3216;
  assign n3218 = ~n3215 & n3217;
  assign n3219 = ~n3214 & n3218;
  assign n3220 = ~n3213 & n3219;
  assign n3221 = n1540 & n2551;
  assign n3222 = n297 & n808;
  assign n3223 = n1927 & ~n3222;
  assign n3224 = ~n2082 & ~n3223;
  assign n3225 = n412 & n2340;
  assign n3226 = n261 & ~n3225;
  assign n3227 = ~n766 & ~n2377;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = n3224 & n3228;
  assign n3230 = ~n1536 & n2212;
  assign n3231 = n497 & ~n3230;
  assign n3232 = ~n402 & ~n3231;
  assign n3233 = n3229 & n3232;
  assign n3234 = n3221 & n3233;
  assign n3235 = n3220 & n3234;
  assign n3236 = n3210 & n3235;
  assign n3237 = n2785 & n3040;
  assign n3238 = n3236 & n3237;
  assign o_38_ = ~n3188 | ~n3238;
  assign n3240 = ~n2733 & ~n2762;
  assign n3241 = ~n667 & n1580;
  assign n3242 = ~n523 & n3241;
  assign n3243 = ~n1185 & n3242;
  assign n3244 = n3240 & n3243;
  assign n3245 = n2076 & n2730;
  assign n3246 = ~n575 & ~n1945;
  assign n3247 = ~n1002 & n3246;
  assign n3248 = ~n419 & n3247;
  assign n3249 = n1097 & n1903;
  assign n3250 = n3248 & n3249;
  assign n3251 = n3245 & n3250;
  assign n3252 = n238 & ~n3251;
  assign n3253 = n3244 & ~n3252;
  assign n3254 = ~n428 & ~n1051;
  assign n3255 = n927 & n3254;
  assign o_39_ = ~n3253 | ~n3255;
  assign n3257 = n71 & ~n2447;
  assign n3258 = ~i_6_ & n2592;
  assign o_40_ = n3257 | n3258;
  assign n3260 = n73 & n217;
  assign o_41_ = n67 & n3260;
  assign o_42_ = n657 & n2180;
  assign n3263 = ~n1684 & n1954;
  assign n3264 = n1222 & ~n2726;
  assign n3265 = n1551 & n3264;
  assign n3266 = n3263 & n3265;
  assign n3267 = ~n2051 & n2189;
  assign n3268 = i_8_ & ~n3267;
  assign n3269 = ~n1007 & ~n1561;
  assign n3270 = ~n1083 & n3269;
  assign n3271 = n2257 & n3270;
  assign n3272 = ~n3268 & n3271;
  assign n3273 = n2120 & n3272;
  assign n3274 = ~n314 & n3273;
  assign n3275 = n200 & ~n3274;
  assign n3276 = ~n1096 & n2365;
  assign n3277 = n612 & ~n1935;
  assign n3278 = n2328 & n3277;
  assign n3279 = n2380 & n2398;
  assign n3280 = ~n2051 & n2122;
  assign n3281 = n3279 & n3280;
  assign n3282 = n3278 & n3281;
  assign n3283 = n3276 & n3282;
  assign n3284 = n2339 & n3283;
  assign n3285 = n318 & ~n3284;
  assign n3286 = ~n2688 & ~n3285;
  assign n3287 = n481 & n3131;
  assign n3288 = n851 & n3287;
  assign n3289 = n3286 & n3288;
  assign n3290 = ~n3275 & n3289;
  assign n3291 = n3158 & n3290;
  assign n3292 = n3266 & n3291;
  assign n3293 = n2256 & ~n2912;
  assign n3294 = ~n2274 & n3293;
  assign o_43_ = ~n3292 | ~n3294;
  assign n3296 = n2202 & n3011;
  assign n3297 = ~n117 & n2258;
  assign n3298 = n3296 & n3297;
  assign n3299 = n3212 & n3298;
  assign n3300 = n2376 & n3299;
  assign n3301 = n232 & ~n3300;
  assign n3302 = ~n2845 & ~n2979;
  assign n3303 = ~n2698 & n3302;
  assign n3304 = ~n2655 & n3303;
  assign n3305 = ~o_16_ & n3304;
  assign n3306 = n2919 & n3305;
  assign n3307 = ~n3301 & n3306;
  assign n3308 = ~n211 & ~n821;
  assign n3309 = i_8_ & ~n3308;
  assign n3310 = ~n1107 & n2235;
  assign n3311 = ~n3309 & n3310;
  assign n3312 = n2813 & n3311;
  assign n3313 = n3165 & n3312;
  assign n3314 = n2114 & n2234;
  assign n3315 = n1512 & n2167;
  assign n3316 = n2213 & n3315;
  assign n3317 = n3314 & n3316;
  assign n3318 = ~n810 & ~n1958;
  assign n3319 = n2271 & n3318;
  assign n3320 = n3317 & n3319;
  assign n3321 = n2109 & n3320;
  assign n3322 = i_8_ & ~n3321;
  assign n3323 = n3144 & ~n3322;
  assign n3324 = n3313 & n3323;
  assign n3325 = n221 & ~n3324;
  assign n3326 = n3292 & ~n3325;
  assign o_44_ = ~n3307 | ~n3326;
  assign n3328 = ~n108 & ~n2469;
  assign o_45_ = ~n2590 | n3328;
endmodule


