// Benchmark "rot" written by ABC on Tue May 16 16:07:52 2017

module rot ( 
    z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r,
    s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4, c0, c1,
    c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2, f3, g0,
    g1, g2, g3, h0, h1, h2, h3, i0, i1, i2, i3, j0, j1, j2, j3, k0, k1, k2,
    k3, l0, l1, l2, l3, m0, m1, m2, m3, n0, n1, n2, n3, o0, o1, o2, o3, p0,
    p1, p2, p3, q0, q1, q2, q3, r0, r1, r2, r3, s0, s1, s2, s3, t0, t1, t2,
    t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2, w3, x0, x1, x2, x3, y0,
    y1, y2, y3,
    z4, z5, z6, z7, a5, a6, a7, a8, b5, b6, b7, b8, c5, c6, c7, c8, d5, d6,
    d7, d8, e5, e6, e7, e8, f4, f5, f6, f7, f8, g4, g5, g6, g7, g8, h4, h5,
    h6, h7, h8, i4, i5, i6, i7, j4, j5, j6, j7, k4, k5, k6, k7, l4, l5, l6,
    l7, m4, m5, m6, m7, n4, n5, n6, n7, o4, o5, o6, o7, p4, p5, p6, p7, q4,
    q5, q6, q7, r4, r5, r6, r7, s4, s5, s6, s7, t4, t5, t6, t7, u4, u5, u6,
    u7, v4, v5, v6, v7, w4, w5, w6, w7, x4, x5, x6, x7, y4, y5, y6, y7  );
  input  z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p,
    q, r, s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4,
    c0, c1, c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2,
    f3, g0, g1, g2, g3, h0, h1, h2, h3, i0, i1, i2, i3, j0, j1, j2, j3, k0,
    k1, k2, k3, l0, l1, l2, l3, m0, m1, m2, m3, n0, n1, n2, n3, o0, o1, o2,
    o3, p0, p1, p2, p3, q0, q1, q2, q3, r0, r1, r2, r3, s0, s1, s2, s3, t0,
    t1, t2, t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2, w3, x0, x1, x2,
    x3, y0, y1, y2, y3;
  output z4, z5, z6, z7, a5, a6, a7, a8, b5, b6, b7, b8, c5, c6, c7, c8, d5,
    d6, d7, d8, e5, e6, e7, e8, f4, f5, f6, f7, f8, g4, g5, g6, g7, g8, h4,
    h5, h6, h7, h8, i4, i5, i6, i7, j4, j5, j6, j7, k4, k5, k6, k7, l4, l5,
    l6, l7, m4, m5, m6, m7, n4, n5, n6, n7, o4, o5, o6, o7, p4, p5, p6, p7,
    q4, q5, q6, q7, r4, r5, r6, r7, s4, s5, s6, s7, t4, t5, t6, t7, u4, u5,
    u6, u7, v4, v5, v6, v7, w4, w5, w6, w7, x4, x5, x6, x7, y4, y5, y6, y7;
  wire n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n278, n279,
    n282, n283, n285, n286, n287, n289, n291, n292, n294, n295, n296, n298,
    n299, n301, n302, n303, n305, n306, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n354, n356, n357, n358, n359, n360, n361, n363, n366,
    n370, n371, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n392, n393, n395, n398, n399,
    n400, n402, n404, n405, n407, n408, n410, n411, n412, n413, n414, n415,
    n416, n418, n419, n420, n421, n422, n423, n424, n427, n428, n429, n430,
    n431, n433, n434, n435, n436, n437, n439, n440, n442, n443, n444, n445,
    n446, n447, n448, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n489, n490, n492, n493, n494, n495, n496,
    n501, n503, n504, n505, n506, n507, n508, n509, n510, n511, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n556, n557, n558, n559, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n579, n583, n584, n585, n586, n587, n589, n590, n591, n592, n594,
    n595, n596, n598, n599, n601, n602, n603, n606, n607, n608, n609, n610,
    n611, n612, n613, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n703, n704, n705, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n733, n734, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n770, n772, n773, n774, n777, n778, n779,
    n781, n782, n784, n785, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n813, n814, n815, n817, n818, n819, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n838, n839, n840, n841, n842, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n869, n870, n871, n872, n873, n874,
    n876, n877, n878, n879, n880, n881, n882, n884, n885, n886, n888, n889,
    n890, n891, n893, n895;
  assign z4 = b4 & v0;
  assign n244 = ~h0 & t0;
  assign n245 = n3 & n244;
  assign n246 = h0 & ~s0;
  assign n247 = u & s0;
  assign n248 = ~n246 & ~n247;
  assign n249 = ~m & ~d0;
  assign n250 = u2 & n249;
  assign n251 = ~w2 & n250;
  assign n252 = x2 & n251;
  assign n253 = n248 & n252;
  assign n254 = ~k & d0;
  assign n255 = u2 & n254;
  assign n256 = ~w2 & n255;
  assign n257 = x2 & n256;
  assign n258 = n248 & n257;
  assign n259 = ~h & u2;
  assign n260 = u3 & n259;
  assign n261 = n248 & n260;
  assign n262 = ~i & u3;
  assign n263 = ~l & ~d0;
  assign n264 = ~j & d0;
  assign n265 = g & ~n264;
  assign n266 = ~n263 & n265;
  assign n267 = ~n262 & n266;
  assign n268 = ~n261 & n267;
  assign n269 = ~n258 & n268;
  assign n270 = ~n253 & n269;
  assign n271 = m2 & y1;
  assign n272 = x1 & n271;
  assign n273 = w2 & n270;
  assign n274 = x2 & ~n272;
  assign n275 = w2 & ~x2;
  assign n276 = ~n274 & ~n275;
  assign d8 = n273 | ~n276;
  assign n278 = ~i2 & ~k2;
  assign n279 = ~d8 & n278;
  assign z5 = n245 | ~n279;
  assign z6 = ~z0 & ~y0;
  assign n282 = k & ~d0;
  assign n283 = m & d0;
  assign z7 = n282 | n283;
  assign n285 = ~x & y;
  assign n286 = e0 & n285;
  assign n287 = n0 & ~n285;
  assign a6 = n286 | n287;
  assign n289 = ~n270 & n272;
  assign a8 = c4 | n289;
  assign n291 = ~c1 & d1;
  assign n292 = c1 & ~d1;
  assign b5 = n291 | n292;
  assign n294 = ~q2 & ~r0;
  assign n295 = m2 & ~n294;
  assign n296 = m1 & m2;
  assign b6 = n295 | n296;
  assign n298 = ~w2 & x2;
  assign n299 = n272 & n298;
  assign b8 = n270 & n299;
  assign n301 = c1 & d1;
  assign n302 = e1 & ~n301;
  assign n303 = ~e1 & n301;
  assign c5 = n302 | n303;
  assign n305 = x1 & ~y1;
  assign n306 = m2 & n305;
  assign c6 = w1 & n306;
  assign n308 = p2 & q2;
  assign n309 = l2 & n308;
  assign n310 = ~f2 & ~h2;
  assign n311 = f2 & ~g2;
  assign n312 = ~h2 & n311;
  assign n313 = ~f2 & ~g2;
  assign n314 = h2 & n313;
  assign n315 = ~n312 & ~n314;
  assign n316 = l2 & ~n315;
  assign n317 = ~z1 & ~n316;
  assign n318 = ~r1 & s1;
  assign n319 = ~p1 & r1;
  assign n320 = ~s1 & n319;
  assign n321 = o2 & n320;
  assign n322 = ~n317 & n321;
  assign n323 = ~n310 & n322;
  assign n324 = o2 & ~p1;
  assign n325 = ~n317 & n324;
  assign n326 = ~n310 & n325;
  assign n327 = n318 & n326;
  assign n328 = ~n323 & ~n327;
  assign n329 = o1 & ~y3;
  assign n330 = n328 & n329;
  assign n331 = ~n309 & n330;
  assign n332 = o1 & ~s1;
  assign n333 = ~y3 & n332;
  assign n334 = ~n309 & n333;
  assign n335 = ~q & o1;
  assign n336 = ~y3 & n335;
  assign n337 = n328 & n336;
  assign n338 = ~s1 & n335;
  assign n339 = ~y3 & n338;
  assign n340 = m1 & n328;
  assign n341 = ~n309 & n340;
  assign n342 = m1 & ~s1;
  assign n343 = ~n309 & n342;
  assign n344 = ~q & m1;
  assign n345 = n328 & n344;
  assign n346 = ~s1 & n344;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n343 & n347;
  assign n349 = ~n341 & n348;
  assign n350 = ~n339 & n349;
  assign n351 = ~n337 & n350;
  assign n352 = ~n334 & n351;
  assign c7 = n331 | ~n352;
  assign n354 = w2 & ~n272;
  assign c8 = ~a4 | n354;
  assign n356 = ~q & l2;
  assign n357 = p & l2;
  assign n358 = ~n & l2;
  assign n359 = ~n356 & ~n358;
  assign n360 = ~n357 & n359;
  assign n361 = ~c1 & l2;
  assign j5 = ~n360 | n361;
  assign n363 = ~d1 & l2;
  assign i5 = ~n360 | n363;
  assign h5 = j5 & i5;
  assign n366 = ~e1 & l2;
  assign g5 = ~n360 | n366;
  assign f5 = j5 & g5;
  assign d5 = h5 & f5;
  assign n370 = ~p2 & q2;
  assign n371 = p2 & ~q2;
  assign e6 = n370 | n371;
  assign n373 = m1 & o1;
  assign n374 = ~y3 & n373;
  assign n375 = c7 & n374;
  assign n376 = i1 & m1;
  assign n377 = c7 & n376;
  assign n378 = n329 & e6;
  assign n379 = ~l2 & o1;
  assign n380 = ~y3 & n379;
  assign n381 = i1 & e6;
  assign n382 = i1 & ~l2;
  assign n383 = ~q & i1;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n381 & n384;
  assign n386 = ~n336 & n385;
  assign n387 = ~n380 & n386;
  assign n388 = ~n378 & n387;
  assign n389 = ~n377 & n388;
  assign d7 = n375 | ~n389;
  assign e5 = i5 & g5;
  assign n392 = ~s & ~l3;
  assign n393 = e4 & i1;
  assign i7 = y3 & n393;
  assign n395 = z3 & i7;
  assign e7 = ~n392 & n395;
  assign e8 = ~w0 & ~x0;
  assign n398 = x & ~y;
  assign n399 = j1 & n398;
  assign n400 = e0 & ~n398;
  assign f4 = n399 | n400;
  assign n402 = m2 & p2;
  assign f6 = n295 | n402;
  assign n404 = m2 & q2;
  assign n405 = ~n296 & ~n402;
  assign f7 = n404 | ~n405;
  assign n407 = p0 & ~y1;
  assign n408 = k1 & y1;
  assign g4 = n407 | n408;
  assign n410 = r0 & ~n308;
  assign n411 = n306 & n410;
  assign n412 = p & ~m2;
  assign n413 = n308 & n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = v3 & n414;
  assign n416 = ~p0 & ~n414;
  assign g6 = n415 | n416;
  assign n418 = ~x1 & n271;
  assign n419 = q & ~m2;
  assign n420 = n308 & n419;
  assign n421 = ~n308 & n418;
  assign n422 = ~n420 & ~n421;
  assign n423 = q3 & n422;
  assign n424 = ~k1 & ~n422;
  assign g7 = n423 | n424;
  assign h4 = v2 | d8;
  assign n427 = p0 & ~n414;
  assign n428 = ~q0 & n427;
  assign n429 = q0 & n416;
  assign n430 = w3 & n414;
  assign n431 = ~n429 & ~n430;
  assign h6 = n428 | ~n431;
  assign n433 = k1 & ~n422;
  assign n434 = ~l1 & n433;
  assign n435 = l1 & n424;
  assign n436 = r3 & n422;
  assign n437 = ~n435 & ~n436;
  assign h7 = n434 | ~n437;
  assign n439 = ~w2 & d8;
  assign n440 = ~w2 & ~x2;
  assign h8 = n439 | n440;
  assign n442 = ~g0 & h0;
  assign n443 = u2 & n442;
  assign n444 = ~s0 & n443;
  assign n445 = ~t & u;
  assign n446 = u2 & n445;
  assign n447 = s0 & n446;
  assign n448 = ~d8 & ~n447;
  assign i4 = n444 | ~n448;
  assign n450 = ~w0 & z6;
  assign n451 = ~e8 & n450;
  assign n452 = z0 & w0;
  assign n453 = ~z0 & ~z6;
  assign n454 = e8 & n453;
  assign n455 = ~n452 & ~n454;
  assign n456 = ~n451 & n455;
  assign n457 = ~x0 & y0;
  assign n458 = u1 & n457;
  assign n459 = ~e8 & n458;
  assign n460 = n456 & n459;
  assign n461 = x0 & ~y0;
  assign n462 = u1 & n461;
  assign n463 = ~z6 & n462;
  assign n464 = n456 & n463;
  assign n465 = x0 & y0;
  assign n466 = u1 & n465;
  assign n467 = ~n456 & n466;
  assign n468 = u1 & z6;
  assign n469 = e8 & n468;
  assign n470 = ~n467 & ~n469;
  assign n471 = ~n464 & n470;
  assign n472 = ~n460 & n471;
  assign n473 = n456 & n472;
  assign n474 = j2 & ~n473;
  assign n475 = ~n3 & ~o3;
  assign n476 = ~t3 & n475;
  assign n477 = a2 & ~n476;
  assign n478 = k0 & l0;
  assign n479 = m0 & n478;
  assign n480 = n477 & n479;
  assign n481 = ~n474 & n480;
  assign n482 = ~n245 & n481;
  assign n483 = j0 & k0;
  assign n484 = l0 & n483;
  assign n485 = m0 & n484;
  assign n486 = ~n474 & n485;
  assign n487 = ~n482 & ~n486;
  assign i6 = l3 & ~n487;
  assign n489 = u2 & ~n248;
  assign n490 = c2 & d8;
  assign j4 = n489 | n490;
  assign n492 = r1 & ~n328;
  assign n493 = t0 & n442;
  assign n494 = ~l3 & n493;
  assign n495 = r0 & ~n492;
  assign n496 = ~n309 & n495;
  assign j6 = n494 | n496;
  assign j7 = ~m1 & ~d8;
  assign k6 = ~k2 & ~m0;
  assign k7 = i1 | n418;
  assign n501 = n & e1;
  assign l5 = n301 & n501;
  assign n503 = ~h3 & i3;
  assign n504 = h3 & ~i3;
  assign n505 = ~n503 & ~n504;
  assign n506 = ~k2 & m2;
  assign n507 = n505 & n506;
  assign n508 = ~i3 & n506;
  assign n509 = ~k2 & p2;
  assign n510 = ~k6 & ~n509;
  assign n511 = ~n508 & n510;
  assign l6 = n507 | ~n511;
  assign n513 = ~n328 & ~j4;
  assign n514 = a & f0;
  assign n515 = r2 & ~n514;
  assign n516 = ~n513 & n515;
  assign n517 = m3 & ~n505;
  assign n518 = b2 & ~d8;
  assign n519 = v1 & n518;
  assign n520 = n517 & ~n519;
  assign n521 = f3 & ~n519;
  assign n522 = e3 & ~n519;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n520 & n523;
  assign n525 = y2 & ~n524;
  assign n526 = ~z3 & ~d8;
  assign n527 = g3 & ~n524;
  assign n528 = ~n492 & n527;
  assign n529 = b2 & ~s1;
  assign n530 = s0 & ~n529;
  assign n531 = n1 & ~n318;
  assign n532 = n1 & ~n518;
  assign n533 = ~n531 & ~n532;
  assign n534 = y3 & n533;
  assign n535 = ~d8 & n534;
  assign n536 = h4 & ~n535;
  assign n537 = n526 & n528;
  assign n538 = n525 & n537;
  assign n539 = u2 & n526;
  assign n540 = n392 & n539;
  assign n541 = u2 & n530;
  assign n542 = n526 & n541;
  assign n543 = n526 & n536;
  assign n544 = n272 & d8;
  assign n545 = ~x2 & ~h8;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n543 & n546;
  assign n548 = ~n542 & n547;
  assign n549 = ~n540 & n548;
  assign n550 = ~n538 & n549;
  assign n551 = ~n516 & ~n550;
  assign n552 = u2 & n551;
  assign n553 = s & ~l3;
  assign n554 = ~n528 & ~n553;
  assign l7 = n552 | ~n554;
  assign n556 = d & e;
  assign n557 = f & n556;
  assign n558 = n318 & ~n557;
  assign n559 = b1 & ~n557;
  assign m5 = n558 | n559;
  assign n561 = ~z2 & ~a3;
  assign n562 = ~b3 & ~c3;
  assign n563 = ~d3 & n562;
  assign n564 = l2 & o0;
  assign n565 = d3 & n564;
  assign n566 = ~c3 & n564;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n563 & n567;
  assign n569 = n561 & n568;
  assign n570 = m3 & ~n492;
  assign n571 = n569 & n570;
  assign n572 = h3 & i3;
  assign n573 = n569 & n572;
  assign n574 = ~n571 & ~n573;
  assign n575 = n244 & n569;
  assign n576 = h3 & ~n574;
  assign n577 = ~n494 & ~n575;
  assign m6 = n576 | ~n577;
  assign n579 = n476 & ~n528;
  assign o7 = ~n533 | n579;
  assign m7 = ~n528 & ~o7;
  assign o4 = w1 & n272;
  assign n583 = n418 & l5;
  assign n584 = ~n & n418;
  assign n585 = n272 & ~o4;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n583 & n586;
  assign n4 = n411 | ~n587;
  assign n589 = g2 & l2;
  assign n590 = ~h2 & ~l2;
  assign n591 = f2 & l2;
  assign n592 = ~n589 & ~n591;
  assign p5 = n590 | ~n592;
  assign n594 = ~g2 & ~l2;
  assign n595 = ~p5 & n594;
  assign n596 = f2 & ~p5;
  assign o5 = n595 | n596;
  assign n598 = ~l2 & ~o5;
  assign n599 = ~p5 & n598;
  assign n5 = a | n599;
  assign n601 = n504 & n574;
  assign n602 = i3 & ~n574;
  assign n603 = ~n575 & ~n602;
  assign n6 = n601 | ~n603;
  assign n7 = n528 & n533;
  assign n606 = ~n492 & ~n569;
  assign n607 = n517 & n606;
  assign n608 = ~n569 & n572;
  assign n609 = ~n607 & ~n608;
  assign n610 = n248 & ~n609;
  assign n611 = z2 & n505;
  assign n612 = z2 & n609;
  assign n613 = ~n610 & ~n612;
  assign o6 = n611 | ~n613;
  assign n615 = ~t1 & t2;
  assign n616 = ~a & n551;
  assign n617 = ~n615 & n616;
  assign n618 = ~n317 & n617;
  assign n619 = ~n589 & n618;
  assign n620 = ~a & n516;
  assign n621 = ~n615 & n620;
  assign n622 = ~n317 & n621;
  assign n623 = ~n589 & n622;
  assign n624 = ~h2 & ~n5;
  assign n625 = n551 & n624;
  assign n626 = ~n615 & n625;
  assign n627 = ~n317 & n626;
  assign n628 = ~f2 & ~n5;
  assign n629 = n551 & n628;
  assign n630 = ~n615 & n629;
  assign n631 = ~n317 & n630;
  assign n632 = n516 & n624;
  assign n633 = ~n615 & n632;
  assign n634 = ~n317 & n633;
  assign n635 = n516 & n628;
  assign n636 = ~n615 & n635;
  assign n637 = ~n317 & n636;
  assign n638 = n551 & ~n5;
  assign n639 = ~n615 & n638;
  assign n640 = n310 & n639;
  assign n641 = n516 & ~n5;
  assign n642 = ~n615 & n641;
  assign n643 = n310 & n642;
  assign n644 = ~n640 & ~n643;
  assign n645 = ~n637 & n644;
  assign n646 = ~n634 & n645;
  assign n647 = ~n631 & n646;
  assign n648 = ~n627 & n647;
  assign n649 = ~n623 & n648;
  assign p4 = n619 | ~n649;
  assign n651 = i0 & ~s0;
  assign n652 = n610 & n651;
  assign n653 = v & s0;
  assign n654 = n610 & n653;
  assign n655 = a3 & ~n492;
  assign n656 = ~n610 & n655;
  assign n657 = ~n505 & ~n609;
  assign n658 = a3 & o6;
  assign n659 = ~n610 & n658;
  assign n660 = ~n657 & ~n659;
  assign n661 = ~n656 & n660;
  assign n662 = ~n654 & n661;
  assign p6 = n652 | ~n662;
  assign n664 = s & ~n530;
  assign n665 = u2 & ~n664;
  assign n666 = a4 & l3;
  assign n667 = ~n528 & n666;
  assign n668 = ~n530 & n667;
  assign n669 = ~n536 & n668;
  assign n670 = n393 & n669;
  assign n671 = a4 & ~n528;
  assign n672 = ~n665 & n671;
  assign n673 = ~n536 & n672;
  assign n674 = n393 & n673;
  assign n675 = a4 & ~n487;
  assign n676 = ~n528 & n675;
  assign n677 = ~n665 & n676;
  assign n678 = ~n536 & n677;
  assign n679 = a4 & i6;
  assign n680 = ~n528 & n679;
  assign n681 = ~n530 & n680;
  assign n682 = ~n536 & n681;
  assign n683 = a4 & ~d8;
  assign n684 = ~n516 & n683;
  assign n685 = n393 & n684;
  assign n686 = a4 & n528;
  assign n687 = ~n536 & n686;
  assign n688 = ~n525 & n687;
  assign n689 = ~n533 & n684;
  assign n690 = n528 & n684;
  assign n691 = ~n487 & n684;
  assign n692 = a4 & ~n533;
  assign n693 = ~n536 & n692;
  assign n694 = ~n691 & ~n693;
  assign n695 = ~n690 & n694;
  assign n696 = ~n689 & n695;
  assign n697 = ~n688 & n696;
  assign n698 = ~n685 & n697;
  assign n699 = ~n682 & n698;
  assign n700 = ~n678 & n699;
  assign n701 = ~n674 & n700;
  assign p7 = n670 | ~n701;
  assign n703 = a1 & t2;
  assign n704 = ~a & n615;
  assign n705 = n310 & n704;
  assign q4 = n703 | n705;
  assign w5 = n3 & ~n487;
  assign n708 = g0 & t0;
  assign n709 = u2 & ~n516;
  assign n710 = n477 & n561;
  assign n711 = ~l2 & n477;
  assign n712 = ~n472 & n711;
  assign n713 = n708 & n712;
  assign n714 = ~l3 & t0;
  assign n715 = n477 & n714;
  assign n716 = ~n709 & n715;
  assign n717 = ~l3 & n244;
  assign n718 = n710 & n717;
  assign n719 = n248 & ~n526;
  assign n720 = ~n505 & n574;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n718 & n721;
  assign n723 = ~n716 & n722;
  assign n724 = ~n713 & n723;
  assign n725 = n244 & w5;
  assign n726 = n477 & n487;
  assign n727 = j0 & n487;
  assign n728 = ~n487 & ~n724;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n726 & n729;
  assign q5 = n725 | ~n730;
  assign q6 = b3 & ~o0;
  assign n733 = ~d4 & ~d8;
  assign n734 = ~n289 & n733;
  assign q7 = ~s1 & ~n734;
  assign n736 = ~o & ~p;
  assign n737 = ~q & n736;
  assign n738 = h2 & n737;
  assign n739 = ~o0 & ~n738;
  assign n740 = a & ~f1;
  assign n741 = ~g1 & n740;
  assign n742 = ~h1 & n741;
  assign n743 = ~q1 & n742;
  assign n744 = ~r1 & n743;
  assign n745 = ~h2 & n744;
  assign n746 = ~n318 & n745;
  assign n747 = ~q1 & ~r1;
  assign n748 = n315 & n747;
  assign n749 = ~n739 & n748;
  assign n750 = ~n318 & n749;
  assign n751 = ~n589 & n750;
  assign n752 = a & ~q1;
  assign n753 = ~r1 & n752;
  assign n754 = ~n739 & n753;
  assign n755 = ~n318 & n754;
  assign n756 = ~n589 & n755;
  assign n757 = ~h2 & n753;
  assign n758 = ~n318 & n757;
  assign n759 = ~n589 & n758;
  assign n760 = ~f1 & ~g1;
  assign n761 = ~h1 & n760;
  assign n762 = ~n739 & n761;
  assign n763 = n589 & n762;
  assign n764 = ~l2 & ~n739;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~n759 & n765;
  assign n767 = ~n756 & n766;
  assign n768 = ~n751 & n767;
  assign r4 = n746 | ~n768;
  assign n770 = ~n494 & n724;
  assign r5 = ~n487 & n770;
  assign n772 = c3 & ~n492;
  assign n773 = ~o0 & n772;
  assign n774 = c3 & q6;
  assign r6 = n773 | n774;
  assign r7 = n318 & ~n734;
  assign n777 = ~a & f0;
  assign n778 = ~a & j4;
  assign n779 = ~n328 & n778;
  assign s4 = n777 | n779;
  assign n781 = j2 & n473;
  assign n782 = ~o3 & n477;
  assign s5 = n781 | n782;
  assign n784 = d3 & ~o0;
  assign n785 = c3 & o0;
  assign s6 = n784 | n785;
  assign n787 = a & n557;
  assign n788 = a & ~n318;
  assign n789 = a & ~n;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n787 & n790;
  assign n792 = o2 & ~n791;
  assign n793 = n2 & ~n791;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n2 & ~n794;
  assign n796 = ~h4 & i4;
  assign n797 = h4 & ~i4;
  assign n798 = ~n796 & ~n797;
  assign n799 = ~i4 & n651;
  assign n800 = n551 & n799;
  assign n801 = ~i4 & n653;
  assign n802 = n551 & n801;
  assign n803 = n2 & ~n551;
  assign n804 = n794 & n803;
  assign n805 = ~n551 & n795;
  assign n806 = n551 & ~n798;
  assign n807 = n525 & n551;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~n805 & n808;
  assign n810 = ~n804 & n809;
  assign n811 = ~n802 & n810;
  assign t4 = n800 | ~n811;
  assign n813 = k0 & ~n710;
  assign n814 = h0 & k0;
  assign n815 = ~l2 & ~n814;
  assign t5 = n813 | ~n815;
  assign n817 = o & ~p;
  assign n818 = n356 & n817;
  assign n819 = ~k2 & n818;
  assign t6 = n781 | n819;
  assign n821 = f3 & ~i3;
  assign n822 = n551 & n821;
  assign n823 = n525 & n822;
  assign n824 = n517 & n823;
  assign n825 = e3 & i3;
  assign n826 = n551 & n825;
  assign n827 = n525 & n826;
  assign n828 = n517 & n827;
  assign n829 = e3 & f3;
  assign n830 = n551 & n829;
  assign n831 = n525 & n830;
  assign n832 = o2 & ~n551;
  assign n833 = ~n795 & n832;
  assign n834 = ~n806 & ~n833;
  assign n835 = ~n831 & n834;
  assign n836 = ~n828 & n835;
  assign u4 = n824 | ~n836;
  assign n838 = l0 & n709;
  assign n839 = l0 & ~n477;
  assign n840 = l0 & ~s0;
  assign n841 = n317 & ~n840;
  assign n842 = ~n839 & n841;
  assign u5 = n838 | ~n842;
  assign u6 = n472 & n708;
  assign n845 = ~n550 & n791;
  assign n846 = ~n514 & n845;
  assign n847 = ~n513 & n846;
  assign n848 = ~n550 & ~n794;
  assign n849 = ~n514 & n848;
  assign n850 = ~n513 & n849;
  assign n851 = n516 & ~n794;
  assign n852 = n516 & n791;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n850 & n853;
  assign v4 = n847 | ~n854;
  assign n856 = ~o & p;
  assign n857 = ~n494 & n856;
  assign n858 = n356 & n857;
  assign n859 = ~n503 & n858;
  assign n860 = p & p2;
  assign n861 = ~n494 & n860;
  assign n862 = n356 & n861;
  assign n863 = ~w1 & ~n494;
  assign n864 = n306 & n863;
  assign n865 = m0 & ~n494;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n862 & n866;
  assign v5 = n859 | ~n867;
  assign n869 = b & ~n551;
  assign n870 = n791 & n869;
  assign n871 = d2 & n551;
  assign n872 = ~b & ~n551;
  assign n873 = ~n791 & n872;
  assign n874 = ~n871 & ~n873;
  assign w4 = n870 | ~n874;
  assign n876 = b & ~n791;
  assign n877 = ~c & ~n551;
  assign n878 = n876 & n877;
  assign n879 = c & ~n551;
  assign n880 = ~n876 & n879;
  assign n881 = e2 & n551;
  assign n882 = ~n880 & ~n881;
  assign x4 = n878 | ~n882;
  assign n884 = k2 & ~n818;
  assign n885 = ~l2 & ~n472;
  assign n886 = n708 & n885;
  assign x5 = n884 | n886;
  assign n888 = r & ~p3;
  assign n889 = s2 & u0;
  assign n890 = r & k3;
  assign n891 = ~n889 & ~n890;
  assign x7 = n888 | ~n891;
  assign n893 = v0 & ~x3;
  assign y4 = a | n893;
  assign n895 = l3 & n708;
  assign y5 = n474 | n895;
  assign y7 = j3 & p3;
  assign d6 = ~p2;
  assign l4 = ~o3;
  assign a5 = m2;
  assign a7 = y0;
  assign b7 = z0;
  assign f8 = w0;
  assign g8 = x0;
  assign k4 = s3;
  assign k5 = l2;
  assign m4 = t3;
  assign s7 = w;
  assign t7 = z;
  assign u7 = a0;
  assign v6 = z6;
  assign v7 = b0;
  assign w6 = y0;
  assign w7 = c0;
  assign x6 = e8;
  assign y6 = w0;
endmodule


