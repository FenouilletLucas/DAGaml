// Benchmark "b9" written by ABC on Tue May 16 16:07:44 2017

module b9 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, p0, q0, r0, s0, t0, u0, v0, w0,
    x0, y0, z0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0;
  output a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, p0, q0, r0, s0, t0, u0, v0,
    w0, x0, y0, z0;
  wire n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n111, n112, n114, n116, n118, n119, n120, n121,
    n122, n124, n126, n127, n128, n129, n130, n131, n133, n134, n135, n136,
    n137, n138, n139, n142, n143, n144, n145, n148, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n163, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180;
  assign n63 = i & d0;
  assign n64 = o0 & n63;
  assign n65 = i & ~c0;
  assign n66 = j0 & n65;
  assign n67 = ~b0 & n66;
  assign n68 = ~e & b0;
  assign n69 = ~c0 & n68;
  assign n70 = j0 & n69;
  assign n71 = ~j & ~e0;
  assign n72 = ~n70 & n71;
  assign n73 = ~n67 & n72;
  assign n74 = ~n64 & n73;
  assign n75 = ~n0 & n73;
  assign h1 = ~n74 & ~n75;
  assign n77 = c0 & j0;
  assign n78 = ~l0 & ~n77;
  assign n79 = b0 & ~n78;
  assign n80 = ~j0 & ~k0;
  assign n81 = c0 & ~k0;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~e & n82;
  assign n84 = ~e & k;
  assign n85 = ~n83 & ~n84;
  assign n86 = ~b0 & ~n84;
  assign n87 = ~n85 & ~n86;
  assign n88 = o0 & n87;
  assign n89 = ~n0 & ~n79;
  assign n90 = ~n79 & ~n88;
  assign b1 = n89 | n90;
  assign n92 = j0 & k0;
  assign n93 = c0 & ~n92;
  assign n94 = ~e0 & ~g0;
  assign n95 = n93 & n94;
  assign n96 = ~b0 & n94;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~e & o0;
  assign n99 = ~n & n98;
  assign n100 = n97 & n99;
  assign n101 = ~j0 & ~l0;
  assign n102 = ~c0 & ~l0;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~s & ~t;
  assign n105 = u & n104;
  assign n106 = b0 & n105;
  assign n107 = n103 & n106;
  assign n108 = ~n100 & ~n107;
  assign n109 = ~n0 & ~n107;
  assign c1 = ~n108 & ~n109;
  assign n111 = a0 & i0;
  assign n112 = m & b0;
  assign e1 = n111 & n112;
  assign n114 = b & w;
  assign f1 = ~x & n114;
  assign n116 = x & n114;
  assign g1 = ~y & n116;
  assign n118 = b0 & j0;
  assign n119 = n71 & ~n118;
  assign n120 = ~n66 & n119;
  assign n121 = ~n64 & n120;
  assign n122 = ~n0 & n120;
  assign j1 = n121 | n122;
  assign n124 = ~p & ~b1;
  assign p0 = ~q | n124;
  assign n126 = e & ~n94;
  assign n127 = e & b0;
  assign n128 = ~c0 & n127;
  assign n129 = j0 & n128;
  assign n130 = k0 & n127;
  assign n131 = ~n129 & ~n130;
  assign q0 = ~n126 & n131;
  assign n133 = ~c0 & j0;
  assign n134 = b0 & n133;
  assign n135 = i & n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~c & ~n63;
  assign n138 = e & n136;
  assign n139 = ~n137 & ~n138;
  assign x0 = n0 & o0;
  assign r0 = ~n139 | ~x0;
  assign n142 = ~b0 & ~l0;
  assign n143 = b0 & ~n77;
  assign n144 = ~n142 & ~n143;
  assign n145 = ~n78 & n144;
  assign s0 = ~v | ~n145;
  assign t0 = v | ~n145;
  assign n148 = b0 & c0;
  assign v0 = ~l0 & ~n148;
  assign n150 = ~p & r;
  assign n151 = ~f0 & ~n150;
  assign n152 = ~h0 & n151;
  assign n153 = o & ~n152;
  assign n154 = d & ~n153;
  assign n155 = ~a & ~z;
  assign n156 = ~a & o;
  assign n157 = o & z;
  assign n158 = ~n156 & ~n157;
  assign n159 = ~n155 & n158;
  assign n160 = ~m0 & n154;
  assign n161 = n154 & n159;
  assign w0 = n160 | n161;
  assign n163 = l & b0;
  assign y0 = n111 & n163;
  assign n165 = ~e & h;
  assign n166 = b0 & n165;
  assign n167 = n82 & n166;
  assign n168 = ~n0 & n167;
  assign n169 = ~o0 & n167;
  assign n170 = ~n168 & ~n169;
  assign n171 = o0 & ~n94;
  assign n172 = o0 & n82;
  assign n173 = b0 & n172;
  assign n174 = ~n171 & ~n173;
  assign n175 = ~e & f;
  assign n176 = n0 & n175;
  assign n177 = ~n174 & n176;
  assign n178 = g & b0;
  assign n179 = l0 & n178;
  assign n180 = ~n177 & ~n179;
  assign z0 = ~n170 | ~n180;
  assign a1 = ~h1;
  assign d1 = ~c1;
  assign u0 = ~v0;
  assign i1 = a1;
endmodule


