// Benchmark "TOP" written by ABC on Sun Apr 24 20:32:56 2016

module TOP ( clock, 
    PCLK, PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_, Pdxport_3_3_,
    Pdxport_4_4_, Pdxport_5_5_, Pdxport_6_6_, Pdxport_7_7_, Pdxport_8_8_,
    Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_, Paport_0_0_, Paport_1_1_,
    Paport_2_2_, Paport_3_3_, Paport_4_4_, Paport_5_5_, Paport_6_6_,
    Paport_7_7_, Paport_8_8_, Paport_9_9_, Paport_10_10_, Paport_11_11_,
    Preset_0_0_, Pready_0_0_,
    PDN, Pnext_0_0_, Pover_0_0_  );
  input  clock;
  input  PCLK, PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_,
    Pdxport_3_3_, Pdxport_4_4_, Pdxport_5_5_, Pdxport_6_6_, Pdxport_7_7_,
    Pdxport_8_8_, Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_,
    Paport_0_0_, Paport_1_1_, Paport_2_2_, Paport_3_3_, Paport_4_4_,
    Paport_5_5_, Paport_6_6_, Paport_7_7_, Paport_8_8_, Paport_9_9_,
    Paport_10_10_, Paport_11_11_, Preset_0_0_, Pready_0_0_;
  output PDN, Pnext_0_0_, Pover_0_0_;
  reg N_N4054, N_N3745, N_N4119, N_N3826, N_N3818, N_N3345, N_N3924,
    N_N3815, N_N3691, N_N3157, N_N3872, N_N3788, N_N3375, N_N3143, N_N4197,
    N_N3843, N_N3426, N_N4118, N_N3580, N_N3175, N_N3071, N_N3808, N_N3923,
    N_N3250, N_N4221, N_N3069, N_N3464, N_N3535, N_N3871, N_N3248, N_N4180,
    N_N3311, N_N3442, N_N3981, N_N3842, N_N3105, N_N4133, N_N4117, N_N3420,
    N_N3761, N_N3062, N_N4071, N_N4227, N_N3807, N_N4145, N_N3922, N_N3516,
    N_N3489, N_N4030, N_N3540, N_N3513, N_N4083, N_N3841, N_N4018, N_N3971,
    N_N4232, N_N4246, N_N3806, N_N3992, N_N4086, N_N4230, N_N4212,
    Pnext_0_0_, N_N3626, N_N3965, N_N3890, NDN3_11, NDN5_10, N_N3786,
    N_N4171, NDN5_16, N_N3799, N_N3844, N_N3196, N_N4126, N_N3681, N_N3679,
    N_N3340, N_N4116, N_N3810, N_N3235, N_N3283, N_N3716, N_N3701, N_N3921,
    N_N3625, N_N3751, N_N3736, N_N3870, N_N4024, N_N3876, N_N3840, N_N4021,
    N_N3932, NLC1_2, N_N3805, N_N3700, N_N3735, NLak3_2, NLak3_9, N_N3906,
    N_N3388, N_N4057, N_N3011, N_N3346, N_N3677, N_N4165, N_N4080, N_N3373,
    N_N3709, N_N4206, N_N3324, N_N3575, N_N4159, NAK5_2, N_N3916, N_N3743,
    N_N4242, N_N3312, N_N3733, N_N3774, N_N4214, N_N3294, N_N3796, N_N3574,
    N_N3791, N_N3480, N_N4243, N_N3940, N_N3509, N_N4015, N_N2989, N_N3919,
    N_N3578, N_N3529, N_N4222, N_N3910, N_N3868, N_N3947, N_N4181, N_N3793,
    N_N3822, N_N3813, N_N4114, N_N4134, N_N3866, N_N4218, N_N3939, N_N3776,
    N_N3387, N_N4194, N_N3821, N_N3882, N_N4167, N_N3800, N_N4237, N_N3417,
    N_N3918, N_N4158, N_N3630, N_N3344, N_N4072, N_N3274, N_N3473, N_N4205,
    N_N4111, N_N3680, N_N3838, N_N3262, N_N4099, N_N3607, N_N3323, N_N3612,
    N_N4079, PDN, N_N3457, N_N3445, N_N3794, N_N3663, N_N3715, N_N4039,
    N_N3280, N_N4239, N_N3988, N_N3433, N_N4075, N_N3468, N_N4045, N_N3482,
    N_N3832, N_N3304, N_N3750, N_N3634, N_N3293, N_N3659, N_N4252, N_N3912,
    N_N3862, N_N3221, N_N3875, N_N3949, N_N3908, N_N3711, N_N3931, N_N3469,
    N_N3436, N_N3974, N_N3905, N_N3741, N_N3369, N_N3164, N_N3500, N_N3996,
    N_N3356, N_N4093, Pover_0_0_, N_N4224, N_N4027, NDN1_4, N_N3384,
    N_N4036, N_N3968, N_N4183, NGFDN_3, N_N4090, N_N4004, N_N3205, N_N4136,
    N_N3303, N_N3533, N_N3336, N_N3961, N_N3331, N_N3203, N_N4236, N_N3884,
    N_N3367, N_N4140, NDN2_2, N_N4106, N_N3100, N_N4193, N_N3470, N_N3424,
    N_N3959, N_N3393, N_N4042, N_N3188, N_N4095, N_N3957, N_N3517, N_N4047,
    N_N3081, N_N3541, N_N4177, NDN3_3, N_N4176, N_N3585, NDN3_8, N_N4209,
    N_N3824, N_N4208, N_N4120, N_N3708, N_N4220, N_N3999, N_N4223, N_N3179,
    N_N4179, N_N3475, N_N4132, N_N4182, N_N3797, N_N3214, N_N4070, N_N4135,
    NLD3_9, NDN5_2, NDN5_3, N_N3778, NDN5_4, N_N3212, NDN5_5, NDN5_6,
    NDN5_7, NDN5_8, N_N4073, NDN5_9, NEN5_9, N_N3684, N_N4056, N_N3713,
    N_N3829, N_N4060, NSr3_2, NSr5_2, NSr5_3, N_N3462, N_N3460, NSr5_4,
    NSr3_9, NSr5_5, NSr5_7, NSr5_8, N_N3998;
  wire n947, n948, n949, n950, n951, n953, n954, n955, n956, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967_1, n968, n969, n970,
    n971, n972_1, n973, n974, n976, n977_1, n978, n979, n980, n981, n982_1,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992_1, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002_1, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022_1, n1023,
    n1024, n1025, n1026, n1027_1, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037_1, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1057_1, n1058, n1060, n1062, n1063, n1064, n1065, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077_1,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087_1,
    n1088, n1089, n1090, n1091, n1092_1, n1093, n1094, n1095, n1096,
    n1097_1, n1098, n1101, n1102, n1103, n1104, n1105, n1106, n1107_1,
    n1108, n1109, n1110, n1111, n1112_1, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122_1, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132_1, n1133, n1134, n1135, n1136,
    n1137_1, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146_1, n1147, n1148, n1149, n1150, n1151_1, n1152, n1153, n1154,
    n1155, n1156_1, n1157, n1158, n1159, n1160, n1161_1, n1162, n1163,
    n1164, n1165, n1166_1, n1167, n1168, n1169, n1170, n1171_1, n1172,
    n1173, n1174, n1175, n1176_1, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231_1, n1232,
    n1233, n1234, n1235, n1236_1, n1237, n1239, n1240, n1241_1, n1242,
    n1244, n1245, n1246_1, n1247, n1248, n1249, n1250, n1251_1, n1252,
    n1253, n1254, n1255, n1256_1, n1257, n1258, n1259, n1260, n1261_1,
    n1262, n1263, n1264, n1265, n1266_1, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1278, n1279, n1280, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301_1, n1302, n1303, n1304,
    n1305, n1306_1, n1307, n1308, n1309, n1310, n1311_1, n1312, n1313,
    n1314, n1315, n1316_1, n1317, n1318, n1319, n1320, n1321_1, n1322,
    n1323, n1324, n1325, n1326_1, n1327, n1328, n1329, n1330, n1331_1,
    n1332, n1333, n1334, n1335, n1336_1, n1337, n1338, n1339, n1340,
    n1341_1, n1342, n1343, n1344, n1345, n1346_1, n1347, n1348, n1349,
    n1350, n1351_1, n1352, n1353, n1354, n1355, n1356_1, n1357, n1358,
    n1359, n1360, n1361_1, n1362, n1363, n1364, n1365, n1366_1, n1367,
    n1368, n1369, n1370, n1371_1, n1372, n1373, n1374, n1375, n1376_1,
    n1377, n1378, n1379, n1380, n1381_1, n1382, n1383, n1384, n1385,
    n1386_1, n1387, n1388, n1389, n1390, n1391_1, n1392, n1393, n1394,
    n1395, n1396_1, n1397, n1398, n1399, n1400, n1401_1, n1402, n1403,
    n1404, n1405, n1406_1, n1407, n1408, n1409, n1410, n1411_1, n1412,
    n1413, n1414, n1415, n1416_1, n1417, n1418, n1419, n1420, n1421_1,
    n1422, n1423, n1424, n1425, n1426_1, n1427, n1428, n1429, n1430,
    n1431_1, n1432, n1433, n1434, n1435, n1436_1, n1437, n1439, n1440,
    n1441_1, n1442, n1445, n1446_1, n1447, n1448, n1451_1, n1452, n1453,
    n1454, n1455, n1457, n1458, n1459, n1461_1, n1462, n1463, n1464,
    n1466_1, n1467, n1468, n1469, n1472, n1473, n1475, n1476_1, n1477,
    n1479, n1480, n1481_1, n1482, n1483, n1484, n1485, n1486_1, n1487,
    n1489, n1490, n1491_1, n1492, n1493, n1494, n1495, n1496_1, n1497,
    n1498, n1499, n1500, n1501_1, n1502, n1503, n1504, n1505, n1506_1,
    n1507, n1508, n1509, n1510, n1511_1, n1512, n1514, n1515, n1516_1,
    n1517, n1520, n1521_1, n1523, n1524, n1525, n1527, n1528, n1529, n1530,
    n1531_1, n1532, n1534, n1535, n1536_1, n1537, n1538, n1539, n1540,
    n1541_1, n1542, n1543, n1544, n1545, n1546_1, n1547, n1548, n1549,
    n1550, n1551_1, n1552, n1553, n1554, n1555, n1556_1, n1557, n1558,
    n1559, n1561_1, n1562, n1563, n1564, n1567, n1568, n1570, n1571_1,
    n1572, n1573, n1574, n1576_1, n1577, n1579, n1580, n1581_1, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1607, n1608, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1631, n1632, n1633, n1634, n1636, n1637,
    n1638, n1639, n1640, n1641, n1643, n1644, n1646, n1647, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1676, n1677, n1679, n1680, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1709, n1710, n1711, n1712, n1713, n1714,
    n1716, n1717, n1719, n1720, n1721, n1722, n1723, n1724, n1726, n1727,
    n1728, n1729, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1757, n1758, n1760, n1761,
    n1762, n1763, n1764, n1765, n1767, n1768, n1769, n1770, n1773, n1774,
    n1775, n1776, n1777, n1778, n1781, n1782, n1783, n1785, n1786, n1787,
    n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1797, n1798, n1799,
    n1800, n1802, n1804, n1807, n1808, n1809, n1810, n1811, n1812, n1815,
    n1816, n1817, n1819, n1820, n1821, n1822, n1825, n1826, n1827, n1828,
    n1829, n1830, n1833, n1834, n1835, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1850, n1851, n1852,
    n1853, n1854, n1856, n1857, n1858, n1859, n1862, n1863, n1864, n1865,
    n1866, n1867, n1870, n1871, n1872, n1874, n1875, n1877, n1878, n1879,
    n1880, n1881, n1884, n1885, n1886, n1888, n1889, n1891, n1892, n1895,
    n1896, n1898, n1899, n1903, n1904, n1906, n1907, n1909, n1910, n1912,
    n1913, n1914, n1915, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1964,
    n1965, n1967, n1969, n1970, n1973, n1975, n1976, n1977, n1978, n1980,
    n1981, n1985, n1986, n1987, n1988, n1989, n1990, n1992, n1993, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2014, n2015, n2017, n2018, n2019, n2020,
    n2021, n2022, n2024, n2025, n2028, n2029, n2031, n2032, n2033, n2034,
    n2035, n2036, n2038, n2039, n2040, n2043, n2044, n2045, n2046, n2048,
    n2049, n2051, n2052, n2053, n2054, n2055, n2056, n2058, n2059, n2060,
    n2061, n2062, n2063, n2065, n2066, n2068, n2069, n2070, n2071, n2073,
    n2074, n2075, n2076, n2077, n2078, n2080, n2081, n2083, n2085, n2086,
    n2087, n2088, n2090, n2092, n2093, n2094, n2095, n2096, n2097, n2100,
    n2101, n2103, n2104, n2105, n2106, n2108, n2109, n2110, n2111, n2112,
    n2113, n2116, n2117, n2120, n2121, n2122, n2123, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2161,
    n2162, n2163, n2164, n2166, n2167, n2169, n2170, n2172, n2173, n2175,
    n2176, n2177, n2178, n2179, n2180, n2182, n2183, n2185, n2186, n2188,
    n2189, n2190, n2191, n2193, n2194, n2197, n2198, n2199, n2200, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2229, n2230, n2232, n2233, n2236,
    n2237, n2239, n2240, n2241, n2243, n2244, n2246, n2247, n2249, n2250,
    n2252, n2255, n2256, n2257, n2258, n2260, n2261, n2263, n2264, n2266,
    n2267, n2268, n2270, n2271, n2272, n2273, n2274, n2275, n2277, n2279,
    n2280, n2283, n2284, n2286, n2287, n2289, n2290, n2292, n2293, n2296,
    n2297, n2298, n2299, n2301, n2302, n2304, n2305, n2307, n2308, n2311,
    n2312, n2314, n2315, n2317, n2318, n2320, n2321, n2323, n2324, n2327,
    n2328, n2330, n2331, n2333, n2334, n2335, n2336, n2338, n2339, n2340,
    n2341, n2342, n2343, n2345, n2346, n2348, n2349, n2351, n2352, n2354,
    n2355, n2356, n2357, n2358, n2359, n2361, n2362, n2364, n2365, n2367,
    n2368, n2371, n2372, n2374, n2375, n2376, n2377, n2378, n2379, n2383,
    n2384, n2385, n2386, n2387, n2388, n2390, n2391, n2393, n2394, n2395,
    n2396, n2398, n2399, n2400, n2401, n2402, n2403, n2406, n2407, n2408,
    n2409, n2412, n2413, n2414, n2416, n2417, n2418, n2419, n2421, n2422,
    n2423, n2424, n2425, n2426, n2430, n2431, n2432, n2433, n2434, n2435,
    n2437, n2438, n2440, n2441, n2442, n2443, n2446, n2447, n2448, n2449,
    n2451, n2452, n2454, n2455, n2456, n2457, n2459, n2460, n2463, n2464,
    n2466, n2467, n2468, n2469, n2470, n2471, n2474, n2475, n2477, n2478,
    n2480, n2481, n2483, n2484, n2486, n2487, n2488, n2489, n2491, n2494,
    n2495, n2497, n2498, n2500, n2501, n2502, n2503, n2505, n2506, n2508,
    n2509, n2512, n2513, n2515, n2516, n2518, n2519, n2520, n2521, n2523,
    n2524, n2527, n2528, n2530, n2531, n2534, n2535, n2536, n2537, n2539,
    n2541, n2542, n2543, n2544, n2546, n2547, n2549, n2551, n2552, n2553,
    n2554, n2556, n2557, n2559, n2560, n2561, n2562, n2564, n2565, n2568,
    n2569, n2571, n2574, n2575, n2577, n2578, n2580, n2581, n2583, n2584,
    n2587, n2588, n2590, n2591, n2593, n2594, n2599, n2600, n2603, n2604,
    n2607, n2612, n2614, n2616, n2617, n2619, n2620, n2622, n2623, n2625,
    n2626, n2628, n2629, n2630, n2631, n2633, n2635, n2636, n2638, n2639,
    n2641, n2644, n2645, n2647, n2648, n2650, n2651, n2653, n2654, n2656,
    n2657, n2659, n2660, n64_1, n69, n74_1, n79, n84_1, n89_1, n94_1, n99,
    n104_1, n109, n114_1, n119_1, n124_1, n129, n134, n139_1, n144_1,
    n149_1, n154_1, n159_1, n164_1, n169_1, n174, n179_1, n184_1, n189_1,
    n194_1, n199_1, n204_1, n209_1, n214_1, n219, n224_1, n229_1, n234_1,
    n239_1, n244_1, n249_1, n254, n259_1, n264_1, n269_1, n274, n279_1,
    n284, n289, n294, n299_1, n304_1, n309, n314, n319_1, n324_1, n329,
    n334, n339_1, n344_1, n349_1, n354, n359, n364, n369_1, n374_1, n378_1,
    n383_1, n388_1, n393_1, n398_1, n403, n408_1, n413_1, n418_1, n423,
    n428_1, n433_1, n438, n443, n448_1, n453, n458_1, n463_1, n468, n473_1,
    n478_1, n483, n488, n493_1, n498, n503, n508_1, n513, n518_1, n523,
    n528_1, n533_1, n538, n543_1, n548, n553_1, n558, n563_1, n568_1,
    n573_1, n578, n583_1, n588, n593, n598, n603, n608, n613_1, n618_1,
    n623_1, n628, n633, n638_1, n643, n648_1, n653_1, n658, n663, n668_1,
    n673, n678_1, n683, n688_1, n693, n698_1, n703_1, n708, n713_1, n718,
    n723, n728, n733, n738, n743, n748_1, n753, n758, n763, n768, n773_1,
    n778_1, n783_1, n788, n793_1, n798, n803_1, n808_1, n813, n818_1,
    n823_1, n828_1, n833, n838_1, n843_1, n848_1, n853, n858_1, n863_1,
    n868, n873_1, n878_1, n883, n888_1, n893, n898, n903, n908, n913,
    n918_1, n923, n928, n933, n937, n942, n947_1, n952, n957_1, n962_1,
    n967, n972, n977, n982, n987_1, n992, n997_1, n1002, n1007_1, n1012_1,
    n1017_1, n1022, n1027, n1032_1, n1037, n1042_1, n1047_1, n1052_1,
    n1057, n1062_1, n1067_1, n1072_1, n1077, n1082_1, n1087, n1092, n1097,
    n1102_1, n1107, n1112, n1117_1, n1122, n1127_1, n1132, n1137, n1141_1,
    n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181_1, n1186_1,
    n1191_1, n1196_1, n1201_1, n1206_1, n1211_1, n1216_1, n1221_1, n1226_1,
    n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271_1,
    n1276_1, n1281, n1286_1, n1291_1, n1296_1, n1301, n1306, n1311, n1316,
    n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366,
    n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416,
    n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466,
    n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1511, n1516,
    n1521, n1526, n1531, n1536, n1541, n1546, n1551, n1556, n1561, n1566,
    n1571, n1576, n1581;
  assign n947 = ~NDN3_3 & ~NSr3_2;
  assign n948 = ~PRESET & ~n947;
  assign n949 = N_N4054 & n948;
  assign n950 = ~PRESET & n947;
  assign n951 = Paport_7_7_ & n950;
  assign n64_1 = n949 | n951;
  assign n953 = ~NLC1_2 & ~PDN;
  assign n954 = Preset_0_0_ & n953;
  assign n955 = ~NDN2_2 & n954;
  assign n956 = ~N_N3745 & ~n955;
  assign n69 = ~PRESET & ~n956;
  assign n958 = Preset_0_0_ & ~NLC1_2;
  assign n959 = NLC1_2 & ~N_N3998;
  assign n960 = ~n958 & ~n959;
  assign n961 = PDN & ~NDN1_4;
  assign n962 = ~PRESET & n961;
  assign n963 = n960 & n962;
  assign n964 = NDN3_3 & ~NDN3_8;
  assign n965 = ~PRESET & ~NLD3_9;
  assign n966 = ~n964 & n965;
  assign n967_1 = ~n961 & n966;
  assign n968 = ~n963 & ~n967_1;
  assign n969 = N_N4119 & ~n968;
  assign n970 = ~PRESET & NLD3_9;
  assign n971 = N_N3535 & n970;
  assign n972_1 = ~PRESET & n964;
  assign n973 = N_N3580 & n972_1;
  assign n974 = ~n971 & ~n973;
  assign n74_1 = n969 | ~n974;
  assign n976 = ~NDN5_10 & ~NSr5_7;
  assign n977_1 = ~PRESET & n976;
  assign n978 = N_N4183 & n976;
  assign n979 = ~NDN5_9 & NEN5_9;
  assign n980 = N_N3826 & n979;
  assign n981 = ~n978 & ~n980;
  assign n982_1 = N_N3679 & n976;
  assign n983 = N_N4021 & n979;
  assign n984 = ~n982_1 & ~n983;
  assign n985 = N_N3799 & n976;
  assign n986 = N_N4024 & n979;
  assign n987 = ~n985 & ~n986;
  assign n988 = N_N3626 & n976;
  assign n989 = N_N3625 & n979;
  assign n990 = ~n988 & ~n989;
  assign n991 = N_N3968 & n976;
  assign n992_1 = N_N3959 & n979;
  assign n993 = ~n991 & ~n992_1;
  assign n994 = n990 & n993;
  assign n995 = n987 & n994;
  assign n996 = N_N3205 & n976;
  assign n997 = N_N3957 & n979;
  assign n998 = ~n996 & ~n997;
  assign n999 = n995 & n998;
  assign n1000 = n984 & n999;
  assign n1001 = N_N3203 & n976;
  assign n1002_1 = N_N3081 & n979;
  assign n1003 = ~n1001 & ~n1002_1;
  assign n1004 = n1000 & n1003;
  assign n1005 = ~n1000 & ~n1003;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n981 & n1006;
  assign n1008 = n981 & ~n1006;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = N_N3890 & n976;
  assign n1011 = N_N3509 & n979;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n984 & ~n999;
  assign n1014 = ~n1000 & ~n1013;
  assign n1015 = ~n1012 & n1014;
  assign n1016 = n1012 & ~n1014;
  assign n1017 = N_N4224 & n976;
  assign n1018 = N_N3829 & n979;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = N_N4086 & n976;
  assign n1021 = N_N3480 & n979;
  assign n1022_1 = ~n1020 & ~n1021;
  assign n1023 = ~n987 & ~n994;
  assign n1024 = ~n995 & ~n1023;
  assign n1025 = ~n1022_1 & n1024;
  assign n1026 = n1022_1 & ~n1024;
  assign n1027_1 = N_N3500 & n976;
  assign n1028 = N_N3684 & n979;
  assign n1029 = ~n1027_1 & ~n1028;
  assign n1030 = ~n990 & ~n993;
  assign n1031 = ~n994 & ~n1030;
  assign n1032 = ~n1029 & n1031;
  assign n1033 = ~n993 & n1029;
  assign n1034 = N_N3971 & n976;
  assign n1035 = N_N3796 & n979;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037_1 = ~n990 & ~n1036;
  assign n1038 = ~n1033 & n1037_1;
  assign n1039 = ~n1032 & ~n1038;
  assign n1040 = ~n1026 & ~n1039;
  assign n1041 = ~n1025 & ~n1040;
  assign n1042 = ~n1019 & ~n1041;
  assign n1043 = n1019 & n1041;
  assign n1044 = ~n995 & ~n998;
  assign n1045 = ~n999 & ~n1044;
  assign n1046 = ~n1043 & n1045;
  assign n1047 = ~n1042 & ~n1046;
  assign n1048 = ~n1016 & ~n1047;
  assign n1049 = ~n1015 & ~n1048;
  assign n1050 = n1009 & n1049;
  assign n1051 = ~n1009 & ~n1049;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n977_1 & ~n1052;
  assign n1054 = ~PRESET & ~n976;
  assign n1055 = N_N3826 & n1054;
  assign n79 = n1053 | n1055;
  assign n1057_1 = N_N3818 & n948;
  assign n1058 = Paport_9_9_ & n950;
  assign n84_1 = n1057_1 | n1058;
  assign n1060 = ~PRESET & ~n955;
  assign n89_1 = N_N3345 & n1060;
  assign n1062 = N_N3924 & ~n968;
  assign n1063 = N_N3981 & n970;
  assign n1064 = N_N3250 & n972_1;
  assign n1065 = ~n1063 & ~n1064;
  assign n94_1 = n1062 | ~n1065;
  assign n1067 = N_N3844 & n976;
  assign n1068 = N_N3529 & n979;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = N_N3701 & n976;
  assign n1071 = N_N3700 & n979;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = n1004 & n1072;
  assign n1074 = ~n1004 & ~n1072;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = ~n1069 & n1075;
  assign n1077_1 = n1069 & ~n1075;
  assign n1078 = ~n1008 & ~n1049;
  assign n1079 = ~n1007 & ~n1078;
  assign n1080 = ~n1077_1 & ~n1079;
  assign n1081 = ~n1076 & ~n1080;
  assign n1082 = N_N4136 & n976;
  assign n1083 = N_N3815 & n979;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = N_N3100 & n976;
  assign n1086 = N_N3585 & n979;
  assign n1087_1 = ~n1085 & ~n1086;
  assign n1088 = n1073 & n1087_1;
  assign n1089 = ~n1073 & ~n1087_1;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n1084 & ~n1090;
  assign n1092_1 = ~n1084 & n1090;
  assign n1093 = ~n1091 & ~n1092_1;
  assign n1094 = ~n1081 & ~n1093;
  assign n1095 = n1081 & n1093;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097_1 = n977_1 & ~n1096;
  assign n1098 = N_N3815 & n1054;
  assign n99 = n1097_1 | n1098;
  assign n104_1 = N_N3691 & n1060;
  assign n1101 = ~NDN5_5 & ~NSr5_5;
  assign n1102 = ~PRESET & n1101;
  assign n1103 = ~N_N3838 & N_N3999;
  assign n1104 = NDN3_8 & NSr3_9;
  assign n1105 = ~NLak3_9 & n1104;
  assign n1106 = NSr5_2 & n1105;
  assign n1107_1 = ~NSr5_4 & NSr5_5;
  assign n1108 = ~n1106 & ~n1107_1;
  assign n1109 = N_N4194 & ~n1108;
  assign n1110 = ~NSr5_7 & NSr5_8;
  assign n1111 = N_N4045 & n1110;
  assign n1112_1 = ~NSr5_2 & NSr5_3;
  assign n1113 = N_N4177 & n1112_1;
  assign n1114 = ~NSr5_3 & NSr5_4;
  assign n1115 = N_N4176 & n1114;
  assign n1116 = ~NSr5_5 & NSr5_7;
  assign n1117 = N_N3457 & n1116;
  assign n1118 = ~n1115 & ~n1117;
  assign n1119 = ~n1113 & n1118;
  assign n1120 = ~n1111 & n1119;
  assign n1121 = ~n1109 & n1120;
  assign n1122_1 = ~N_N3999 & n1121;
  assign n1123 = N_N4070 & ~n1108;
  assign n1124 = N_N3808 & n1112_1;
  assign n1125 = N_N3806 & n1116;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n1123 & n1126;
  assign n1128 = N_N3807 & n1114;
  assign n1129 = N_N3805 & n1110;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = n1127 & n1130;
  assign n1132_1 = N_N4179 & ~n1108;
  assign n1133 = N_N3872 & n1112_1;
  assign n1134 = N_N3870 & n1110;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = N_N4030 & n1116;
  assign n1137_1 = N_N3871 & n1114;
  assign n1138 = ~n1136 & ~n1137_1;
  assign n1139 = n1135 & n1138;
  assign n1140 = ~n1132_1 & n1139;
  assign n1141 = N_N4206 & ~n1108;
  assign n1142 = N_N3813 & n1112_1;
  assign n1143 = N_N3188 & n1110;
  assign n1144 = N_N4239 & n1114;
  assign n1145 = N_N3436 & n1116;
  assign n1146_1 = ~n1144 & ~n1145;
  assign n1147 = ~n1143 & n1146_1;
  assign n1148 = ~n1142 & n1147;
  assign n1149 = ~n1141 & n1148;
  assign n1150 = n1140 & n1149;
  assign n1151_1 = n1131 & n1150;
  assign n1152 = N_N4220 & ~n1108;
  assign n1153 = N_N3922 & n1116;
  assign n1154 = N_N3921 & n1110;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156_1 = N_N3924 & n1112_1;
  assign n1157 = N_N3923 & n1114;
  assign n1158 = ~n1156_1 & ~n1157;
  assign n1159 = n1155 & n1158;
  assign n1160 = ~n1152 & n1159;
  assign n1161_1 = N_N3906 & ~n1108;
  assign n1162 = N_N3939 & n1114;
  assign n1163 = N_N3940 & n1112_1;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = N_N3304 & n1116;
  assign n1166_1 = N_N3303 & n1110;
  assign n1167 = ~n1165 & ~n1166_1;
  assign n1168 = n1164 & n1167;
  assign n1169 = ~n1161_1 & n1168;
  assign n1170 = N_N4120 & ~n1108;
  assign n1171_1 = N_N4116 & n1110;
  assign n1172 = N_N4117 & n1116;
  assign n1173 = ~n1171_1 & ~n1172;
  assign n1174 = N_N4119 & n1112_1;
  assign n1175 = N_N4118 & n1114;
  assign n1176_1 = ~n1174 & ~n1175;
  assign n1177 = n1173 & n1176_1;
  assign n1178 = ~n1170 & n1177;
  assign n1179 = n1169 & n1178;
  assign n1180 = N_N4237 & ~n1108;
  assign n1181 = N_N3433 & n1116;
  assign n1182 = N_N4208 & n1114;
  assign n1183 = N_N3659 & n1110;
  assign n1184 = N_N4209 & n1112_1;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = ~n1182 & n1185;
  assign n1187 = ~n1181 & n1186;
  assign n1188 = ~n1180 & n1187;
  assign n1189 = N_N4242 & ~n1108;
  assign n1190 = N_N4047 & n1110;
  assign n1191 = N_N3800 & n1112_1;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = N_N3164 & n1116;
  assign n1194 = N_N4252 & n1114;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1192 & n1195;
  assign n1197 = ~n1189 & n1196;
  assign n1198 = n1188 & n1197;
  assign n1199 = n1179 & n1198;
  assign n1200 = n1160 & n1199;
  assign n1201 = N_N4057 & ~n1108;
  assign n1202 = N_N3367 & n1110;
  assign n1203 = N_N3918 & n1114;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = N_N3221 & n1116;
  assign n1206 = N_N3919 & n1112_1;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = n1204 & n1207;
  assign n1209 = ~n1201 & n1208;
  assign n1210 = N_N4165 & ~n1108;
  assign n1211 = N_N3868 & n1112_1;
  assign n1212 = N_N4099 & n1114;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = N_N3711 & n1116;
  assign n1215 = N_N3424 & n1110;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = n1213 & n1216;
  assign n1218 = ~n1210 & n1217;
  assign n1219 = N_N4132 & ~n1108;
  assign n1220 = N_N3842 & n1114;
  assign n1221 = N_N3840 & n1110;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = N_N3841 & n1116;
  assign n1224 = N_N3843 & n1112_1;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n1222 & n1225;
  assign n1227 = ~n1219 & n1226;
  assign n1228 = n1218 & n1227;
  assign n1229 = n1209 & n1228;
  assign n1230 = n1200 & n1229;
  assign n1231_1 = n1151_1 & n1230;
  assign n1232 = n1122_1 & n1231_1;
  assign n1233 = ~n1103 & ~n1232;
  assign n1234 = N_N4027 & n1233;
  assign n1235 = n1102 & n1234;
  assign n1236_1 = ~PRESET & ~n1101;
  assign n1237 = N_N3157 & n1236_1;
  assign n109 = n1235 | n1237;
  assign n1239 = N_N3872 & ~n968;
  assign n1240 = N_N3761 & n970;
  assign n1241_1 = N_N3248 & n972_1;
  assign n1242 = ~n1240 & ~n1241_1;
  assign n114_1 = n1239 | ~n1242;
  assign n1244 = N_N4042 & n976;
  assign n1245 = N_N3824 & n979;
  assign n1246_1 = ~n1244 & ~n1245;
  assign n1247 = N_N3736 & n976;
  assign n1248 = N_N3735 & n979;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = n1088 & n1249;
  assign n1251_1 = n1246_1 & n1250;
  assign n1252 = ~n1246_1 & ~n1250;
  assign n1253 = ~n1251_1 & ~n1252;
  assign n1254 = N_N4140 & n976;
  assign n1255 = N_N3788 & n979;
  assign n1256_1 = ~n1254 & ~n1255;
  assign n1257 = ~n1088 & ~n1249;
  assign n1258 = ~n1250 & ~n1257;
  assign n1259 = ~n1081 & ~n1091;
  assign n1260 = ~n1092_1 & ~n1259;
  assign n1261_1 = ~n1258 & n1260;
  assign n1262 = n1258 & ~n1260;
  assign n1263 = N_N3810 & n976;
  assign n1264 = N_N3947 & n979;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266_1 = ~n1262 & n1265;
  assign n1267 = ~n1261_1 & ~n1266_1;
  assign n1268 = n1256_1 & ~n1267;
  assign n1269 = ~n1256_1 & n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1253 & n1270;
  assign n1272 = n1253 & ~n1270;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = n977_1 & ~n1273;
  assign n1275 = N_N3788 & n1054;
  assign n119_1 = n1274 | n1275;
  assign n124_1 = N_N3375 & n1060;
  assign n1278 = N_N3996 & n1233;
  assign n1279 = n1102 & n1278;
  assign n1280 = N_N3143 & n1236_1;
  assign n129 = n1279 | n1280;
  assign n1282 = N_N4214 & N_N3462;
  assign n1283 = ~N_N3575 & n1282;
  assign n1284 = ~n1112_1 & ~n1116;
  assign n1285 = ~n1110 & n1284;
  assign n1286 = ~n1114 & n1285;
  assign n1287 = n1108 & n1286;
  assign n1288 = N_N3460 & n1233;
  assign n1289 = ~n1287 & n1288;
  assign n1290 = ~N_N4214 & n1289;
  assign n1291 = ~n1283 & ~n1290;
  assign n1292 = ~PRESET & n1291;
  assign n1293 = N_N4197 & n1292;
  assign n1294 = ~PRESET & n1283;
  assign n1295 = N_N3470 & ~n1108;
  assign n1296 = N_N3473 & n1116;
  assign n1297 = N_N3469 & n1112_1;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = N_N4194 & n1110;
  assign n1300 = N_N3468 & n1114;
  assign n1301_1 = ~n1299 & ~n1300;
  assign n1302 = n1298 & n1301_1;
  assign n1303 = ~n1295 & n1302;
  assign n1304 = N_N3500 & ~n1108;
  assign n1305 = N_N4120 & n1110;
  assign n1306_1 = N_N3708 & n1112_1;
  assign n1307 = ~n1305 & ~n1306_1;
  assign n1308 = N_N3175 & n1116;
  assign n1309 = N_N2989 & n1114;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311_1 = n1307 & n1310;
  assign n1312 = ~n1304 & n1311_1;
  assign n1313 = N_N3971 & ~n1108;
  assign n1314 = N_N3388 & n1112_1;
  assign n1315 = N_N3906 & n1110;
  assign n1316_1 = ~n1314 & ~n1315;
  assign n1317 = ~n1313 & n1316_1;
  assign n1318 = N_N3745 & n1114;
  assign n1319 = N_N3387 & n1116;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321_1 = n1317 & n1320;
  assign n1322 = N_N3965 & ~n1321_1;
  assign n1323 = ~n1312 & n1322;
  assign n1324 = n1312 & ~n1322;
  assign n1325 = N_N4027 & ~n1324;
  assign n1326_1 = ~n1323 & ~n1325;
  assign n1327 = N_N3992 & ~n1326_1;
  assign n1328 = ~N_N3992 & n1326_1;
  assign n1329 = N_N4086 & ~n1108;
  assign n1330 = N_N3345 & n1114;
  assign n1331_1 = N_N3344 & n1116;
  assign n1332 = N_N3346 & n1112_1;
  assign n1333 = N_N4057 & n1110;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1331_1 & n1334;
  assign n1336_1 = ~n1330 & n1335;
  assign n1337 = ~n1329 & n1336_1;
  assign n1338 = ~n1328 & ~n1337;
  assign n1339 = ~n1327 & ~n1338;
  assign n1340 = N_N3996 & ~n1339;
  assign n1341_1 = ~N_N3996 & n1339;
  assign n1342 = N_N4224 & ~n1108;
  assign n1343 = N_N4222 & n1114;
  assign n1344 = N_N4223 & n1112_1;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346_1 = N_N4220 & n1110;
  assign n1347 = N_N4221 & n1116;
  assign n1348 = ~n1346_1 & ~n1347;
  assign n1349 = n1345 & n1348;
  assign n1350 = ~n1342 & n1349;
  assign n1351_1 = ~n1341_1 & ~n1350;
  assign n1352 = ~n1340 & ~n1351_1;
  assign n1353 = N_N4018 & ~n1352;
  assign n1354 = ~N_N4018 & n1352;
  assign n1355 = N_N3890 & ~n1108;
  assign n1356_1 = N_N3323 & n1116;
  assign n1357 = N_N4165 & n1110;
  assign n1358 = ~n1356_1 & ~n1357;
  assign n1359 = N_N3691 & n1114;
  assign n1360 = N_N3324 & n1112_1;
  assign n1361_1 = ~n1359 & ~n1360;
  assign n1362 = n1358 & n1361_1;
  assign n1363 = ~n1355 & n1362;
  assign n1364 = ~n1354 & ~n1363;
  assign n1365 = ~n1353 & ~n1364;
  assign n1366_1 = N_N3974 & ~n1365;
  assign n1367 = ~N_N3974 & n1365;
  assign n1368 = N_N4183 & ~n1108;
  assign n1369 = N_N4180 & n1116;
  assign n1370 = N_N4181 & n1114;
  assign n1371_1 = ~n1369 & ~n1370;
  assign n1372 = N_N4179 & n1110;
  assign n1373 = N_N4182 & n1112_1;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = n1371_1 & n1374;
  assign n1376_1 = ~n1368 & n1375;
  assign n1377 = ~n1367 & ~n1376_1;
  assign n1378 = ~n1366_1 & ~n1377;
  assign n1379 = N_N4083 & ~n1378;
  assign n1380 = ~N_N4083 & n1378;
  assign n1381_1 = N_N3844 & ~n1108;
  assign n1382 = N_N3312 & n1112_1;
  assign n1383 = N_N3375 & n1114;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = N_N4206 & n1110;
  assign n1386_1 = N_N3988 & n1116;
  assign n1387 = ~n1385 & ~n1386_1;
  assign n1388 = n1384 & n1387;
  assign n1389 = ~n1381_1 & n1388;
  assign n1390 = ~n1380 & ~n1389;
  assign n1391_1 = ~n1379 & ~n1390;
  assign n1392 = N_N3949 & ~n1391_1;
  assign n1393 = ~N_N3949 & n1391_1;
  assign n1394 = N_N4136 & ~n1108;
  assign n1395 = N_N4135 & n1112_1;
  assign n1396_1 = N_N4132 & n1110;
  assign n1397 = ~n1395 & ~n1396_1;
  assign n1398 = N_N4133 & n1116;
  assign n1399 = N_N4134 & n1114;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401_1 = n1397 & n1400;
  assign n1402 = ~n1394 & n1401_1;
  assign n1403 = ~n1393 & ~n1402;
  assign n1404 = ~n1392 & ~n1403;
  assign n1405 = N_N4145 & ~n1404;
  assign n1406_1 = ~N_N4145 & n1404;
  assign n1407 = N_N3810 & ~n1108;
  assign n1408 = N_N3426 & n1114;
  assign n1409 = N_N3293 & n1116;
  assign n1410 = N_N3294 & n1112_1;
  assign n1411_1 = N_N4242 & n1110;
  assign n1412 = ~n1410 & ~n1411_1;
  assign n1413 = ~n1409 & n1412;
  assign n1414 = ~n1408 & n1413;
  assign n1415 = ~n1407 & n1414;
  assign n1416_1 = ~n1406_1 & ~n1415;
  assign n1417 = ~n1405 & ~n1416_1;
  assign n1418 = N_N3912 & ~n1417;
  assign n1419 = ~N_N3912 & n1417;
  assign n1420 = N_N4140 & ~n1108;
  assign n1421_1 = N_N4070 & n1110;
  assign n1422 = N_N4072 & n1114;
  assign n1423 = N_N4073 & n1112_1;
  assign n1424 = N_N4071 & n1116;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426_1 = ~n1422 & n1425;
  assign n1427 = ~n1421_1 & n1426_1;
  assign n1428 = ~n1420 & n1427;
  assign n1429 = ~n1419 & ~n1428;
  assign n1430 = ~n1418 & ~n1429;
  assign n1431_1 = N_N4197 & ~n1430;
  assign n1432 = ~N_N4197 & n1430;
  assign n1433 = ~n1431_1 & ~n1432;
  assign n1434 = n1303 & ~n1433;
  assign n1435 = ~n1303 & n1433;
  assign n1436_1 = ~n1434 & ~n1435;
  assign n1437 = n1294 & n1436_1;
  assign n134 = n1293 | n1437;
  assign n1439 = N_N3843 & ~n968;
  assign n1440 = N_N3105 & n972_1;
  assign n1441_1 = N_N3489 & n970;
  assign n1442 = ~n1440 & ~n1441_1;
  assign n139_1 = n1439 | ~n1442;
  assign n144_1 = N_N3426 & n1060;
  assign n1445 = N_N4118 & ~n968;
  assign n1446_1 = N_N4232 & n972_1;
  assign n1447 = N_N3179 & n970;
  assign n1448 = ~n1446_1 & ~n1447;
  assign n149_1 = n1445 | ~n1448;
  assign n154_1 = N_N3580 & n948;
  assign n1451_1 = ~NDN5_2 & ~NSr5_2;
  assign n1452 = ~PRESET & n1451_1;
  assign n1453 = n1234 & n1452;
  assign n1454 = ~PRESET & ~n1451_1;
  assign n1455 = N_N3175 & n1454;
  assign n159_1 = n1453 | n1455;
  assign n1457 = N_N3071 & n1236_1;
  assign n1458 = N_N3974 & n1233;
  assign n1459 = n1102 & n1458;
  assign n164_1 = n1457 | n1459;
  assign n1461_1 = N_N3808 & ~n968;
  assign n1462 = N_N3062 & n972_1;
  assign n1463 = N_N3513 & n970;
  assign n1464 = ~n1462 & ~n1463;
  assign n169_1 = n1461_1 | ~n1464;
  assign n1466_1 = N_N3923 & ~n968;
  assign n1467 = N_N3475 & n970;
  assign n1468 = N_N4230 & n972_1;
  assign n1469 = ~n1467 & ~n1468;
  assign n174 = n1466_1 | ~n1469;
  assign n179_1 = N_N3250 & n948;
  assign n1472 = n1278 & n1452;
  assign n1473 = N_N4221 & n1454;
  assign n184_1 = n1472 | n1473;
  assign n1475 = N_N3949 & n1233;
  assign n1476_1 = n1102 & n1475;
  assign n1477 = N_N3069 & n1236_1;
  assign n189_1 = n1476_1 | n1477;
  assign n1479 = ~PRESET & n979;
  assign n1480 = n1029 & ~n1031;
  assign n1481_1 = ~n1032 & ~n1480;
  assign n1482 = ~n1037_1 & ~n1481_1;
  assign n1483 = n1037_1 & n1481_1;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = n1479 & n1484;
  assign n1486_1 = ~PRESET & ~n979;
  assign n1487 = N_N3464 & n1486_1;
  assign n194_1 = n1485 | n1487;
  assign n1489 = ~NDN5_6 & n1105;
  assign n1490 = ~PRESET & n1489;
  assign n1491_1 = N_N3940 & n1489;
  assign n1492 = N_N3939 & n979;
  assign n1493 = ~n1491_1 & ~n1492;
  assign n1494 = N_N3906 & n1489;
  assign n1495 = N_N3910 & n979;
  assign n1496_1 = ~n1494 & ~n1495;
  assign n1497 = ~n1493 & ~n1496_1;
  assign n1498 = N_N4119 & n1489;
  assign n1499 = N_N4118 & n979;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501_1 = N_N4120 & n1489;
  assign n1502 = N_N3157 & n979;
  assign n1503 = ~n1501_1 & ~n1502;
  assign n1504 = n1500 & n1503;
  assign n1505 = ~n1500 & ~n1503;
  assign n1506_1 = ~n1504 & ~n1505;
  assign n1507 = ~n1497 & n1506_1;
  assign n1508 = n1497 & ~n1506_1;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = n1490 & ~n1509;
  assign n1511_1 = ~PRESET & ~n1489;
  assign n1512 = N_N3535 & n1511_1;
  assign n199_1 = n1510 | n1512;
  assign n1514 = N_N3871 & ~n968;
  assign n1515 = N_N3214 & n970;
  assign n1516_1 = N_N3786 & n972_1;
  assign n1517 = ~n1515 & ~n1516_1;
  assign n204_1 = n1514 | ~n1517;
  assign n209_1 = N_N3248 & n948;
  assign n1520 = N_N4180 & n1454;
  assign n1521_1 = n1452 & n1458;
  assign n214_1 = n1520 | n1521_1;
  assign n1523 = N_N3311 & n1236_1;
  assign n1524 = N_N3912 & n1233;
  assign n1525 = n1102 & n1524;
  assign n219 = n1523 | n1525;
  assign n1527 = ~n1042 & ~n1043;
  assign n1528 = ~n1045 & ~n1527;
  assign n1529 = n1045 & n1527;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531_1 = n1479 & n1530;
  assign n1532 = N_N3442 & n1486_1;
  assign n224_1 = n1531_1 | n1532;
  assign n1534 = N_N4220 & n1489;
  assign n1535 = N_N3143 & n979;
  assign n1536_1 = ~n1534 & ~n1535;
  assign n1537 = N_N3924 & n1489;
  assign n1538 = N_N3923 & n979;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = N_N4057 & n1489;
  assign n1541_1 = N_N3793 & n979;
  assign n1542 = ~n1540 & ~n1541_1;
  assign n1543 = n1497 & ~n1504;
  assign n1544 = ~n1505 & ~n1543;
  assign n1545 = ~n1542 & ~n1544;
  assign n1546_1 = n1542 & n1544;
  assign n1547 = N_N3919 & n1489;
  assign n1548 = N_N3918 & n979;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1546_1 & ~n1549;
  assign n1551_1 = ~n1545 & ~n1550;
  assign n1552 = n1539 & n1551_1;
  assign n1553 = ~n1539 & ~n1551_1;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = n1536_1 & n1554;
  assign n1556_1 = ~n1536_1 & ~n1554;
  assign n1557 = ~n1555 & ~n1556_1;
  assign n1558 = n1490 & ~n1557;
  assign n1559 = N_N3981 & n1511_1;
  assign n229_1 = n1558 | n1559;
  assign n1561_1 = N_N3842 & ~n968;
  assign n1562 = N_N3196 & n972_1;
  assign n1563 = N_N3212 & n970;
  assign n1564 = ~n1562 & ~n1563;
  assign n234_1 = n1561_1 | ~n1564;
  assign n239_1 = N_N3105 & n948;
  assign n1567 = n1452 & n1475;
  assign n1568 = N_N4133 & n1454;
  assign n244_1 = n1567 | n1568;
  assign n1570 = ~NDN5_3 & ~NSr5_3;
  assign n1571_1 = ~PRESET & n1570;
  assign n1572 = n1234 & n1571_1;
  assign n1573 = ~PRESET & ~n1570;
  assign n1574 = N_N4117 & n1573;
  assign n249_1 = n1572 | n1574;
  assign n1576_1 = ~n1052 & n1479;
  assign n1577 = N_N3420 & n1486_1;
  assign n254 = n1576_1 | n1577;
  assign n1579 = N_N4179 & n1489;
  assign n1580 = N_N3071 & n979;
  assign n1581_1 = ~n1579 & ~n1580;
  assign n1582 = N_N3872 & n1489;
  assign n1583 = N_N3871 & n979;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1581_1 & n1584;
  assign n1586 = ~n1581_1 & ~n1584;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = N_N3868 & n1489;
  assign n1589 = N_N4099 & n979;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = N_N4165 & n1489;
  assign n1592 = N_N3776 & n979;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = ~n1590 & ~n1593;
  assign n1595 = n1590 & n1593;
  assign n1596 = ~n1536_1 & ~n1552;
  assign n1597 = ~n1553 & ~n1596;
  assign n1598 = ~n1595 & ~n1597;
  assign n1599 = ~n1594 & ~n1598;
  assign n1600 = ~n1587 & n1599;
  assign n1601 = n1587 & ~n1599;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = n1490 & n1602;
  assign n1604 = N_N3761 & n1511_1;
  assign n259_1 = n1603 | n1604;
  assign n264_1 = N_N3062 & n948;
  assign n1607 = N_N4071 & n1454;
  assign n1608 = n1452 & n1524;
  assign n269_1 = n1607 | n1608;
  assign n1610 = N_N4095 & ~n1108;
  assign n1611 = N_N3905 & n1112_1;
  assign n1612 = N_N3663 & n1116;
  assign n1613 = N_N4237 & n1110;
  assign n1614 = N_N3445 & n1114;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = ~n1611 & n1616;
  assign n1618 = ~n1610 & n1617;
  assign n1619 = ~n1303 & ~n1432;
  assign n1620 = ~n1431_1 & ~n1619;
  assign n1621 = ~n1618 & n1620;
  assign n1622 = n1618 & ~n1620;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = n1294 & ~n1623;
  assign n1625 = ~N_N4227 & n1624;
  assign n1626 = n1283 & n1623;
  assign n1627 = ~n1291 & ~n1626;
  assign n1628 = ~PRESET & N_N4227;
  assign n1629 = ~n1627 & n1628;
  assign n274 = n1625 | n1629;
  assign n1631 = N_N3807 & ~n968;
  assign n1632 = N_N3713 & n970;
  assign n1633 = N_N3235 & n972_1;
  assign n1634 = ~n1632 & ~n1633;
  assign n279_1 = n1631 | ~n1634;
  assign n1636 = N_N4145 & n1292;
  assign n1637 = ~n1405 & ~n1406_1;
  assign n1638 = n1415 & n1637;
  assign n1639 = ~n1415 & ~n1637;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = n1294 & ~n1640;
  assign n284 = n1636 | n1641;
  assign n1643 = n1278 & n1571_1;
  assign n1644 = N_N3922 & n1573;
  assign n289 = n1643 | n1644;
  assign n1646 = ~n1096 & n1479;
  assign n1647 = N_N3516 & n1486_1;
  assign n294 = n1646 | n1647;
  assign n1649 = N_N3813 & n1489;
  assign n1650 = N_N4239 & n979;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = N_N4206 & n1489;
  assign n1653 = N_N3630 & n979;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1651 & ~n1654;
  assign n1656 = n1651 & n1654;
  assign n1657 = ~n1585 & ~n1599;
  assign n1658 = ~n1586 & ~n1657;
  assign n1659 = ~n1656 & ~n1658;
  assign n1660 = ~n1655 & ~n1659;
  assign n1661 = N_N4132 & n1489;
  assign n1662 = N_N3069 & n979;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = N_N3843 & n1489;
  assign n1665 = N_N3842 & n979;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = n1663 & n1666;
  assign n1668 = ~n1663 & ~n1666;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = ~n1660 & ~n1669;
  assign n1671 = n1660 & n1669;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = n1490 & ~n1672;
  assign n1674 = N_N3489 & n1511_1;
  assign n299_1 = n1673 | n1674;
  assign n1676 = n1458 & n1571_1;
  assign n1677 = N_N4030 & n1573;
  assign n304_1 = n1676 | n1677;
  assign n1679 = ~n1273 & n1479;
  assign n1680 = N_N3540 & n1486_1;
  assign n309 = n1679 | n1680;
  assign n1682 = N_N4070 & n1489;
  assign n1683 = N_N3311 & n979;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = N_N3808 & n1489;
  assign n1686 = N_N3807 & n979;
  assign n1687 = ~n1685 & ~n1686;
  assign n1688 = n1684 & n1687;
  assign n1689 = ~n1684 & ~n1687;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = N_N4242 & n1489;
  assign n1692 = N_N3607 & n979;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = n1660 & ~n1668;
  assign n1695 = ~n1667 & ~n1694;
  assign n1696 = ~n1693 & n1695;
  assign n1697 = n1693 & ~n1695;
  assign n1698 = N_N3800 & n1489;
  assign n1699 = N_N4252 & n979;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = ~n1697 & ~n1700;
  assign n1702 = ~n1696 & ~n1701;
  assign n1703 = ~n1690 & n1702;
  assign n1704 = n1690 & ~n1702;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = n1490 & n1705;
  assign n1707 = N_N3513 & n1511_1;
  assign n314 = n1706 | n1707;
  assign n1709 = N_N4083 & n1292;
  assign n1710 = ~n1379 & ~n1380;
  assign n1711 = n1389 & n1710;
  assign n1712 = ~n1389 & ~n1710;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = n1294 & ~n1713;
  assign n319_1 = n1709 | n1714;
  assign n1716 = n1475 & n1571_1;
  assign n1717 = N_N3841 & n1573;
  assign n324_1 = n1716 | n1717;
  assign n1719 = N_N4018 & n1292;
  assign n1720 = ~n1353 & ~n1354;
  assign n1721 = n1363 & n1720;
  assign n1722 = ~n1363 & ~n1720;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = n1294 & ~n1723;
  assign n329 = n1719 | n1724;
  assign n1726 = N_N3971 & ~n968;
  assign n1727 = N_N3680 & n970;
  assign n1728 = N_N3681 & n972_1;
  assign n1729 = ~n1727 & ~n1728;
  assign n334 = n1726 | ~n1729;
  assign n339_1 = N_N4232 & n948;
  assign n1732 = ~n1233 & ~n1287;
  assign n1733 = N_N3460 & ~n1732;
  assign n1734 = ~N_N3578 & ~n1733;
  assign n1735 = n1292 & ~n1734;
  assign n1736 = n1233 & n1734;
  assign n1737 = ~PRESET & n1736;
  assign n1738 = ~n1735 & ~n1737;
  assign n1739 = N_N4246 & ~n1738;
  assign n1740 = ~N_N3961 & N_N4060;
  assign n1741 = ~N_N4126 & n1740;
  assign n1742 = ~N_N4004 & n1741;
  assign n1743 = ~N_N4171 & n1742;
  assign n1744 = ~N_N4036 & n1743;
  assign n1745 = ~N_N4212 & n1744;
  assign n1746 = ~N_N4093 & n1745;
  assign n1747 = ~N_N4246 & n1746;
  assign n1748 = N_N4246 & ~n1746;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n1294 & ~n1749;
  assign n1751 = ~n1233 & n1734;
  assign n1752 = ~n1290 & ~n1751;
  assign n1753 = ~PRESET & ~n1752;
  assign n1754 = ~n1197 & n1753;
  assign n1755 = ~n1750 & ~n1754;
  assign n344_1 = n1739 | ~n1755;
  assign n1757 = N_N3806 & n1573;
  assign n1758 = n1524 & n1571_1;
  assign n349_1 = n1757 | n1758;
  assign n1760 = N_N3992 & n1292;
  assign n1761 = ~n1327 & ~n1328;
  assign n1762 = n1337 & n1761;
  assign n1763 = ~n1337 & ~n1761;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = n1294 & ~n1764;
  assign n354 = n1760 | n1765;
  assign n1767 = N_N4086 & ~n968;
  assign n1768 = N_N3716 & n972_1;
  assign n1769 = N_N3715 & n970;
  assign n1770 = ~n1768 & ~n1769;
  assign n359 = n1767 | ~n1770;
  assign n364 = N_N4230 & n948;
  assign n1773 = N_N4212 & ~n1738;
  assign n1774 = N_N4212 & ~n1744;
  assign n1775 = ~n1745 & ~n1774;
  assign n1776 = n1294 & ~n1775;
  assign n1777 = ~n1149 & n1753;
  assign n1778 = ~n1776 & ~n1777;
  assign n369_1 = n1773 | ~n1778;
  assign n1441 = NDN5_9 & n965;
  assign n1781 = ~NDN5_16 & NLD3_9;
  assign n1782 = ~PRESET & Pnext_0_0_;
  assign n1783 = ~n1781 & n1782;
  assign n374_1 = n1441 | n1783;
  assign n1785 = ~NDN5_7 & ~NSr5_7;
  assign n1786 = ~PRESET & n1785;
  assign n1787 = N_N3965 & n1233;
  assign n1788 = n1786 & n1787;
  assign n1789 = ~PRESET & ~n1785;
  assign n1790 = N_N3626 & n1789;
  assign n378_1 = n1788 | n1790;
  assign n1792 = N_N3965 & n1292;
  assign n1793 = ~N_N3965 & n1321_1;
  assign n1794 = n1294 & ~n1322;
  assign n1795 = ~n1793 & n1794;
  assign n383_1 = n1792 | n1795;
  assign n1797 = N_N3890 & ~n968;
  assign n1798 = N_N3750 & n970;
  assign n1799 = N_N3751 & n972_1;
  assign n1800 = ~n1798 & ~n1799;
  assign n388_1 = n1797 | ~n1800;
  assign n1802 = ~PRESET & ~NGFDN_3;
  assign n393_1 = NDN3_11 & n1802;
  assign n1804 = ~NDN5_10 & NSr5_7;
  assign n398_1 = n965 & ~n1804;
  assign n403 = N_N3786 & n948;
  assign n1807 = N_N4171 & ~n1738;
  assign n1808 = N_N4171 & ~n1742;
  assign n1809 = ~n1743 & ~n1808;
  assign n1810 = n1294 & ~n1809;
  assign n1811 = ~n1218 & n1753;
  assign n1812 = ~n1810 & ~n1811;
  assign n408_1 = n1807 | ~n1812;
  assign n413_1 = NDN5_16 & n965;
  assign n1815 = N_N3992 & n1233;
  assign n1816 = n1786 & n1815;
  assign n1817 = N_N3799 & n1789;
  assign n418_1 = n1816 | n1817;
  assign n1819 = N_N3844 & ~n968;
  assign n1820 = N_N3875 & n970;
  assign n1821 = N_N3876 & n972_1;
  assign n1822 = ~n1820 & ~n1821;
  assign n423 = n1819 | ~n1822;
  assign n428_1 = N_N3196 & n948;
  assign n1825 = n1294 & n1741;
  assign n1826 = n1294 & ~n1740;
  assign n1827 = n1738 & ~n1826;
  assign n1828 = N_N4126 & ~n1827;
  assign n1829 = ~n1209 & n1753;
  assign n1830 = ~n1828 & ~n1829;
  assign n433_1 = n1825 | ~n1830;
  assign n438 = N_N3681 & n948;
  assign n1833 = N_N4018 & n1233;
  assign n1834 = n1786 & n1833;
  assign n1835 = N_N3679 & n1789;
  assign n443 = n1834 | n1835;
  assign n1837 = N_N3340 & n1735;
  assign n1838 = ~N_N3369 & n1747;
  assign n1839 = ~N_N3283 & n1838;
  assign n1840 = ~N_N3340 & n1283;
  assign n1841 = n1839 & n1840;
  assign n1842 = n1283 & ~n1839;
  assign n1843 = ~n1736 & ~n1842;
  assign n1844 = N_N3340 & ~n1843;
  assign n1845 = ~n1188 & ~n1752;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = ~n1841 & n1846;
  assign n1848 = ~PRESET & ~n1847;
  assign n448_1 = n1837 | n1848;
  assign n1850 = ~NDN5_4 & ~NSr5_4;
  assign n1851 = ~PRESET & n1850;
  assign n1852 = n1234 & n1851;
  assign n1853 = ~PRESET & ~n1850;
  assign n1854 = N_N4116 & n1853;
  assign n453 = n1852 | n1854;
  assign n1856 = N_N3810 & ~n968;
  assign n1857 = N_N3931 & n970;
  assign n1858 = N_N3932 & n972_1;
  assign n1859 = ~n1857 & ~n1858;
  assign n458_1 = n1856 | ~n1859;
  assign n463_1 = N_N3235 & n948;
  assign n1862 = N_N3283 & ~n1738;
  assign n1863 = N_N3283 & ~n1838;
  assign n1864 = ~n1839 & ~n1863;
  assign n1865 = n1294 & ~n1864;
  assign n1866 = ~n1121 & n1753;
  assign n1867 = ~n1865 & ~n1866;
  assign n468 = n1862 | ~n1867;
  assign n473_1 = N_N3716 & n948;
  assign n1870 = N_N4083 & n1233;
  assign n1871 = n1786 & n1870;
  assign n1872 = N_N3701 & n1789;
  assign n478_1 = n1871 | n1872;
  assign n1874 = n1278 & n1851;
  assign n1875 = N_N3921 & n1853;
  assign n483 = n1874 | n1875;
  assign n1877 = ~NDN5_8 & ~NSr5_8;
  assign n1878 = ~PRESET & n1877;
  assign n1879 = n1787 & n1878;
  assign n1880 = ~PRESET & ~n1877;
  assign n1881 = N_N3625 & n1880;
  assign n488 = n1879 | n1881;
  assign n493_1 = N_N3751 & n948;
  assign n1884 = N_N3736 & n1789;
  assign n1885 = N_N4145 & n1233;
  assign n1886 = n1786 & n1885;
  assign n498 = n1884 | n1886;
  assign n1888 = n1458 & n1851;
  assign n1889 = N_N3870 & n1853;
  assign n503 = n1888 | n1889;
  assign n1891 = n1815 & n1878;
  assign n1892 = N_N4024 & n1880;
  assign n508_1 = n1891 | n1892;
  assign n513 = N_N3876 & n948;
  assign n1895 = n1475 & n1851;
  assign n1896 = N_N3840 & n1853;
  assign n518_1 = n1895 | n1896;
  assign n1898 = n1833 & n1878;
  assign n1899 = N_N4021 & n1880;
  assign n523 = n1898 | n1899;
  assign n528_1 = N_N3932 & n948;
  assign n533_1 = ~PRESET & ~PDN;
  assign n1903 = n1524 & n1851;
  assign n1904 = N_N3805 & n1853;
  assign n538 = n1903 | n1904;
  assign n1906 = n1870 & n1878;
  assign n1907 = N_N3700 & n1880;
  assign n543_1 = n1906 | n1907;
  assign n1909 = n1878 & n1885;
  assign n1910 = N_N3735 & n1880;
  assign n548 = n1909 | n1910;
  assign n1912 = Pready_0_0_ & ~NLak3_2;
  assign n1913 = ~PDN & n1912;
  assign n1914 = n960 & n1913;
  assign n1915 = NSr3_2 & n1914;
  assign n553_1 = ~PRESET & n1915;
  assign n1917 = N_N4205 & ~N_N3336;
  assign n1918 = ~N_N4205 & N_N3336;
  assign n1919 = ~N_N3882 & N_N3884;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~N_N4015 & N_N3908;
  assign n1922 = N_N4054 & ~N_N3489;
  assign n1923 = N_N4015 & ~N_N3908;
  assign n1924 = ~N_N4243 & N_N3862;
  assign n1925 = ~N_N3761 & N_N4056;
  assign n1926 = N_N4243 & ~N_N3862;
  assign n1927 = ~N_N3574 & N_N3832;
  assign n1928 = ~N_N3981 & N_N3778;
  assign n1929 = N_N3574 & ~N_N3832;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = N_N3535 & ~N_N3797;
  assign n1932 = N_N3916 & ~N_N4111;
  assign n1933 = ~n1931 & n1932;
  assign n1934 = N_N3733 & ~N_N3794;
  assign n1935 = ~N_N3535 & N_N3797;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1933 & n1936;
  assign n1938 = ~N_N3733 & N_N3794;
  assign n1939 = N_N3981 & ~N_N3778;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n1937 & n1940;
  assign n1942 = n1930 & ~n1941;
  assign n1943 = N_N3761 & ~N_N4056;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1927 & n1944;
  assign n1946 = ~n1926 & ~n1945;
  assign n1947 = ~n1925 & n1946;
  assign n1948 = ~N_N4054 & N_N3489;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1924 & n1949;
  assign n1951 = ~n1923 & ~n1950;
  assign n1952 = ~n1922 & n1951;
  assign n1953 = ~N_N3818 & N_N3513;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = ~n1921 & n1954;
  assign n1956 = N_N3818 & ~N_N3513;
  assign n1957 = N_N3882 & ~N_N3884;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = ~n1955 & n1958;
  assign n1960 = n1920 & ~n1959;
  assign n1961 = NLD3_9 & ~n1960;
  assign n1962 = ~n1917 & n1961;
  assign n558 = ~PRESET & n1962;
  assign n1964 = N_N3906 & n948;
  assign n1965 = Pdxport_0_0_ & n950;
  assign n563_1 = n1964 | n1965;
  assign n1967 = ~N_N3388 & ~n955;
  assign n568_1 = ~PRESET & ~n1967;
  assign n1969 = N_N4057 & n948;
  assign n1970 = Pdxport_2_2_ & n950;
  assign n573_1 = n1969 | n1970;
  assign n578 = N_N3011 & n948;
  assign n1973 = ~N_N3346 & ~n955;
  assign n583_1 = ~PRESET & ~n1973;
  assign n1975 = n1493 & n1496_1;
  assign n1976 = ~n1497 & ~n1975;
  assign n1977 = n1479 & n1976;
  assign n1978 = N_N3677 & n1486_1;
  assign n588 = n1977 | n1978;
  assign n1980 = N_N4165 & n948;
  assign n1981 = Pdxport_4_4_ & n950;
  assign n593 = n1980 | n1981;
  assign n598 = N_N4080 & n948;
  assign n603 = N_N3373 & n948;
  assign n1985 = ~n1545 & ~n1546_1;
  assign n1986 = n1549 & ~n1985;
  assign n1987 = ~n1549 & n1985;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = n1479 & n1988;
  assign n1990 = N_N3709 & n1486_1;
  assign n608 = n1989 | n1990;
  assign n1992 = N_N4206 & n948;
  assign n1993 = Pdxport_6_6_ & n950;
  assign n613_1 = n1992 | n1993;
  assign n618_1 = N_N3324 & n1060;
  assign n1996 = N_N4093 & ~n1745;
  assign n1997 = ~n1746 & ~n1996;
  assign n1998 = N_N4004 & ~n1741;
  assign n1999 = ~n1742 & ~n1998;
  assign n2000 = ~N_N3283 & ~N_N3369;
  assign n2001 = ~N_N4246 & n2000;
  assign n2002 = ~N_N4126 & ~N_N3961;
  assign n2003 = n2001 & n2002;
  assign n2004 = n1840 & n2003;
  assign n2005 = n1999 & n2004;
  assign n2006 = ~N_N4212 & ~N_N4036;
  assign n2007 = ~N_N4060 & n2006;
  assign n2008 = ~N_N4171 & n2007;
  assign n2009 = n2005 & n2008;
  assign n2010 = n1997 & n2009;
  assign n623_1 = ~PRESET & n2010;
  assign n628 = N_N4159 & n948;
  assign n633 = ~PRESET & ~n1733;
  assign n2014 = N_N3916 & n948;
  assign n2015 = Paport_0_0_ & n950;
  assign n638_1 = n2014 | n2015;
  assign n2017 = ~n1594 & ~n1595;
  assign n2018 = n1597 & ~n2017;
  assign n2019 = ~n1597 & n2017;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = n1479 & n2020;
  assign n2022 = N_N3743 & n1486_1;
  assign n643 = n2021 | n2022;
  assign n2024 = N_N4242 & n948;
  assign n2025 = Pdxport_8_8_ & n950;
  assign n648_1 = n2024 | n2025;
  assign n653_1 = N_N3312 & n1060;
  assign n2028 = N_N3733 & n948;
  assign n2029 = Paport_2_2_ & n950;
  assign n658 = n2028 | n2029;
  assign n2031 = n1655 & ~n1658;
  assign n2032 = n1656 & n1658;
  assign n2033 = n1660 & ~n2032;
  assign n2034 = ~n2031 & ~n2033;
  assign n2035 = n1479 & ~n2034;
  assign n2036 = N_N3774 & n1486_1;
  assign n663 = n2035 | n2036;
  assign n2038 = N_N4214 & ~n2010;
  assign n2039 = ~n1290 & ~n2038;
  assign n2040 = N_N3462 & ~n2039;
  assign n668_1 = ~PRESET & n2040;
  assign n673 = N_N3294 & n1060;
  assign n2043 = n990 & n1036;
  assign n2044 = ~n1037_1 & ~n2043;
  assign n2045 = n977_1 & n2044;
  assign n2046 = N_N3796 & n1054;
  assign n678_1 = n2045 | n2046;
  assign n2048 = N_N3574 & n948;
  assign n2049 = Paport_4_4_ & n950;
  assign n683 = n2048 | n2049;
  assign n2051 = ~n1696 & ~n1697;
  assign n2052 = n1700 & ~n2051;
  assign n2053 = ~n1700 & n2051;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n1479 & n2054;
  assign n2056 = N_N3791 & n1486_1;
  assign n688_1 = n2055 | n2056;
  assign n2058 = ~n1025 & ~n1026;
  assign n2059 = n1039 & ~n2058;
  assign n2060 = ~n1039 & n2058;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = n977_1 & n2061;
  assign n2063 = N_N3480 & n1054;
  assign n693 = n2062 | n2063;
  assign n2065 = N_N4243 & n948;
  assign n2066 = Paport_6_6_ & n950;
  assign n698_1 = n2065 | n2066;
  assign n2068 = N_N3940 & ~n968;
  assign n2069 = N_N4111 & n970;
  assign n2070 = N_N4218 & n972_1;
  assign n2071 = ~n2069 & ~n2070;
  assign n703_1 = n2068 | ~n2071;
  assign n2073 = ~n1015 & ~n1016;
  assign n2074 = ~n1047 & ~n2073;
  assign n2075 = n1047 & n2073;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = n977_1 & ~n2076;
  assign n2078 = N_N3509 & n1054;
  assign n708 = n2077 | n2078;
  assign n2080 = N_N4015 & n948;
  assign n2081 = Paport_8_8_ & n950;
  assign n713_1 = n2080 | n2081;
  assign n2083 = ~N_N2989 & ~n955;
  assign n718 = ~PRESET & ~n2083;
  assign n2085 = N_N3919 & ~n968;
  assign n2086 = N_N3794 & n970;
  assign n2087 = N_N3417 & n972_1;
  assign n2088 = ~n2086 & ~n2087;
  assign n723 = n2085 | ~n2088;
  assign n2090 = ~PRESET & n1733;
  assign n728 = N_N3578 & n2090;
  assign n2092 = ~n1076 & ~n1077_1;
  assign n2093 = n1079 & ~n2092;
  assign n2094 = ~n1079 & n2092;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = n977_1 & n2095;
  assign n2097 = N_N3529 & n1054;
  assign n733 = n2096 | n2097;
  assign n738 = N_N4222 & n1060;
  assign n2100 = n1102 & n1787;
  assign n2101 = N_N3910 & n1236_1;
  assign n743 = n2100 | n2101;
  assign n2103 = N_N3868 & ~n968;
  assign n2104 = N_N3832 & n970;
  assign n2105 = N_N3262 & n972_1;
  assign n2106 = ~n2104 & ~n2105;
  assign n748_1 = n2103 | ~n2106;
  assign n2108 = ~n1261_1 & ~n1262;
  assign n2109 = ~n1265 & ~n2108;
  assign n2110 = n1265 & n2108;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = n977_1 & ~n2111;
  assign n2113 = N_N3947 & n1054;
  assign n753 = n2112 | n2113;
  assign n758 = N_N4181 & n1060;
  assign n2116 = n1102 & n1815;
  assign n2117 = N_N3793 & n1236_1;
  assign n763 = n2116 | n2117;
  assign n768 = N_N3822 & n948;
  assign n2120 = N_N3813 & ~n968;
  assign n2121 = N_N3862 & n970;
  assign n2122 = N_N3280 & n972_1;
  assign n2123 = ~n2121 & ~n2122;
  assign n773_1 = n2120 | ~n2123;
  assign n2125 = N_N3470 & n976;
  assign n2126 = N_N3274 & n979;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = n1253 & ~n1268;
  assign n2129 = ~n1269 & ~n2128;
  assign n2130 = n2127 & n2129;
  assign n2131 = ~n2127 & ~n2129;
  assign n2132 = N_N3482 & n976;
  assign n2133 = N_N4075 & n979;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~n1251_1 & ~n2134;
  assign n2136 = n1251_1 & n2134;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2131 & ~n2137;
  assign n2139 = ~n2130 & ~n2138;
  assign n2140 = N_N4039 & n976;
  assign n2141 = N_N3612 & n979;
  assign n2142 = ~n2140 & ~n2141;
  assign n2143 = N_N4095 & n976;
  assign n2144 = N_N4167 & n979;
  assign n2145 = ~n2143 & ~n2144;
  assign n2146 = ~n2142 & n2145;
  assign n2147 = n2142 & ~n2145;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = ~n2136 & n2148;
  assign n2150 = n2136 & ~n2148;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = n2139 & n2151;
  assign n2153 = ~n2139 & ~n2151;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = n1479 & ~n2154;
  assign n2156 = N_N4114 & n1486_1;
  assign n778_1 = n2155 | n2156;
  assign n783_1 = N_N4134 & n1060;
  assign n788 = N_N3866 & n948;
  assign n793_1 = N_N4218 & n948;
  assign n2161 = N_N3939 & ~n968;
  assign n2162 = N_N3741 & n972_1;
  assign n2163 = N_N3677 & n970;
  assign n2164 = ~n2162 & ~n2163;
  assign n798 = n2161 | ~n2164;
  assign n2166 = n1102 & n1833;
  assign n2167 = N_N3776 & n1236_1;
  assign n803_1 = n2166 | n2167;
  assign n2169 = n1452 & n1787;
  assign n2170 = N_N3387 & n1454;
  assign n808_1 = n2169 | n2170;
  assign n2172 = N_N4194 & n948;
  assign n2173 = Pdxport_10_10_ & n950;
  assign n813 = n2172 | n2173;
  assign n2175 = ~n2130 & ~n2131;
  assign n2176 = ~n2137 & n2175;
  assign n2177 = n2137 & ~n2175;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = n1479 & ~n2178;
  assign n2180 = N_N3821 & n1486_1;
  assign n818_1 = n2179 | n2180;
  assign n2182 = N_N3882 & n948;
  assign n2183 = Paport_10_10_ & n950;
  assign n823_1 = n2182 | n2183;
  assign n2185 = n977_1 & ~n2154;
  assign n2186 = N_N4167 & n1054;
  assign n828_1 = n2185 | n2186;
  assign n2188 = N_N3800 & ~n968;
  assign n2189 = N_N3908 & n970;
  assign n2190 = N_N3634 & n972_1;
  assign n2191 = ~n2189 & ~n2190;
  assign n833 = n2188 | ~n2191;
  assign n2193 = N_N4237 & n948;
  assign n2194 = Pdxport_11_11_ & n950;
  assign n838_1 = n2193 | n2194;
  assign n843_1 = N_N3417 & n948;
  assign n2197 = N_N3918 & ~n968;
  assign n2198 = N_N3356 & n972_1;
  assign n2199 = N_N3709 & n970;
  assign n2200 = ~n2198 & ~n2199;
  assign n848_1 = n2197 | ~n2200;
  assign n2202 = N_N4177 & n1489;
  assign n2203 = N_N4176 & n979;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = ~n1688 & ~n1702;
  assign n2206 = ~n1689 & ~n2205;
  assign n2207 = ~n2204 & ~n2206;
  assign n2208 = n2204 & n2206;
  assign n2209 = N_N4194 & n1489;
  assign n2210 = N_N4193 & n979;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n2208 & ~n2211;
  assign n2213 = ~n2207 & ~n2212;
  assign n2214 = N_N4237 & n1489;
  assign n2215 = N_N4236 & n979;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = N_N4209 & n1489;
  assign n2218 = N_N4208 & n979;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = ~n2216 & n2219;
  assign n2221 = n2216 & ~n2219;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = n2213 & n2222;
  assign n2224 = ~n2213 & ~n2222;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = n1479 & n2225;
  assign n2227 = N_N4158 & n1486_1;
  assign n853 = n2226 | n2227;
  assign n2229 = n1102 & n1870;
  assign n2230 = N_N3630 & n1236_1;
  assign n858_1 = n2229 | n2230;
  assign n2232 = N_N3344 & n1454;
  assign n2233 = n1452 & n1815;
  assign n863_1 = n2232 | n2233;
  assign n868 = N_N4072 & n1060;
  assign n2236 = n977_1 & ~n2178;
  assign n2237 = N_N3274 & n1054;
  assign n873_1 = n2236 | n2237;
  assign n2239 = N_N3473 & n1454;
  assign n2240 = N_N4197 & n1233;
  assign n2241 = n1452 & n2240;
  assign n878_1 = n2239 | n2241;
  assign n2243 = N_N4205 & n948;
  assign n2244 = Paport_11_11_ & n950;
  assign n883 = n2243 | n2244;
  assign n2246 = n1490 & n1976;
  assign n2247 = N_N4111 & n1511_1;
  assign n888_1 = n2246 | n2247;
  assign n2249 = n1479 & n2044;
  assign n2250 = N_N3680 & n1486_1;
  assign n893 = n2249 | n2250;
  assign n2252 = ~N_N3838 & ~n1289;
  assign n898 = ~PRESET & ~n2252;
  assign n903 = N_N3262 & n948;
  assign n2255 = N_N4099 & ~n968;
  assign n2256 = N_N3384 & n972_1;
  assign n2257 = N_N3743 & n970;
  assign n2258 = ~n2256 & ~n2257;
  assign n908 = n2255 | ~n2258;
  assign n2260 = N_N3607 & n1236_1;
  assign n2261 = n1102 & n1885;
  assign n913 = n2260 | n2261;
  assign n2263 = N_N3323 & n1454;
  assign n2264 = n1452 & n1833;
  assign n918_1 = n2263 | n2264;
  assign n2266 = N_N4227 & n1233;
  assign n2267 = n1878 & n2266;
  assign n2268 = N_N3612 & n1880;
  assign n923 = n2267 | n2268;
  assign n2270 = ~n2207 & ~n2208;
  assign n2271 = n2211 & ~n2270;
  assign n2272 = ~n2211 & n2270;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = n1479 & n2273;
  assign n2275 = N_N4079 & n1486_1;
  assign n928 = n2274 | n2275;
  assign n2277 = ~NGFDN_3 & ~n958;
  assign n933 = n533_1 & ~n2277;
  assign n2279 = N_N3457 & n1573;
  assign n2280 = n1571_1 & n2240;
  assign n937 = n2279 | n2280;
  assign n942 = N_N3445 & n1060;
  assign n2283 = n1490 & n1988;
  assign n2284 = N_N3794 & n1511_1;
  assign n947_1 = n2283 | n2284;
  assign n2286 = N_N3663 & n1454;
  assign n2287 = n1452 & n2266;
  assign n952 = n2286 | n2287;
  assign n2289 = n1479 & n2061;
  assign n2290 = N_N3715 & n1486_1;
  assign n957_1 = n2289 | n2290;
  assign n2292 = n1786 & n2266;
  assign n2293 = N_N4039 & n1789;
  assign n962_1 = n2292 | n2293;
  assign n967 = N_N3280 & n948;
  assign n2296 = N_N4239 & ~n968;
  assign n2297 = N_N4090 & n972_1;
  assign n2298 = N_N3774 & n970;
  assign n2299 = ~n2297 & ~n2298;
  assign n972 = n2296 | ~n2299;
  assign n2301 = n1452 & n1870;
  assign n2302 = N_N3988 & n1454;
  assign n977 = n2301 | n2302;
  assign n2304 = N_N3433 & n1573;
  assign n2305 = n1571_1 & n2266;
  assign n982 = n2304 | n2305;
  assign n2307 = n1878 & n2240;
  assign n2308 = N_N4075 & n1880;
  assign n987_1 = n2307 | n2308;
  assign n992 = N_N3468 & n1060;
  assign n2311 = N_N4045 & n1853;
  assign n2312 = n1851 & n2240;
  assign n997_1 = n2311 | n2312;
  assign n2314 = N_N3482 & n1789;
  assign n2315 = n1786 & n2240;
  assign n1002 = n2314 | n2315;
  assign n2317 = n1490 & n2020;
  assign n2318 = N_N3832 & n1511_1;
  assign n1007_1 = n2317 | n2318;
  assign n2320 = n1571_1 & n1787;
  assign n2321 = N_N3304 & n1573;
  assign n1012_1 = n2320 | n2321;
  assign n2323 = n1479 & ~n2076;
  assign n2324 = N_N3750 & n1486_1;
  assign n1017_1 = n2323 | n2324;
  assign n1022 = N_N3634 & n948;
  assign n2327 = N_N3293 & n1454;
  assign n2328 = n1452 & n1885;
  assign n1027 = n2327 | n2328;
  assign n2330 = n1851 & n2266;
  assign n2331 = N_N3659 & n1853;
  assign n1032_1 = n2330 | n2331;
  assign n2333 = N_N4252 & ~n968;
  assign n2334 = N_N3533 & n972_1;
  assign n2335 = N_N3791 & n970;
  assign n2336 = ~n2334 & ~n2335;
  assign n1037 = n2333 | ~n2336;
  assign n2338 = N_N3912 & n1292;
  assign n2339 = ~n1418 & ~n1419;
  assign n2340 = n1428 & n2339;
  assign n2341 = ~n1428 & ~n2339;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = n1294 & ~n2342;
  assign n1042_1 = n2338 | n2343;
  assign n2345 = n1490 & ~n2034;
  assign n2346 = N_N3862 & n1511_1;
  assign n1047_1 = n2345 | n2346;
  assign n2348 = n1571_1 & n1815;
  assign n2349 = N_N3221 & n1573;
  assign n1052_1 = n2348 | n2349;
  assign n2351 = n1479 & n2095;
  assign n2352 = N_N3875 & n1486_1;
  assign n1057 = n2351 | n2352;
  assign n2354 = N_N3949 & n1292;
  assign n2355 = ~n1392 & ~n1393;
  assign n2356 = n1402 & n2355;
  assign n2357 = ~n1402 & ~n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = n1294 & ~n2358;
  assign n1062_1 = n2354 | n2359;
  assign n2361 = n1490 & n2054;
  assign n2362 = N_N3908 & n1511_1;
  assign n1067_1 = n2361 | n2362;
  assign n2364 = n1571_1 & n1833;
  assign n2365 = N_N3711 & n1573;
  assign n1072_1 = n2364 | n2365;
  assign n2367 = n1479 & ~n2111;
  assign n2368 = N_N3931 & n1486_1;
  assign n1077 = n2367 | n2368;
  assign n1082_1 = N_N3469 & n1060;
  assign n2371 = n1571_1 & n1870;
  assign n2372 = N_N3436 & n1573;
  assign n1087 = n2371 | n2372;
  assign n2374 = N_N3974 & n1292;
  assign n2375 = ~n1366_1 & ~n1367;
  assign n2376 = n1376_1 & n2375;
  assign n2377 = ~n1376_1 & ~n2375;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = n1294 & ~n2378;
  assign n1092 = n2374 | n2379;
  assign n1097 = N_N3905 & n1060;
  assign n1102_1 = N_N3741 & n948;
  assign n2383 = N_N3369 & ~n1738;
  assign n2384 = N_N3369 & ~n1747;
  assign n2385 = ~n1838 & ~n2384;
  assign n2386 = n1294 & ~n2385;
  assign n2387 = ~n1131 & n1753;
  assign n2388 = ~n2386 & ~n2387;
  assign n1107 = n2383 | ~n2388;
  assign n2390 = N_N3164 & n1573;
  assign n2391 = n1571_1 & n1885;
  assign n1112 = n2390 | n2391;
  assign n2393 = N_N3500 & ~n968;
  assign n2394 = N_N3331 & n972_1;
  assign n2395 = N_N3464 & n970;
  assign n2396 = ~n2394 & ~n2395;
  assign n1117_1 = n2393 | ~n2396;
  assign n2398 = N_N3996 & n1292;
  assign n2399 = ~n1340 & ~n1341_1;
  assign n2400 = n1350 & n2399;
  assign n2401 = ~n1350 & ~n2399;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = n1294 & ~n2402;
  assign n1122 = n2398 | n2403;
  assign n1127_1 = N_N3356 & n948;
  assign n2406 = N_N4093 & ~n1738;
  assign n2407 = n1294 & ~n1997;
  assign n2408 = ~n1227 & n1753;
  assign n2409 = ~n2407 & ~n2408;
  assign n1132 = n2406 | ~n2409;
  assign n1176 = ~NSr3_9 & n1802;
  assign n2412 = ~NDN3_11 & NGFDN_3;
  assign n2413 = ~PRESET & Pover_0_0_;
  assign n2414 = ~n2412 & n2413;
  assign n1137 = n1176 | n2414;
  assign n2416 = N_N4224 & ~n968;
  assign n2417 = N_N4106 & n972_1;
  assign n2418 = N_N3442 & n970;
  assign n2419 = ~n2417 & ~n2418;
  assign n1141_1 = n2416 | ~n2419;
  assign n2421 = N_N4027 & n1292;
  assign n2422 = ~n1323 & n1325;
  assign n2423 = ~n1323 & ~n1324;
  assign n2424 = ~N_N4027 & ~n2423;
  assign n2425 = n1294 & ~n2424;
  assign n2426 = ~n2422 & n2425;
  assign n1146 = n2421 | n2426;
  assign n1151 = NDN1_4 & n533_1;
  assign n1156 = N_N3384 & n948;
  assign n2430 = N_N4036 & ~n1738;
  assign n2431 = N_N4036 & ~n1743;
  assign n2432 = ~n1744 & ~n2431;
  assign n2433 = n1294 & ~n2432;
  assign n2434 = ~n1140 & n1753;
  assign n2435 = ~n2433 & ~n2434;
  assign n1161 = n2430 | ~n2435;
  assign n2437 = n1234 & n1786;
  assign n2438 = N_N3968 & n1789;
  assign n1166 = n2437 | n2438;
  assign n2440 = N_N4183 & ~n968;
  assign n2441 = N_N3393 & n972_1;
  assign n2442 = N_N3420 & n970;
  assign n2443 = ~n2441 & ~n2442;
  assign n1171 = n2440 | ~n2443;
  assign n1181_1 = N_N4090 & n948;
  assign n2446 = N_N4004 & ~n1738;
  assign n2447 = n1294 & ~n1999;
  assign n2448 = ~n1160 & n1753;
  assign n2449 = ~n2447 & ~n2448;
  assign n1186_1 = n2446 | ~n2449;
  assign n2451 = n1278 & n1786;
  assign n2452 = N_N3205 & n1789;
  assign n1191_1 = n2451 | n2452;
  assign n2454 = N_N4136 & ~n968;
  assign n2455 = N_N3517 & n972_1;
  assign n2456 = N_N3516 & n970;
  assign n2457 = ~n2455 & ~n2456;
  assign n1196_1 = n2454 | ~n2457;
  assign n2459 = n1787 & n1851;
  assign n2460 = N_N3303 & n1853;
  assign n1201_1 = n2459 | n2460;
  assign n1206_1 = N_N3533 & n948;
  assign n2463 = N_N3336 & n1511_1;
  assign n2464 = n1490 & n2225;
  assign n1211_1 = n2463 | n2464;
  assign n2466 = ~n1178 & n1753;
  assign n2467 = ~N_N4060 & n1294;
  assign n2468 = n1738 & ~n2467;
  assign n2469 = N_N3961 & ~n2468;
  assign n2470 = n1294 & n1740;
  assign n2471 = ~n2469 & ~n2470;
  assign n1216_1 = n2466 | ~n2471;
  assign n1221_1 = N_N3331 & n948;
  assign n2474 = n1458 & n1786;
  assign n2475 = N_N3203 & n1789;
  assign n1226_1 = n2474 | n2475;
  assign n2477 = N_N4236 & n1236_1;
  assign n2478 = n1102 & n2266;
  assign n1231 = n2477 | n2478;
  assign n2480 = n1490 & n2273;
  assign n2481 = N_N3884 & n1511_1;
  assign n1236 = n2480 | n2481;
  assign n2483 = n1815 & n1851;
  assign n2484 = N_N3367 & n1853;
  assign n1241 = n2483 | n2484;
  assign n2486 = N_N4140 & ~n968;
  assign n2487 = N_N3540 & n970;
  assign n2488 = N_N3541 & n972_1;
  assign n2489 = ~n2487 & ~n2488;
  assign n1246 = n2486 | ~n2489;
  assign n2491 = NDN2_2 & ~n954;
  assign n1251 = ~PRESET & n2491;
  assign n1256 = N_N4106 & n948;
  assign n2494 = n1475 & n1786;
  assign n2495 = N_N3100 & n1789;
  assign n1261 = n2494 | n2495;
  assign n2497 = N_N4193 & n1236_1;
  assign n2498 = n1102 & n2240;
  assign n1266 = n2497 | n2498;
  assign n2500 = N_N3470 & ~n968;
  assign n2501 = N_N3821 & n970;
  assign n2502 = N_N3822 & n972_1;
  assign n2503 = ~n2501 & ~n2502;
  assign n1271_1 = n2500 | ~n2503;
  assign n2505 = n1833 & n1851;
  assign n2506 = N_N3424 & n1853;
  assign n1276_1 = n2505 | n2506;
  assign n2508 = n1234 & n1878;
  assign n2509 = N_N3959 & n1880;
  assign n1281 = n2508 | n2509;
  assign n1286_1 = N_N3393 & n948;
  assign n2512 = n1524 & n1786;
  assign n2513 = N_N4042 & n1789;
  assign n1291_1 = n2512 | n2513;
  assign n2515 = n1851 & n1870;
  assign n2516 = N_N3188 & n1853;
  assign n1296_1 = n2515 | n2516;
  assign n2518 = N_N4095 & ~n968;
  assign n2519 = N_N4114 & n970;
  assign n2520 = N_N3866 & n972_1;
  assign n2521 = ~n2519 & ~n2520;
  assign n1301 = n2518 | ~n2521;
  assign n2523 = n1278 & n1878;
  assign n2524 = N_N3957 & n1880;
  assign n1306 = n2523 | n2524;
  assign n1311 = N_N3517 & n948;
  assign n2527 = n1851 & n1885;
  assign n2528 = N_N4047 & n1853;
  assign n1316 = n2527 | n2528;
  assign n2530 = n1458 & n1878;
  assign n2531 = N_N3081 & n1880;
  assign n1321 = n2530 | n2531;
  assign n1326 = N_N3541 & n948;
  assign n2534 = N_N4177 & ~n968;
  assign n2535 = N_N3011 & n972_1;
  assign n2536 = N_N3884 & n970;
  assign n2537 = ~n2535 & ~n2536;
  assign n1331 = n2534 | ~n2537;
  assign n2539 = ~NDN3_3 & NSr3_2;
  assign n1336 = n1802 & ~n2539;
  assign n2541 = N_N4176 & ~n968;
  assign n2542 = N_N4079 & n970;
  assign n2543 = N_N4080 & n972_1;
  assign n2544 = ~n2542 & ~n2543;
  assign n1341 = n2541 | ~n2544;
  assign n2546 = n1475 & n1878;
  assign n2547 = N_N3585 & n1880;
  assign n1346 = n2546 | n2547;
  assign n2549 = ~NDN3_3 & ~NDN3_8;
  assign n1351 = n1802 & ~n2549;
  assign n2551 = N_N4209 & ~n968;
  assign n2552 = N_N3336 & n970;
  assign n2553 = N_N3373 & n972_1;
  assign n2554 = ~n2552 & ~n2553;
  assign n1356 = n2551 | ~n2554;
  assign n2556 = n1524 & n1878;
  assign n2557 = N_N3824 & n1880;
  assign n1361 = n2556 | n2557;
  assign n2559 = N_N4208 & ~n968;
  assign n2560 = N_N4158 & n970;
  assign n2561 = N_N4159 & n972_1;
  assign n2562 = ~n2560 & ~n2561;
  assign n1366 = n2559 | ~n2562;
  assign n2564 = N_N4120 & n948;
  assign n2565 = Pdxport_1_1_ & n950;
  assign n1371 = n2564 | n2565;
  assign n1376 = N_N3708 & n1060;
  assign n2568 = N_N4220 & n948;
  assign n2569 = Pdxport_3_3_ & n950;
  assign n1381 = n2568 | n2569;
  assign n2571 = ~N_N3999 & ~n1289;
  assign n1386 = n2090 & ~n2571;
  assign n1391 = N_N4223 & n1060;
  assign n2574 = n1479 & ~n1509;
  assign n2575 = N_N3179 & n1486_1;
  assign n1396 = n2574 | n2575;
  assign n2577 = N_N4179 & n948;
  assign n2578 = Pdxport_5_5_ & n950;
  assign n1401 = n2577 | n2578;
  assign n2580 = n1479 & ~n1557;
  assign n2581 = N_N3475 & n1486_1;
  assign n1406 = n2580 | n2581;
  assign n2583 = N_N4132 & n948;
  assign n2584 = Pdxport_7_7_ & n950;
  assign n1411 = n2583 | n2584;
  assign n1416 = N_N4182 & n1060;
  assign n2587 = N_N3797 & n948;
  assign n2588 = Paport_1_1_ & n950;
  assign n1421 = n2587 | n2588;
  assign n2590 = n1479 & n1602;
  assign n2591 = N_N3214 & n1486_1;
  assign n1426 = n2590 | n2591;
  assign n2593 = N_N4070 & n948;
  assign n2594 = Pdxport_9_9_ & n950;
  assign n1431 = n2593 | n2594;
  assign n1436 = N_N4135 & n1060;
  assign n1446 = ~PRESET & ~NSr5_2;
  assign n1451 = ~PRESET & ~NSr5_3;
  assign n2599 = N_N3778 & n948;
  assign n2600 = Paport_3_3_ & n950;
  assign n1456 = n2599 | n2600;
  assign n1461 = ~PRESET & ~NSr5_4;
  assign n2603 = n1479 & ~n1672;
  assign n2604 = N_N3212 & n1486_1;
  assign n1466 = n2603 | n2604;
  assign n1471 = ~PRESET & ~NSr5_5;
  assign n2607 = ~NDN5_6 & ~n1105;
  assign n1476 = n965 & ~n2607;
  assign n1481 = ~PRESET & ~NSr5_7;
  assign n1486 = ~PRESET & ~NSr5_8;
  assign n1491 = N_N4073 & n1060;
  assign n2612 = NEN5_9 & n965;
  assign n1496 = n1441 | n2612;
  assign n2614 = ~NSr5_8 & n965;
  assign n1501 = n2612 | n2614;
  assign n2616 = n977_1 & n1484;
  assign n2617 = N_N3684 & n1054;
  assign n1506 = n2616 | n2617;
  assign n2619 = N_N4056 & n948;
  assign n2620 = Paport_5_5_ & n950;
  assign n1511 = n2619 | n2620;
  assign n2622 = n1479 & n1705;
  assign n2623 = N_N3713 & n1486_1;
  assign n1516 = n2622 | n2623;
  assign n2625 = n977_1 & n1530;
  assign n2626 = N_N3829 & n1054;
  assign n1521 = n2625 | n2626;
  assign n2628 = ~N_N4060 & ~n1738;
  assign n2629 = N_N4060 & n1294;
  assign n2630 = ~n1169 & n1753;
  assign n2631 = ~n2629 & ~n2630;
  assign n1526 = ~n2628 & n2631;
  assign n2633 = NSr3_2 & ~n1914;
  assign n1531 = ~n533_1 | n2633;
  assign n2635 = NAK5_2 & n1105;
  assign n2636 = NSr5_2 & ~n2635;
  assign n1536 = ~n965 | n2636;
  assign n2638 = NAK5_2 & ~NSr5_2;
  assign n2639 = NSr5_3 & ~n2638;
  assign n1541 = ~n965 | n2639;
  assign n2641 = N_N3462 & ~n2010;
  assign n1546 = ~n2090 | n2641;
  assign n1551 = n1287 | n1546;
  assign n2644 = NAK5_2 & ~NSr5_3;
  assign n2645 = NSr5_4 & ~n2644;
  assign n1556 = ~n965 | n2645;
  assign n2647 = NDN3_8 & n1962;
  assign n2648 = NSr3_9 & ~n2647;
  assign n1561 = ~n533_1 | n2648;
  assign n2650 = NAK5_2 & ~NSr5_4;
  assign n2651 = NSr5_5 & ~n2650;
  assign n1566 = ~n965 | n2651;
  assign n2653 = NAK5_2 & ~NSr5_5;
  assign n2654 = NSr5_7 & ~n2653;
  assign n1571 = ~n965 | n2654;
  assign n2656 = NAK5_2 & ~NSr5_7;
  assign n2657 = n965 & n2656;
  assign n1576 = ~n2614 & ~n2657;
  assign n2659 = ~N_N3998 & ~n953;
  assign n2660 = ~n954 & ~n2659;
  assign n1581 = PRESET | n2660;
  always @ (posedge clock) begin
    N_N4054 <= n64_1;
    N_N3745 <= n69;
    N_N4119 <= n74_1;
    N_N3826 <= n79;
    N_N3818 <= n84_1;
    N_N3345 <= n89_1;
    N_N3924 <= n94_1;
    N_N3815 <= n99;
    N_N3691 <= n104_1;
    N_N3157 <= n109;
    N_N3872 <= n114_1;
    N_N3788 <= n119_1;
    N_N3375 <= n124_1;
    N_N3143 <= n129;
    N_N4197 <= n134;
    N_N3843 <= n139_1;
    N_N3426 <= n144_1;
    N_N4118 <= n149_1;
    N_N3580 <= n154_1;
    N_N3175 <= n159_1;
    N_N3071 <= n164_1;
    N_N3808 <= n169_1;
    N_N3923 <= n174;
    N_N3250 <= n179_1;
    N_N4221 <= n184_1;
    N_N3069 <= n189_1;
    N_N3464 <= n194_1;
    N_N3535 <= n199_1;
    N_N3871 <= n204_1;
    N_N3248 <= n209_1;
    N_N4180 <= n214_1;
    N_N3311 <= n219;
    N_N3442 <= n224_1;
    N_N3981 <= n229_1;
    N_N3842 <= n234_1;
    N_N3105 <= n239_1;
    N_N4133 <= n244_1;
    N_N4117 <= n249_1;
    N_N3420 <= n254;
    N_N3761 <= n259_1;
    N_N3062 <= n264_1;
    N_N4071 <= n269_1;
    N_N4227 <= n274;
    N_N3807 <= n279_1;
    N_N4145 <= n284;
    N_N3922 <= n289;
    N_N3516 <= n294;
    N_N3489 <= n299_1;
    N_N4030 <= n304_1;
    N_N3540 <= n309;
    N_N3513 <= n314;
    N_N4083 <= n319_1;
    N_N3841 <= n324_1;
    N_N4018 <= n329;
    N_N3971 <= n334;
    N_N4232 <= n339_1;
    N_N4246 <= n344_1;
    N_N3806 <= n349_1;
    N_N3992 <= n354;
    N_N4086 <= n359;
    N_N4230 <= n364;
    N_N4212 <= n369_1;
    Pnext_0_0_ <= n374_1;
    N_N3626 <= n378_1;
    N_N3965 <= n383_1;
    N_N3890 <= n388_1;
    NDN3_11 <= n393_1;
    NDN5_10 <= n398_1;
    N_N3786 <= n403;
    N_N4171 <= n408_1;
    NDN5_16 <= n413_1;
    N_N3799 <= n418_1;
    N_N3844 <= n423;
    N_N3196 <= n428_1;
    N_N4126 <= n433_1;
    N_N3681 <= n438;
    N_N3679 <= n443;
    N_N3340 <= n448_1;
    N_N4116 <= n453;
    N_N3810 <= n458_1;
    N_N3235 <= n463_1;
    N_N3283 <= n468;
    N_N3716 <= n473_1;
    N_N3701 <= n478_1;
    N_N3921 <= n483;
    N_N3625 <= n488;
    N_N3751 <= n493_1;
    N_N3736 <= n498;
    N_N3870 <= n503;
    N_N4024 <= n508_1;
    N_N3876 <= n513;
    N_N3840 <= n518_1;
    N_N4021 <= n523;
    N_N3932 <= n528_1;
    NLC1_2 <= n533_1;
    N_N3805 <= n538;
    N_N3700 <= n543_1;
    N_N3735 <= n548;
    NLak3_2 <= n553_1;
    NLak3_9 <= n558;
    N_N3906 <= n563_1;
    N_N3388 <= n568_1;
    N_N4057 <= n573_1;
    N_N3011 <= n578;
    N_N3346 <= n583_1;
    N_N3677 <= n588;
    N_N4165 <= n593;
    N_N4080 <= n598;
    N_N3373 <= n603;
    N_N3709 <= n608;
    N_N4206 <= n613_1;
    N_N3324 <= n618_1;
    N_N3575 <= n623_1;
    N_N4159 <= n628;
    NAK5_2 <= n633;
    N_N3916 <= n638_1;
    N_N3743 <= n643;
    N_N4242 <= n648_1;
    N_N3312 <= n653_1;
    N_N3733 <= n658;
    N_N3774 <= n663;
    N_N4214 <= n668_1;
    N_N3294 <= n673;
    N_N3796 <= n678_1;
    N_N3574 <= n683;
    N_N3791 <= n688_1;
    N_N3480 <= n693;
    N_N4243 <= n698_1;
    N_N3940 <= n703_1;
    N_N3509 <= n708;
    N_N4015 <= n713_1;
    N_N2989 <= n718;
    N_N3919 <= n723;
    N_N3578 <= n728;
    N_N3529 <= n733;
    N_N4222 <= n738;
    N_N3910 <= n743;
    N_N3868 <= n748_1;
    N_N3947 <= n753;
    N_N4181 <= n758;
    N_N3793 <= n763;
    N_N3822 <= n768;
    N_N3813 <= n773_1;
    N_N4114 <= n778_1;
    N_N4134 <= n783_1;
    N_N3866 <= n788;
    N_N4218 <= n793_1;
    N_N3939 <= n798;
    N_N3776 <= n803_1;
    N_N3387 <= n808_1;
    N_N4194 <= n813;
    N_N3821 <= n818_1;
    N_N3882 <= n823_1;
    N_N4167 <= n828_1;
    N_N3800 <= n833;
    N_N4237 <= n838_1;
    N_N3417 <= n843_1;
    N_N3918 <= n848_1;
    N_N4158 <= n853;
    N_N3630 <= n858_1;
    N_N3344 <= n863_1;
    N_N4072 <= n868;
    N_N3274 <= n873_1;
    N_N3473 <= n878_1;
    N_N4205 <= n883;
    N_N4111 <= n888_1;
    N_N3680 <= n893;
    N_N3838 <= n898;
    N_N3262 <= n903;
    N_N4099 <= n908;
    N_N3607 <= n913;
    N_N3323 <= n918_1;
    N_N3612 <= n923;
    N_N4079 <= n928;
    PDN <= n933;
    N_N3457 <= n937;
    N_N3445 <= n942;
    N_N3794 <= n947_1;
    N_N3663 <= n952;
    N_N3715 <= n957_1;
    N_N4039 <= n962_1;
    N_N3280 <= n967;
    N_N4239 <= n972;
    N_N3988 <= n977;
    N_N3433 <= n982;
    N_N4075 <= n987_1;
    N_N3468 <= n992;
    N_N4045 <= n997_1;
    N_N3482 <= n1002;
    N_N3832 <= n1007_1;
    N_N3304 <= n1012_1;
    N_N3750 <= n1017_1;
    N_N3634 <= n1022;
    N_N3293 <= n1027;
    N_N3659 <= n1032_1;
    N_N4252 <= n1037;
    N_N3912 <= n1042_1;
    N_N3862 <= n1047_1;
    N_N3221 <= n1052_1;
    N_N3875 <= n1057;
    N_N3949 <= n1062_1;
    N_N3908 <= n1067_1;
    N_N3711 <= n1072_1;
    N_N3931 <= n1077;
    N_N3469 <= n1082_1;
    N_N3436 <= n1087;
    N_N3974 <= n1092;
    N_N3905 <= n1097;
    N_N3741 <= n1102_1;
    N_N3369 <= n1107;
    N_N3164 <= n1112;
    N_N3500 <= n1117_1;
    N_N3996 <= n1122;
    N_N3356 <= n1127_1;
    N_N4093 <= n1132;
    Pover_0_0_ <= n1137;
    N_N4224 <= n1141_1;
    N_N4027 <= n1146;
    NDN1_4 <= n1151;
    N_N3384 <= n1156;
    N_N4036 <= n1161;
    N_N3968 <= n1166;
    N_N4183 <= n1171;
    NGFDN_3 <= n1176;
    N_N4090 <= n1181_1;
    N_N4004 <= n1186_1;
    N_N3205 <= n1191_1;
    N_N4136 <= n1196_1;
    N_N3303 <= n1201_1;
    N_N3533 <= n1206_1;
    N_N3336 <= n1211_1;
    N_N3961 <= n1216_1;
    N_N3331 <= n1221_1;
    N_N3203 <= n1226_1;
    N_N4236 <= n1231;
    N_N3884 <= n1236;
    N_N3367 <= n1241;
    N_N4140 <= n1246;
    NDN2_2 <= n1251;
    N_N4106 <= n1256;
    N_N3100 <= n1261;
    N_N4193 <= n1266;
    N_N3470 <= n1271_1;
    N_N3424 <= n1276_1;
    N_N3959 <= n1281;
    N_N3393 <= n1286_1;
    N_N4042 <= n1291_1;
    N_N3188 <= n1296_1;
    N_N4095 <= n1301;
    N_N3957 <= n1306;
    N_N3517 <= n1311;
    N_N4047 <= n1316;
    N_N3081 <= n1321;
    N_N3541 <= n1326;
    N_N4177 <= n1331;
    NDN3_3 <= n1336;
    N_N4176 <= n1341;
    N_N3585 <= n1346;
    NDN3_8 <= n1351;
    N_N4209 <= n1356;
    N_N3824 <= n1361;
    N_N4208 <= n1366;
    N_N4120 <= n1371;
    N_N3708 <= n1376;
    N_N4220 <= n1381;
    N_N3999 <= n1386;
    N_N4223 <= n1391;
    N_N3179 <= n1396;
    N_N4179 <= n1401;
    N_N3475 <= n1406;
    N_N4132 <= n1411;
    N_N4182 <= n1416;
    N_N3797 <= n1421;
    N_N3214 <= n1426;
    N_N4070 <= n1431;
    N_N4135 <= n1436;
    NLD3_9 <= n1441;
    NDN5_2 <= n1446;
    NDN5_3 <= n1451;
    N_N3778 <= n1456;
    NDN5_4 <= n1461;
    N_N3212 <= n1466;
    NDN5_5 <= n1471;
    NDN5_6 <= n1476;
    NDN5_7 <= n1481;
    NDN5_8 <= n1486;
    N_N4073 <= n1491;
    NDN5_9 <= n1496;
    NEN5_9 <= n1501;
    N_N3684 <= n1506;
    N_N4056 <= n1511;
    N_N3713 <= n1516;
    N_N3829 <= n1521;
    N_N4060 <= n1526;
    NSr3_2 <= n1531;
    NSr5_2 <= n1536;
    NSr5_3 <= n1541;
    N_N3462 <= n1546;
    N_N3460 <= n1551;
    NSr5_4 <= n1556;
    NSr3_9 <= n1561;
    NSr5_5 <= n1566;
    NSr5_7 <= n1571;
    NSr5_8 <= n1576;
    N_N3998 <= n1581;
  end
endmodule


