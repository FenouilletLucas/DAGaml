// Benchmark "alu4_cl" written by ABC on Tue May 16 16:07:44 2017

module alu4_cl ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    o, p, q, r, s, t, u, v  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output o, p, q, r, s, t, u, v;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
    n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n668, n669, n670, n671, n672,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996;
  assign n23 = ~a & e;
  assign n24 = i & ~k;
  assign n25 = l & n24;
  assign n26 = a & ~e;
  assign n27 = k & ~l;
  assign n28 = i & n27;
  assign n29 = ~i & ~k;
  assign n30 = k & l;
  assign n31 = ~n29 & ~n30;
  assign n32 = ~i & j;
  assign n33 = i & k;
  assign n34 = i & j;
  assign n35 = ~j & l;
  assign n36 = ~n & n35;
  assign n37 = n33 & n36;
  assign n38 = n & ~n27;
  assign n39 = n32 & n38;
  assign n40 = n27 & n34;
  assign n41 = ~n39 & ~n40;
  assign n42 = ~n37 & n41;
  assign n43 = ~n & n29;
  assign n44 = ~l & n43;
  assign n45 = ~j & n43;
  assign n46 = ~n44 & ~n45;
  assign n47 = a & e;
  assign n48 = ~i & n27;
  assign n49 = ~i & ~j;
  assign n50 = ~k & l;
  assign n51 = n34 & n50;
  assign n52 = n49 & n50;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~j & n48;
  assign n55 = n & ~n53;
  assign n56 = ~n54 & ~n55;
  assign n57 = ~k & ~l;
  assign n58 = i & ~j;
  assign n59 = ~n & n58;
  assign n60 = n57 & n59;
  assign n61 = k & n58;
  assign n62 = n & n61;
  assign n63 = ~n60 & ~n62;
  assign n64 = ~a & ~e;
  assign n65 = n & n32;
  assign n66 = n27 & n65;
  assign n67 = n23 & n66;
  assign n68 = n26 & n65;
  assign n69 = ~e & ~n42;
  assign n70 = ~a & ~n46;
  assign n71 = n47 & ~n56;
  assign n72 = ~n63 & ~n64;
  assign n73 = ~n71 & ~n72;
  assign n74 = ~n70 & n73;
  assign n75 = ~n69 & n74;
  assign n76 = ~n68 & n75;
  assign n77 = ~n67 & n76;
  assign n78 = ~i & k;
  assign n79 = i & n57;
  assign n80 = ~n78 & ~n79;
  assign n81 = a & ~n77;
  assign n82 = ~l & ~n78;
  assign n83 = ~i & l;
  assign n84 = a & l;
  assign n85 = ~k & ~n49;
  assign n86 = j & n;
  assign n87 = n83 & n86;
  assign n88 = ~k & n87;
  assign n89 = ~j & n;
  assign n90 = n28 & n89;
  assign n91 = n & n27;
  assign n92 = n47 & n91;
  assign n93 = n58 & n92;
  assign n94 = n81 & n91;
  assign n95 = n34 & n94;
  assign n96 = n77 & n91;
  assign n97 = n49 & n96;
  assign n98 = a & n87;
  assign n99 = ~n77 & n87;
  assign n100 = ~n98 & ~n99;
  assign n101 = ~n97 & n100;
  assign n102 = ~n95 & n101;
  assign n103 = ~n93 & n102;
  assign n104 = n47 & n88;
  assign n105 = n90 & n103;
  assign n106 = ~n104 & ~n105;
  assign n107 = ~j & ~l;
  assign n108 = j & n29;
  assign n109 = k & n34;
  assign n110 = ~k & n34;
  assign n111 = l & n110;
  assign n112 = j & n48;
  assign n113 = ~n111 & ~n112;
  assign n114 = n & n107;
  assign n115 = ~n77 & n114;
  assign n116 = k & n115;
  assign n117 = i & n116;
  assign n118 = n106 & n117;
  assign n119 = n77 & n114;
  assign n120 = k & n119;
  assign n121 = i & n120;
  assign n122 = ~n106 & n121;
  assign n123 = ~n103 & n114;
  assign n124 = k & n123;
  assign n125 = ~a & n124;
  assign n126 = ~i & n125;
  assign n127 = n & ~n34;
  assign n128 = n77 & n127;
  assign n129 = k & n128;
  assign n130 = l & n129;
  assign n131 = a & n130;
  assign n132 = n & n29;
  assign n133 = n77 & n132;
  assign n134 = a & n133;
  assign n135 = ~j & n134;
  assign n136 = ~n77 & n132;
  assign n137 = ~l & n136;
  assign n138 = j & n137;
  assign n139 = n & ~n77;
  assign n140 = l & n139;
  assign n141 = ~a & n140;
  assign n142 = ~n85 & n141;
  assign n143 = n & ~n103;
  assign n144 = l & n143;
  assign n145 = n108 & n144;
  assign n146 = n106 & n145;
  assign n147 = n & n103;
  assign n148 = l & n147;
  assign n149 = n108 & n148;
  assign n150 = ~n106 & n149;
  assign n151 = n103 & n114;
  assign n152 = a & n151;
  assign n153 = ~i & n152;
  assign n154 = n & n58;
  assign n155 = ~k & n154;
  assign n156 = n23 & n155;
  assign n157 = n26 & n155;
  assign n158 = l & n;
  assign n159 = ~a & n158;
  assign n160 = n109 & n159;
  assign n161 = n24 & n114;
  assign n162 = e & n161;
  assign n163 = ~l & n132;
  assign n164 = a & n163;
  assign n165 = n34 & n91;
  assign n166 = n103 & n165;
  assign n167 = n & ~n113;
  assign n168 = n77 & n167;
  assign n169 = ~n166 & ~n168;
  assign n170 = ~n164 & n169;
  assign n171 = ~n162 & n170;
  assign n172 = ~n160 & n171;
  assign n173 = ~n157 & n172;
  assign n174 = ~n156 & n173;
  assign n175 = ~n153 & n174;
  assign n176 = ~n150 & n175;
  assign n177 = ~n146 & n176;
  assign n178 = ~n142 & n177;
  assign n179 = ~n138 & n178;
  assign n180 = ~n135 & n179;
  assign n181 = ~n131 & n180;
  assign n182 = ~n126 & n181;
  assign n183 = ~n122 & n182;
  assign n184 = ~n118 & n183;
  assign n185 = ~j & k;
  assign n186 = n & n57;
  assign n187 = n34 & n186;
  assign n188 = ~n & n83;
  assign n189 = n185 & n188;
  assign n190 = ~n187 & ~n189;
  assign n191 = ~j & ~n;
  assign n192 = n25 & n191;
  assign n193 = n23 & n192;
  assign n194 = l & n191;
  assign n195 = n26 & n194;
  assign n196 = ~e & ~n;
  assign n197 = ~j & n196;
  assign n198 = n28 & n197;
  assign n199 = ~n & ~n77;
  assign n200 = ~j & n199;
  assign n201 = ~n31 & n200;
  assign n202 = ~n & n77;
  assign n203 = ~j & n202;
  assign n204 = ~n80 & n203;
  assign n205 = j & ~n;
  assign n206 = n33 & n205;
  assign n207 = n81 & n206;
  assign n208 = ~n82 & n205;
  assign n209 = n47 & n208;
  assign n210 = n64 & n205;
  assign n211 = n48 & n210;
  assign n212 = e & ~n;
  assign n213 = j & n212;
  assign n214 = n83 & n213;
  assign n215 = n43 & ~n77;
  assign n216 = e & n215;
  assign n217 = ~n & ~n85;
  assign n218 = n84 & n217;
  assign n219 = n & n184;
  assign n220 = ~m & n219;
  assign n221 = n & ~n184;
  assign n222 = m & n221;
  assign n223 = n190 & ~n222;
  assign n224 = ~n220 & n223;
  assign n225 = ~n218 & n224;
  assign n226 = ~n216 & n225;
  assign n227 = ~n214 & n226;
  assign n228 = ~n211 & n227;
  assign n229 = ~n209 & n228;
  assign n230 = ~n207 & n229;
  assign n231 = ~n204 & n230;
  assign n232 = ~n201 & n231;
  assign n233 = ~n198 & n232;
  assign n234 = ~n195 & n233;
  assign o = n193 | ~n234;
  assign n236 = ~b & f;
  assign n237 = b & ~f;
  assign n238 = ~b & ~f;
  assign n239 = b & f;
  assign n240 = ~j & n27;
  assign n241 = n & n240;
  assign n242 = n56 & ~n241;
  assign n243 = ~i & n;
  assign n244 = n27 & n243;
  assign n245 = ~n23 & n244;
  assign n246 = j & n245;
  assign n247 = n236 & n246;
  assign n248 = ~n23 & n243;
  assign n249 = j & n248;
  assign n250 = n237 & n249;
  assign n251 = n & n238;
  assign n252 = ~i & n251;
  assign n253 = n23 & n252;
  assign n254 = j & n253;
  assign n255 = n & n239;
  assign n256 = ~i & n255;
  assign n257 = n27 & n256;
  assign n258 = n23 & n257;
  assign n259 = n185 & n243;
  assign n260 = n84 & n259;
  assign n261 = ~f & ~n42;
  assign n262 = ~b & ~n46;
  assign n263 = n239 & ~n242;
  assign n264 = ~n63 & ~n238;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n262 & n265;
  assign n267 = ~n261 & n266;
  assign n268 = ~n260 & n267;
  assign n269 = ~n258 & n268;
  assign n270 = ~n254 & n269;
  assign n271 = ~n250 & n270;
  assign n272 = ~n247 & n271;
  assign n273 = b & n91;
  assign n274 = i & n273;
  assign n275 = f & n274;
  assign n276 = ~j & n275;
  assign n277 = n91 & ~n272;
  assign n278 = b & n277;
  assign n279 = i & n278;
  assign n280 = j & n279;
  assign n281 = n49 & n91;
  assign n282 = n272 & n281;
  assign n283 = n87 & ~n272;
  assign n284 = b & n87;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n282 & n285;
  assign n287 = ~n280 & n286;
  assign n288 = ~n276 & n287;
  assign n289 = n88 & n239;
  assign n290 = n90 & n288;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n77 & ~n106;
  assign n293 = ~j & n24;
  assign n294 = l & n49;
  assign n295 = n30 & ~n34;
  assign n296 = ~n294 & ~n295;
  assign n297 = ~k & n49;
  assign n298 = n296 & ~n297;
  assign n299 = ~n103 & ~n106;
  assign n300 = j & ~k;
  assign n301 = n83 & n300;
  assign n302 = a & ~n103;
  assign n303 = ~n288 & ~n302;
  assign n304 = n288 & n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~l & n32;
  assign n307 = ~n111 & ~n306;
  assign n308 = n103 & n288;
  assign n309 = ~a & ~b;
  assign n310 = ~n34 & n57;
  assign n311 = n77 & n272;
  assign n312 = n114 & ~n272;
  assign n313 = n33 & n312;
  assign n314 = ~n292 & n313;
  assign n315 = n291 & n314;
  assign n316 = n114 & n272;
  assign n317 = n33 & n316;
  assign n318 = n292 & n317;
  assign n319 = n291 & n318;
  assign n320 = ~n292 & n317;
  assign n321 = ~n291 & n320;
  assign n322 = n292 & n313;
  assign n323 = ~n291 & n322;
  assign n324 = n & n293;
  assign n325 = l & n324;
  assign n326 = n47 & n325;
  assign n327 = n238 & n326;
  assign n328 = b & n324;
  assign n329 = ~f & n328;
  assign n330 = ~n47 & n329;
  assign n331 = n & n272;
  assign n332 = ~n81 & n331;
  assign n333 = b & n332;
  assign n334 = ~n298 & n333;
  assign n335 = n & ~n272;
  assign n336 = n81 & n335;
  assign n337 = b & n336;
  assign n338 = ~n298 & n337;
  assign n339 = n & n301;
  assign n340 = ~n288 & n339;
  assign n341 = n291 & n340;
  assign n342 = ~n299 & n341;
  assign n343 = n288 & n339;
  assign n344 = ~n291 & n343;
  assign n345 = ~n299 & n344;
  assign n346 = n291 & n343;
  assign n347 = n299 & n346;
  assign n348 = ~n291 & n340;
  assign n349 = n299 & n348;
  assign n350 = n & n109;
  assign n351 = ~l & n350;
  assign n352 = ~n103 & n351;
  assign n353 = ~n288 & n352;
  assign n354 = b & n114;
  assign n355 = n305 & n354;
  assign n356 = ~i & n355;
  assign n357 = ~b & n114;
  assign n358 = ~n305 & n357;
  assign n359 = n78 & n358;
  assign n360 = n & ~n296;
  assign n361 = ~n272 & n360;
  assign n362 = ~n81 & n361;
  assign n363 = ~b & n362;
  assign n364 = n272 & n360;
  assign n365 = n81 & n364;
  assign n366 = ~b & n365;
  assign n367 = n47 & n324;
  assign n368 = n239 & n367;
  assign n369 = ~n47 & n324;
  assign n370 = n236 & n369;
  assign n371 = ~n307 & n335;
  assign n372 = ~n77 & n371;
  assign n373 = ~l & n335;
  assign n374 = n108 & n373;
  assign n375 = b & n350;
  assign n376 = n84 & n375;
  assign n377 = n308 & n351;
  assign n378 = n309 & n350;
  assign n379 = l & n378;
  assign n380 = f & n161;
  assign n381 = b & n;
  assign n382 = n310 & n381;
  assign n383 = n167 & n311;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n380 & n384;
  assign n386 = ~n379 & n385;
  assign n387 = ~n377 & n386;
  assign n388 = ~n376 & n387;
  assign n389 = ~n374 & n388;
  assign n390 = ~n372 & n389;
  assign n391 = ~n370 & n390;
  assign n392 = ~n368 & n391;
  assign n393 = ~n366 & n392;
  assign n394 = ~n363 & n393;
  assign n395 = ~n359 & n394;
  assign n396 = ~n356 & n395;
  assign n397 = ~n353 & n396;
  assign n398 = ~n349 & n397;
  assign n399 = ~n347 & n398;
  assign n400 = ~n345 & n399;
  assign n401 = ~n342 & n400;
  assign n402 = ~n338 & n401;
  assign n403 = ~n334 & n402;
  assign n404 = ~n330 & n403;
  assign n405 = ~n327 & n404;
  assign n406 = ~n323 & n405;
  assign n407 = ~n321 & n406;
  assign n408 = ~n319 & n407;
  assign n409 = ~n315 & n408;
  assign n410 = ~m & ~n184;
  assign n411 = ~n & ~n272;
  assign n412 = b & n411;
  assign n413 = j & n412;
  assign n414 = n33 & n413;
  assign n415 = n208 & n239;
  assign n416 = n48 & n205;
  assign n417 = n238 & n416;
  assign n418 = f & ~n;
  assign n419 = j & n418;
  assign n420 = n83 & n419;
  assign n421 = n192 & n236;
  assign n422 = n194 & n237;
  assign n423 = ~f & ~n;
  assign n424 = ~j & n423;
  assign n425 = n28 & n424;
  assign n426 = ~j & n411;
  assign n427 = ~n31 & n426;
  assign n428 = ~n & n272;
  assign n429 = ~j & n428;
  assign n430 = ~n80 & n429;
  assign n431 = b & n217;
  assign n432 = l & n431;
  assign n433 = n43 & ~n272;
  assign n434 = f & n433;
  assign n435 = n & n410;
  assign n436 = n409 & n435;
  assign n437 = n & ~n410;
  assign n438 = ~n409 & n437;
  assign n439 = n190 & ~n438;
  assign n440 = ~n436 & n439;
  assign n441 = ~n434 & n440;
  assign n442 = ~n432 & n441;
  assign n443 = ~n430 & n442;
  assign n444 = ~n427 & n443;
  assign n445 = ~n425 & n444;
  assign n446 = ~n422 & n445;
  assign n447 = ~n421 & n446;
  assign n448 = ~n420 & n447;
  assign n449 = ~n417 & n448;
  assign n450 = ~n415 & n449;
  assign p = n414 | ~n450;
  assign n452 = n23 & ~n237;
  assign n453 = ~n236 & ~n452;
  assign n454 = ~c & ~g;
  assign n455 = c & g;
  assign n456 = ~c & g;
  assign n457 = n & n456;
  assign n458 = ~i & n457;
  assign n459 = n27 & n458;
  assign n460 = n453 & n459;
  assign n461 = j & n460;
  assign n462 = c & ~g;
  assign n463 = n & n462;
  assign n464 = ~i & n463;
  assign n465 = n453 & n464;
  assign n466 = j & n465;
  assign n467 = n & n454;
  assign n468 = ~i & n467;
  assign n469 = ~n453 & n468;
  assign n470 = j & n469;
  assign n471 = n & n455;
  assign n472 = ~i & n471;
  assign n473 = n27 & n472;
  assign n474 = ~n453 & n473;
  assign n475 = b & n259;
  assign n476 = l & n475;
  assign n477 = ~g & ~n42;
  assign n478 = ~c & ~n46;
  assign n479 = ~n63 & ~n454;
  assign n480 = ~n242 & n455;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n478 & n481;
  assign n483 = ~n477 & n482;
  assign n484 = ~n476 & n483;
  assign n485 = ~n474 & n484;
  assign n486 = ~n470 & n485;
  assign n487 = ~n466 & n486;
  assign n488 = ~n461 & n487;
  assign n489 = c & l;
  assign n490 = n47 & ~n238;
  assign n491 = ~n239 & ~n490;
  assign n492 = c & n91;
  assign n493 = i & n492;
  assign n494 = g & n493;
  assign n495 = ~j & n494;
  assign n496 = n91 & ~n488;
  assign n497 = c & n496;
  assign n498 = i & n497;
  assign n499 = j & n498;
  assign n500 = n281 & n488;
  assign n501 = n87 & ~n488;
  assign n502 = c & n87;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n500 & n503;
  assign n505 = ~n499 & n504;
  assign n506 = ~n495 & n505;
  assign n507 = b & n302;
  assign n508 = b & ~n288;
  assign n509 = ~n288 & n302;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n507 & n510;
  assign n512 = n506 & ~n511;
  assign n513 = ~n506 & n511;
  assign n514 = ~n512 & ~n513;
  assign n515 = b & n81;
  assign n516 = b & ~n272;
  assign n517 = n81 & ~n272;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n515 & n518;
  assign n520 = ~n291 & n292;
  assign n521 = ~n272 & n292;
  assign n522 = ~n272 & ~n291;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n520 & n523;
  assign n525 = n88 & n455;
  assign n526 = n90 & n506;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~n488 & ~n527;
  assign n529 = n488 & n527;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n291 & n299;
  assign n532 = ~n288 & n299;
  assign n533 = ~n288 & ~n291;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n531 & n534;
  assign n536 = n308 & n506;
  assign n537 = ~c & n309;
  assign n538 = n311 & n488;
  assign n539 = n324 & ~n491;
  assign n540 = l & n539;
  assign n541 = n454 & n540;
  assign n542 = n350 & ~n506;
  assign n543 = ~l & n542;
  assign n544 = ~n308 & n543;
  assign n545 = ~c & n114;
  assign n546 = ~n514 & n545;
  assign n547 = n78 & n546;
  assign n548 = n & ~n488;
  assign n549 = ~c & n548;
  assign n550 = n519 & n549;
  assign n551 = ~n296 & n550;
  assign n552 = n & n488;
  assign n553 = ~c & n552;
  assign n554 = ~n519 & n553;
  assign n555 = ~n296 & n554;
  assign n556 = c & n552;
  assign n557 = ~n298 & n556;
  assign n558 = n519 & n557;
  assign n559 = c & n548;
  assign n560 = ~n298 & n559;
  assign n561 = ~n519 & n560;
  assign n562 = c & n114;
  assign n563 = n514 & n562;
  assign n564 = ~i & n563;
  assign n565 = n33 & n114;
  assign n566 = n530 & n565;
  assign n567 = n524 & n566;
  assign n568 = ~n530 & n565;
  assign n569 = ~n524 & n568;
  assign n570 = n324 & n491;
  assign n571 = c & n570;
  assign n572 = ~g & n571;
  assign n573 = ~c & n570;
  assign n574 = g & n573;
  assign n575 = n339 & ~n527;
  assign n576 = n506 & n575;
  assign n577 = n535 & n576;
  assign n578 = n339 & n527;
  assign n579 = ~n506 & n578;
  assign n580 = n535 & n579;
  assign n581 = n506 & n578;
  assign n582 = ~n535 & n581;
  assign n583 = ~n506 & n575;
  assign n584 = ~n535 & n583;
  assign n585 = n455 & n539;
  assign n586 = ~n307 & n548;
  assign n587 = ~n311 & n586;
  assign n588 = ~l & n548;
  assign n589 = n108 & n588;
  assign n590 = n351 & n536;
  assign n591 = n350 & n537;
  assign n592 = l & n591;
  assign n593 = n350 & n489;
  assign n594 = ~n309 & n593;
  assign n595 = g & n161;
  assign n596 = c & n;
  assign n597 = n310 & n596;
  assign n598 = n167 & n538;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n595 & n599;
  assign n601 = ~n594 & n600;
  assign n602 = ~n592 & n601;
  assign n603 = ~n590 & n602;
  assign n604 = ~n589 & n603;
  assign n605 = ~n587 & n604;
  assign n606 = ~n585 & n605;
  assign n607 = ~n584 & n606;
  assign n608 = ~n582 & n607;
  assign n609 = ~n580 & n608;
  assign n610 = ~n577 & n609;
  assign n611 = ~n574 & n610;
  assign n612 = ~n572 & n611;
  assign n613 = ~n569 & n612;
  assign n614 = ~n567 & n613;
  assign n615 = ~n564 & n614;
  assign n616 = ~n561 & n615;
  assign n617 = ~n558 & n616;
  assign n618 = ~n555 & n617;
  assign n619 = ~n551 & n618;
  assign n620 = ~n547 & n619;
  assign n621 = ~n544 & n620;
  assign n622 = ~n541 & n621;
  assign n623 = ~n409 & n410;
  assign n624 = g & ~n;
  assign n625 = ~j & n624;
  assign n626 = ~c & n625;
  assign n627 = n25 & n626;
  assign n628 = ~n & ~n488;
  assign n629 = j & n628;
  assign n630 = n33 & n629;
  assign n631 = c & n630;
  assign n632 = ~g & ~n;
  assign n633 = ~j & n632;
  assign n634 = n28 & n633;
  assign n635 = ~n & n488;
  assign n636 = ~j & n635;
  assign n637 = ~n80 & n636;
  assign n638 = ~j & n628;
  assign n639 = ~n31 & n638;
  assign n640 = n205 & n454;
  assign n641 = n48 & n640;
  assign n642 = j & n624;
  assign n643 = n83 & n642;
  assign n644 = n208 & n455;
  assign n645 = ~n & n489;
  assign n646 = ~g & n645;
  assign n647 = ~j & n646;
  assign n648 = n43 & ~n488;
  assign n649 = g & n648;
  assign n650 = n217 & n489;
  assign n651 = n & n623;
  assign n652 = n622 & n651;
  assign n653 = n & ~n623;
  assign n654 = ~n622 & n653;
  assign n655 = n190 & ~n654;
  assign n656 = ~n652 & n655;
  assign n657 = ~n650 & n656;
  assign n658 = ~n649 & n657;
  assign n659 = ~n647 & n658;
  assign n660 = ~n644 & n659;
  assign n661 = ~n643 & n660;
  assign n662 = ~n641 & n661;
  assign n663 = ~n639 & n662;
  assign n664 = ~n637 & n663;
  assign n665 = ~n634 & n664;
  assign n666 = ~n631 & n665;
  assign q = n627 | ~n666;
  assign n668 = c & n453;
  assign n669 = ~g & n453;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~n462 & n670;
  assign n672 = ~d & ~h;
  assign t = d & h;
  assign n674 = h & n;
  assign n675 = ~i & n674;
  assign n676 = ~d & n675;
  assign n677 = ~n671 & n676;
  assign n678 = n27 & n677;
  assign n679 = j & n678;
  assign n680 = ~h & n;
  assign n681 = ~i & n680;
  assign n682 = d & n681;
  assign n683 = ~n671 & n682;
  assign n684 = j & n683;
  assign n685 = ~i & ~n;
  assign n686 = ~d & n685;
  assign n687 = ~k & n686;
  assign n688 = ~l & n687;
  assign n689 = ~j & n687;
  assign n690 = n & n672;
  assign n691 = ~i & n690;
  assign n692 = n671 & n691;
  assign n693 = j & n692;
  assign n694 = n & t;
  assign n695 = ~i & n694;
  assign n696 = n671 & n695;
  assign n697 = n27 & n696;
  assign n698 = n243 & n489;
  assign n699 = n185 & n698;
  assign n700 = ~n53 & n694;
  assign n701 = ~i & t;
  assign n702 = n240 & n701;
  assign n703 = n240 & n694;
  assign n704 = ~h & ~n42;
  assign n705 = ~n63 & ~n672;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n703 & n706;
  assign n708 = ~n702 & n707;
  assign n709 = ~n700 & n708;
  assign n710 = ~n699 & n709;
  assign n711 = ~n697 & n710;
  assign n712 = ~n693 & n711;
  assign n713 = ~n689 & n712;
  assign n714 = ~n688 & n713;
  assign n715 = ~n684 & n714;
  assign n716 = ~n679 & n715;
  assign n717 = d & ~n716;
  assign n718 = d & l;
  assign n719 = c & ~n511;
  assign n720 = c & ~n506;
  assign n721 = ~n506 & ~n511;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~n719 & n722;
  assign n724 = n91 & t;
  assign n725 = n58 & n724;
  assign n726 = n91 & n717;
  assign n727 = n34 & n726;
  assign n728 = n91 & n716;
  assign n729 = n49 & n728;
  assign n730 = d & n87;
  assign n731 = n87 & ~n716;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n729 & n732;
  assign n734 = ~n727 & n733;
  assign n735 = ~n725 & n734;
  assign n736 = ~n527 & ~n535;
  assign n737 = ~n506 & ~n535;
  assign n738 = ~n506 & ~n527;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = n88 & t;
  assign n742 = n90 & n735;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n454 & ~n491;
  assign n745 = ~n455 & ~n744;
  assign n746 = ~n524 & ~n527;
  assign n747 = ~n488 & ~n524;
  assign n748 = ~n528 & ~n747;
  assign n749 = ~n746 & n748;
  assign n750 = n716 & ~n743;
  assign n751 = ~n716 & n743;
  assign n752 = ~n750 & ~n751;
  assign n753 = c & ~n519;
  assign n754 = c & ~n488;
  assign n755 = ~n488 & ~n519;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n753 & n756;
  assign n758 = n716 & ~n757;
  assign n759 = ~n716 & n757;
  assign n760 = ~n758 & ~n759;
  assign n761 = n538 & n716;
  assign n762 = d & n;
  assign n763 = ~l & n762;
  assign n764 = n735 & n763;
  assign n765 = n723 & n764;
  assign n766 = n49 & n765;
  assign n767 = ~n735 & n763;
  assign n768 = ~n723 & n767;
  assign n769 = n49 & n768;
  assign n770 = ~d & n241;
  assign n771 = ~i & n770;
  assign n772 = ~n735 & n771;
  assign n773 = n723 & n772;
  assign n774 = n735 & n771;
  assign n775 = ~n723 & n774;
  assign n776 = n & n108;
  assign n777 = l & n776;
  assign n778 = ~n743 & n777;
  assign n779 = n735 & n778;
  assign n780 = n740 & n779;
  assign n781 = n743 & n777;
  assign n782 = ~n735 & n781;
  assign n783 = n740 & n782;
  assign n784 = n735 & n781;
  assign n785 = ~n740 & n784;
  assign n786 = ~n735 & n778;
  assign n787 = ~n740 & n786;
  assign n788 = n325 & ~n745;
  assign n789 = n672 & n788;
  assign n790 = i & n241;
  assign n791 = ~n752 & n790;
  assign n792 = n749 & n791;
  assign n793 = n752 & n790;
  assign n794 = ~n749 & n793;
  assign n795 = n351 & ~n735;
  assign n796 = ~n536 & n795;
  assign n797 = n351 & n735;
  assign n798 = n536 & n797;
  assign n799 = d & n324;
  assign n800 = n745 & n799;
  assign n801 = ~h & n800;
  assign n802 = ~d & n324;
  assign n803 = n745 & n802;
  assign n804 = h & n803;
  assign n805 = ~d & n591;
  assign n806 = l & n805;
  assign n807 = n324 & ~n745;
  assign n808 = t & n807;
  assign n809 = n760 & n762;
  assign n810 = ~n298 & n809;
  assign n811 = ~l & n324;
  assign n812 = h & n811;
  assign n813 = ~d & n;
  assign n814 = ~n760 & n813;
  assign n815 = ~n296 & n814;
  assign n816 = ~n716 & n776;
  assign n817 = ~l & n816;
  assign n818 = n350 & n718;
  assign n819 = ~n537 & n818;
  assign n820 = n & ~n307;
  assign n821 = ~n716 & n820;
  assign n822 = ~n538 & n821;
  assign n823 = n310 & n762;
  assign n824 = n167 & n761;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n822 & n825;
  assign n827 = ~n819 & n826;
  assign n828 = ~n817 & n827;
  assign n829 = ~n815 & n828;
  assign n830 = ~n812 & n829;
  assign n831 = ~n810 & n830;
  assign n832 = ~n808 & n831;
  assign n833 = ~n806 & n832;
  assign n834 = ~n804 & n833;
  assign n835 = ~n801 & n834;
  assign n836 = ~n798 & n835;
  assign n837 = ~n796 & n836;
  assign n838 = ~n794 & n837;
  assign n839 = ~n792 & n838;
  assign n840 = ~n789 & n839;
  assign n841 = ~n787 & n840;
  assign n842 = ~n785 & n841;
  assign n843 = ~n783 & n842;
  assign n844 = ~n780 & n843;
  assign n845 = ~n775 & n844;
  assign n846 = ~n773 & n845;
  assign n847 = ~n769 & n846;
  assign n848 = ~n766 & n847;
  assign n849 = ~n622 & n623;
  assign n850 = h & ~n;
  assign n851 = ~j & n850;
  assign n852 = n25 & n851;
  assign n853 = ~d & n852;
  assign n854 = ~h & ~n;
  assign n855 = ~j & n854;
  assign n856 = n28 & n855;
  assign n857 = ~n & n716;
  assign n858 = ~j & n857;
  assign n859 = ~n80 & n858;
  assign n860 = ~n & ~n716;
  assign n861 = ~j & n860;
  assign n862 = ~n31 & n861;
  assign n863 = n208 & t;
  assign n864 = n416 & n672;
  assign n865 = n206 & n717;
  assign n866 = j & n850;
  assign n867 = n83 & n866;
  assign n868 = ~n & n718;
  assign n869 = ~h & n868;
  assign n870 = ~j & n869;
  assign n871 = n43 & ~n716;
  assign n872 = h & n871;
  assign n873 = n217 & n718;
  assign n874 = n & n849;
  assign n875 = n848 & n874;
  assign n876 = n & ~n849;
  assign n877 = ~n848 & n876;
  assign n878 = n190 & ~n877;
  assign n879 = ~n875 & n878;
  assign n880 = ~n873 & n879;
  assign n881 = ~n872 & n880;
  assign n882 = ~n870 & n881;
  assign n883 = ~n867 & n882;
  assign n884 = ~n865 & n883;
  assign n885 = ~n864 & n884;
  assign n886 = ~n863 & n885;
  assign n887 = ~n862 & n886;
  assign n888 = ~n859 & n887;
  assign n889 = ~n856 & n888;
  assign r = n853 | ~n889;
  assign s = n672 | t;
  assign n892 = ~l & n;
  assign n893 = n185 & n892;
  assign n894 = i & n893;
  assign n895 = ~n716 & n894;
  assign n896 = ~n749 & n895;
  assign n897 = ~n743 & n894;
  assign n898 = ~n749 & n897;
  assign n899 = ~n34 & n158;
  assign n900 = k & n899;
  assign n901 = ~n757 & n900;
  assign n902 = ~n716 & n901;
  assign n903 = ~n716 & n897;
  assign n904 = ~i & n893;
  assign n905 = d & n904;
  assign n906 = ~n723 & n905;
  assign n907 = ~n735 & n893;
  assign n908 = ~i & n907;
  assign n909 = ~n723 & n908;
  assign n910 = d & n900;
  assign n911 = ~n757 & n910;
  assign n912 = d & n908;
  assign n913 = n158 & ~n757;
  assign n914 = n49 & n913;
  assign n915 = ~n716 & n914;
  assign n916 = d & n158;
  assign n917 = ~n757 & n916;
  assign n918 = n49 & n917;
  assign n919 = n158 & n293;
  assign n920 = ~n672 & n919;
  assign n921 = ~n745 & n920;
  assign n922 = n717 & n900;
  assign n923 = n108 & n158;
  assign n924 = ~n743 & n923;
  assign n925 = ~n740 & n924;
  assign n926 = n158 & ~n735;
  assign n927 = n108 & n926;
  assign n928 = ~n740 & n927;
  assign n929 = ~n743 & n927;
  assign n930 = n109 & n158;
  assign n931 = n537 & n930;
  assign n932 = ~d & n931;
  assign n933 = n & n761;
  assign n934 = ~l & n933;
  assign n935 = n32 & n934;
  assign n936 = k & n935;
  assign n937 = n34 & n892;
  assign n938 = n735 & n937;
  assign n939 = n536 & n938;
  assign n940 = n158 & n717;
  assign n941 = n49 & n940;
  assign n942 = t & n919;
  assign n943 = n & n110;
  assign n944 = ~l & n943;
  assign n945 = ~n848 & n874;
  assign n946 = n110 & n933;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~n944 & n947;
  assign n949 = ~n942 & n948;
  assign n950 = ~n941 & n949;
  assign n951 = ~n939 & n950;
  assign n952 = ~n936 & n951;
  assign n953 = ~n932 & n952;
  assign n954 = ~n929 & n953;
  assign n955 = ~n928 & n954;
  assign n956 = ~n925 & n955;
  assign n957 = ~n922 & n956;
  assign n958 = ~n921 & n957;
  assign n959 = ~n918 & n958;
  assign n960 = ~n915 & n959;
  assign n961 = ~n912 & n960;
  assign n962 = ~n911 & n961;
  assign n963 = ~n909 & n962;
  assign n964 = ~n906 & n963;
  assign n965 = ~n903 & n964;
  assign n966 = ~n902 & n965;
  assign n967 = ~n898 & n966;
  assign u = n896 | ~n967;
  assign n969 = ~e & s;
  assign n970 = ~f & n969;
  assign n971 = n537 & n970;
  assign n972 = ~g & n971;
  assign n973 = n455 & n970;
  assign n974 = n309 & n973;
  assign n975 = n47 & s;
  assign n976 = n238 & n975;
  assign n977 = n454 & n976;
  assign n978 = n239 & s;
  assign n979 = n47 & n978;
  assign n980 = n454 & n979;
  assign n981 = n64 & s;
  assign n982 = n239 & n981;
  assign n983 = n454 & n982;
  assign n984 = n455 & s;
  assign n985 = n47 & n984;
  assign n986 = n238 & n985;
  assign n987 = n239 & n984;
  assign n988 = n47 & n987;
  assign n989 = n64 & n984;
  assign n990 = n239 & n989;
  assign n991 = ~n988 & ~n990;
  assign n992 = ~n986 & n991;
  assign n993 = ~n983 & n992;
  assign n994 = ~n980 & n993;
  assign n995 = ~n977 & n994;
  assign n996 = ~n974 & n995;
  assign v = n972 | ~n996;
endmodule


