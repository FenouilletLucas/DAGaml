// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:10 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_;
  wire n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
    n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
    n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
    n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
    n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
  assign n21 = ~i_0_ & ~i_1_;
  assign n22 = i_2_ & n21;
  assign n23 = ~i_9_ & n22;
  assign n24 = ~i_6_ & ~i_7_;
  assign n25 = i_8_ & n24;
  assign n26 = ~i_3_ & i_4_;
  assign n27 = ~i_5_ & n26;
  assign n28 = n25 & n27;
  assign n29 = n23 & n28;
  assign n30 = ~i_6_ & i_7_;
  assign n31 = i_8_ & n30;
  assign n32 = i_9_ & n31;
  assign n33 = ~i_0_ & i_1_;
  assign n34 = ~i_2_ & n33;
  assign n35 = ~i_3_ & ~i_4_;
  assign n36 = ~i_5_ & n35;
  assign n37 = n34 & n36;
  assign n38 = n32 & n37;
  assign n39 = ~n29 & ~n38;
  assign n40 = ~i_2_ & n21;
  assign n41 = ~i_9_ & n40;
  assign n42 = ~i_8_ & n24;
  assign n43 = i_3_ & i_4_;
  assign n44 = ~i_5_ & n43;
  assign n45 = n42 & n44;
  assign n46 = i_5_ & n35;
  assign n47 = i_6_ & i_7_;
  assign n48 = i_8_ & n47;
  assign n49 = n46 & n48;
  assign n50 = ~n45 & ~n49;
  assign n51 = n41 & ~n50;
  assign n52 = i_0_ & ~i_1_;
  assign n53 = ~i_9_ & n52;
  assign n54 = i_2_ & n53;
  assign n55 = i_5_ & n26;
  assign n56 = n48 & n55;
  assign n57 = n54 & n56;
  assign n58 = ~i_9_ & n34;
  assign n59 = ~i_8_ & n30;
  assign n60 = n36 & n59;
  assign n61 = n58 & n60;
  assign n62 = ~n57 & ~n61;
  assign n63 = ~n51 & n62;
  assign n64 = i_0_ & i_1_;
  assign n65 = ~i_9_ & n64;
  assign n66 = i_2_ & n65;
  assign n67 = ~i_8_ & n47;
  assign n68 = n55 & n67;
  assign n69 = n25 & n36;
  assign n70 = ~n68 & ~n69;
  assign n71 = n66 & ~n70;
  assign n72 = i_9_ & n59;
  assign n73 = i_2_ & n52;
  assign n74 = i_5_ & n43;
  assign n75 = n73 & n74;
  assign n76 = n72 & n75;
  assign n77 = i_6_ & ~i_7_;
  assign n78 = i_9_ & n77;
  assign n79 = ~i_8_ & n78;
  assign n80 = n22 & n46;
  assign n81 = n79 & n80;
  assign n82 = ~n76 & ~n81;
  assign n83 = ~n71 & n82;
  assign n84 = n63 & n83;
  assign n85 = n39 & n84;
  assign n86 = ~i_2_ & n52;
  assign n87 = n55 & n86;
  assign n88 = n79 & n87;
  assign n89 = i_9_ & n48;
  assign n90 = n46 & n86;
  assign n91 = n89 & n90;
  assign n92 = ~n88 & ~n91;
  assign n93 = ~i_2_ & n64;
  assign n94 = n74 & n93;
  assign n95 = i_9_ & n67;
  assign n96 = ~n72 & ~n95;
  assign n97 = n94 & ~n96;
  assign n98 = i_8_ & n77;
  assign n99 = i_9_ & n98;
  assign n100 = n34 & n74;
  assign n101 = n99 & n100;
  assign n102 = i_9_ & n25;
  assign n103 = n36 & n73;
  assign n104 = n102 & n103;
  assign n105 = ~n101 & ~n104;
  assign n106 = ~n97 & n105;
  assign n107 = n92 & n106;
  assign n108 = n85 & n107;
  assign n109 = n27 & n30;
  assign n110 = i_8_ & n109;
  assign n111 = n41 & n110;
  assign n112 = n42 & n55;
  assign n113 = i_2_ & n33;
  assign n114 = ~i_9_ & n113;
  assign n115 = n112 & n114;
  assign n116 = ~n111 & ~n115;
  assign n117 = ~i_2_ & n53;
  assign n118 = n26 & n98;
  assign n119 = i_5_ & n118;
  assign n120 = n117 & n119;
  assign n121 = n25 & n46;
  assign n122 = ~i_2_ & n65;
  assign n123 = n121 & n122;
  assign n124 = i_3_ & ~i_4_;
  assign n125 = i_5_ & n124;
  assign n126 = n59 & n125;
  assign n127 = n54 & n126;
  assign n128 = ~n123 & ~n127;
  assign n129 = ~n120 & n128;
  assign n130 = n46 & n73;
  assign n131 = n32 & n130;
  assign n132 = n54 & n112;
  assign n133 = ~n131 & ~n132;
  assign n134 = n34 & n55;
  assign n135 = n99 & n134;
  assign n136 = n133 & ~n135;
  assign n137 = n129 & n136;
  assign n138 = n116 & n137;
  assign n139 = n44 & n48;
  assign n140 = n30 & n55;
  assign n141 = n25 & n55;
  assign n142 = ~n140 & ~n141;
  assign n143 = ~n139 & n142;
  assign n144 = n54 & ~n143;
  assign n145 = ~i_5_ & n124;
  assign n146 = n86 & n145;
  assign n147 = n22 & n145;
  assign n148 = ~n146 & ~n147;
  assign n149 = n79 & ~n148;
  assign n150 = n34 & n44;
  assign n151 = n32 & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = n27 & n34;
  assign n154 = n72 & n153;
  assign n155 = ~i_5_ & n118;
  assign n156 = n41 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = n152 & n157;
  assign n159 = ~n144 & n158;
  assign n160 = n138 & n159;
  assign n161 = n108 & n160;
  assign n162 = n55 & n113;
  assign n163 = ~n95 & ~n99;
  assign n164 = n162 & ~n163;
  assign n165 = n43 & n113;
  assign n166 = i_5_ & n165;
  assign n167 = n79 & n166;
  assign n168 = n30 & n145;
  assign n169 = ~i_8_ & n168;
  assign n170 = n58 & n169;
  assign n171 = n55 & n59;
  assign n172 = n23 & n171;
  assign n173 = ~n170 & ~n172;
  assign n174 = ~n167 & n173;
  assign n175 = n46 & n113;
  assign n176 = n32 & n175;
  assign n177 = n40 & n55;
  assign n178 = n102 & n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = n44 & n93;
  assign n181 = n99 & n180;
  assign n182 = n179 & ~n181;
  assign n183 = ~i_8_ & n77;
  assign n184 = n125 & n183;
  assign n185 = ~n121 & ~n184;
  assign n186 = n117 & ~n185;
  assign n187 = n34 & n145;
  assign n188 = n72 & n187;
  assign n189 = ~n186 & ~n188;
  assign n190 = n182 & n189;
  assign n191 = n174 & n190;
  assign n192 = ~n164 & n191;
  assign n193 = n161 & n192;
  assign n194 = n47 & n125;
  assign n195 = i_8_ & n194;
  assign n196 = n54 & n195;
  assign n197 = n22 & n27;
  assign n198 = n79 & n197;
  assign n199 = n98 & n125;
  assign n200 = n23 & n199;
  assign n201 = ~n198 & ~n200;
  assign n202 = ~n196 & n201;
  assign n203 = i_9_ & n42;
  assign n204 = n113 & n125;
  assign n205 = n203 & n204;
  assign n206 = n202 & ~n205;
  assign n207 = n55 & n183;
  assign n208 = n48 & n74;
  assign n209 = ~n207 & ~n208;
  assign n210 = n114 & ~n209;
  assign n211 = n22 & n44;
  assign n212 = n99 & n211;
  assign n213 = n36 & n67;
  assign n214 = n58 & n213;
  assign n215 = ~n212 & ~n214;
  assign n216 = ~n210 & n215;
  assign n217 = n206 & n216;
  assign n218 = n74 & n183;
  assign n219 = n117 & n218;
  assign n220 = n27 & n183;
  assign n221 = n66 & n220;
  assign n222 = ~n219 & ~n221;
  assign n223 = n25 & n74;
  assign n224 = n54 & n223;
  assign n225 = n67 & n74;
  assign n226 = n41 & n225;
  assign n227 = ~n224 & ~n226;
  assign n228 = n222 & n227;
  assign n229 = n36 & n77;
  assign n230 = ~i_8_ & n229;
  assign n231 = n122 & n230;
  assign n232 = n40 & n145;
  assign n233 = n72 & n232;
  assign n234 = n78 & n130;
  assign n235 = n55 & n73;
  assign n236 = n203 & n235;
  assign n237 = ~n234 & ~n236;
  assign n238 = ~n233 & n237;
  assign n239 = ~n231 & n238;
  assign n240 = n228 & n239;
  assign n241 = n217 & n240;
  assign n242 = n46 & n67;
  assign n243 = n27 & n67;
  assign n244 = ~n242 & ~n243;
  assign n245 = n122 & ~n244;
  assign n246 = n86 & n125;
  assign n247 = n102 & n246;
  assign n248 = ~n245 & ~n247;
  assign n249 = i_2_ & n64;
  assign n250 = n44 & n249;
  assign n251 = n72 & n250;
  assign n252 = n79 & n232;
  assign n253 = ~n251 & ~n252;
  assign n254 = n32 & n90;
  assign n255 = n30 & n125;
  assign n256 = n23 & n255;
  assign n257 = ~n254 & ~n256;
  assign n258 = n253 & n257;
  assign n259 = n248 & n258;
  assign n260 = i_8_ & n229;
  assign n261 = n122 & n260;
  assign n262 = n32 & n211;
  assign n263 = ~n261 & ~n262;
  assign n264 = n27 & n73;
  assign n265 = n34 & n125;
  assign n266 = ~n264 & ~n265;
  assign n267 = n32 & ~n266;
  assign n268 = n58 & n68;
  assign n269 = ~n267 & ~n268;
  assign n270 = n263 & n269;
  assign n271 = n259 & n270;
  assign n272 = ~n195 & ~n208;
  assign n273 = n122 & ~n272;
  assign n274 = n89 & n264;
  assign n275 = n22 & n242;
  assign n276 = ~n274 & ~n275;
  assign n277 = ~n273 & n276;
  assign n278 = n25 & n44;
  assign n279 = ~n243 & ~n278;
  assign n280 = n54 & ~n279;
  assign n281 = ~n117 & ~n122;
  assign n282 = n45 & ~n281;
  assign n283 = n102 & n130;
  assign n284 = ~n282 & ~n283;
  assign n285 = ~n280 & n284;
  assign n286 = n277 & n285;
  assign n287 = n271 & n286;
  assign n288 = n241 & n287;
  assign n289 = n193 & n288;
  assign n290 = n117 & n230;
  assign n291 = n75 & n99;
  assign n292 = n32 & n197;
  assign n293 = n46 & n59;
  assign n294 = n114 & n293;
  assign n295 = ~n292 & ~n294;
  assign n296 = ~n291 & n295;
  assign n297 = ~n290 & n296;
  assign n298 = n23 & n155;
  assign n299 = n44 & n86;
  assign n300 = n79 & n299;
  assign n301 = n58 & n171;
  assign n302 = ~n300 & ~n301;
  assign n303 = ~n298 & n302;
  assign n304 = n113 & n145;
  assign n305 = n36 & n113;
  assign n306 = n93 & n145;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~n304 & n307;
  assign n309 = n89 & ~n308;
  assign n310 = n303 & ~n309;
  assign n311 = n297 & n310;
  assign n312 = n203 & n304;
  assign n313 = n122 & n223;
  assign n314 = n44 & n59;
  assign n315 = n41 & n314;
  assign n316 = ~n313 & ~n315;
  assign n317 = ~n312 & n316;
  assign n318 = n74 & n86;
  assign n319 = n95 & n318;
  assign n320 = n22 & n74;
  assign n321 = n72 & n320;
  assign n322 = n28 & n114;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~n319 & n323;
  assign n325 = n317 & n324;
  assign n326 = n27 & n40;
  assign n327 = n32 & n326;
  assign n328 = n74 & n249;
  assign n329 = n55 & n249;
  assign n330 = ~n328 & ~n329;
  assign n331 = n27 & n93;
  assign n332 = ~n246 & ~n331;
  assign n333 = n330 & n332;
  assign n334 = n32 & ~n333;
  assign n335 = ~n327 & ~n334;
  assign n336 = n325 & n335;
  assign n337 = n311 & n336;
  assign n338 = n41 & n278;
  assign n339 = n102 & n305;
  assign n340 = n145 & n183;
  assign n341 = n23 & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = ~n338 & n342;
  assign n344 = n79 & n103;
  assign n345 = n343 & ~n344;
  assign n346 = n66 & n169;
  assign n347 = n117 & n199;
  assign n348 = ~n346 & ~n347;
  assign n349 = n95 & n100;
  assign n350 = n31 & n46;
  assign n351 = n66 & n350;
  assign n352 = ~n349 & ~n351;
  assign n353 = n348 & n352;
  assign n354 = n42 & n145;
  assign n355 = n54 & n354;
  assign n356 = n31 & n74;
  assign n357 = n58 & n356;
  assign n358 = ~n355 & ~n357;
  assign n359 = n95 & n180;
  assign n360 = n34 & n46;
  assign n361 = n89 & n360;
  assign n362 = ~n359 & ~n361;
  assign n363 = n358 & n362;
  assign n364 = n37 & n203;
  assign n365 = n40 & n44;
  assign n366 = n102 & n365;
  assign n367 = ~n364 & ~n366;
  assign n368 = n89 & n211;
  assign n369 = n66 & n225;
  assign n370 = ~n368 & ~n369;
  assign n371 = n367 & n370;
  assign n372 = n363 & n371;
  assign n373 = n353 & n372;
  assign n374 = n345 & n373;
  assign n375 = n337 & n374;
  assign n376 = n44 & n183;
  assign n377 = n31 & n44;
  assign n378 = n46 & n183;
  assign n379 = ~n207 & ~n378;
  assign n380 = ~n377 & n379;
  assign n381 = ~n376 & n380;
  assign n382 = n23 & ~n381;
  assign n383 = ~n246 & ~n264;
  assign n384 = ~n211 & n383;
  assign n385 = n95 & ~n384;
  assign n386 = n98 & n145;
  assign n387 = ~n60 & ~n386;
  assign n388 = i_8_ & n168;
  assign n389 = n387 & ~n388;
  assign n390 = ~n109 & n389;
  assign n391 = n117 & ~n390;
  assign n392 = ~n385 & ~n391;
  assign n393 = n67 & n124;
  assign n394 = ~i_5_ & n393;
  assign n395 = n41 & n394;
  assign n396 = n392 & ~n395;
  assign n397 = ~n382 & n396;
  assign n398 = ~n32 & ~n95;
  assign n399 = n55 & n93;
  assign n400 = n44 & n73;
  assign n401 = n32 & n400;
  assign n402 = ~n399 & ~n401;
  assign n403 = ~n398 & ~n402;
  assign n404 = n23 & n356;
  assign n405 = n122 & n213;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n403 & n406;
  assign n408 = ~n305 & ~n328;
  assign n409 = ~n90 & n408;
  assign n410 = n203 & ~n409;
  assign n411 = n40 & n74;
  assign n412 = n99 & n411;
  assign n413 = ~n150 & ~n232;
  assign n414 = n95 & ~n413;
  assign n415 = ~n412 & ~n414;
  assign n416 = ~n410 & n415;
  assign n417 = n407 & n416;
  assign n418 = n44 & n67;
  assign n419 = n66 & n418;
  assign n420 = n125 & n249;
  assign n421 = n79 & n420;
  assign n422 = ~n419 & ~n421;
  assign n423 = n87 & n99;
  assign n424 = n27 & n249;
  assign n425 = n102 & n424;
  assign n426 = ~n423 & ~n425;
  assign n427 = n22 & n36;
  assign n428 = ~n146 & ~n427;
  assign n429 = n102 & ~n428;
  assign n430 = n426 & ~n429;
  assign n431 = ~i_8_ & n194;
  assign n432 = n58 & n431;
  assign n433 = n53 & n68;
  assign n434 = ~n432 & ~n433;
  assign n435 = n430 & n434;
  assign n436 = n422 & n435;
  assign n437 = n417 & n436;
  assign n438 = n74 & n98;
  assign n439 = n25 & n145;
  assign n440 = n48 & n145;
  assign n441 = ~n220 & ~n440;
  assign n442 = ~n439 & n441;
  assign n443 = ~n438 & n442;
  assign n444 = n114 & ~n443;
  assign n445 = n79 & n134;
  assign n446 = ~n203 & ~n445;
  assign n447 = n27 & n113;
  assign n448 = n22 & n55;
  assign n449 = ~n100 & ~n134;
  assign n450 = ~n448 & n449;
  assign n451 = ~n447 & n450;
  assign n452 = ~n446 & ~n451;
  assign n453 = n42 & n74;
  assign n454 = ~n393 & ~n453;
  assign n455 = n66 & ~n454;
  assign n456 = ~i_8_ & n109;
  assign n457 = n122 & n456;
  assign n458 = ~n455 & ~n457;
  assign n459 = ~n452 & n458;
  assign n460 = ~n444 & n459;
  assign n461 = n437 & n460;
  assign n462 = n397 & n461;
  assign n463 = n375 & n462;
  assign o_0_ = ~n289 | ~n463;
  assign n465 = n122 & n220;
  assign n466 = n93 & n125;
  assign n467 = n99 & n466;
  assign n468 = n95 & n265;
  assign n469 = ~n467 & ~n468;
  assign n470 = ~n465 & n469;
  assign n471 = n54 & n418;
  assign n472 = n470 & ~n471;
  assign n473 = n102 & n197;
  assign n474 = n36 & n40;
  assign n475 = ~n235 & ~n474;
  assign n476 = n89 & ~n475;
  assign n477 = ~n473 & ~n476;
  assign n478 = n23 & n218;
  assign n479 = ~i_5_ & n165;
  assign n480 = n99 & n479;
  assign n481 = n40 & n125;
  assign n482 = ~n153 & ~n481;
  assign n483 = n32 & ~n482;
  assign n484 = ~n480 & ~n483;
  assign n485 = ~n478 & n484;
  assign n486 = n477 & n485;
  assign n487 = n472 & n486;
  assign n488 = n49 & n66;
  assign n489 = n79 & n235;
  assign n490 = ~n488 & ~n489;
  assign n491 = n102 & n250;
  assign n492 = n36 & n42;
  assign n493 = n41 & n492;
  assign n494 = ~n491 & ~n493;
  assign n495 = n490 & n494;
  assign n496 = i_8_ & n140;
  assign n497 = n58 & n496;
  assign n498 = n23 & n195;
  assign n499 = ~n497 & ~n498;
  assign n500 = n495 & n499;
  assign n501 = n46 & n249;
  assign n502 = n95 & n501;
  assign n503 = n32 & n75;
  assign n504 = n42 & n46;
  assign n505 = n23 & n504;
  assign n506 = ~n503 & ~n505;
  assign n507 = ~n502 & n506;
  assign n508 = n72 & n264;
  assign n509 = n32 & n365;
  assign n510 = ~n508 & ~n509;
  assign n511 = n36 & n249;
  assign n512 = n79 & n511;
  assign n513 = n117 & n492;
  assign n514 = ~n512 & ~n513;
  assign n515 = n510 & n514;
  assign n516 = n507 & n515;
  assign n517 = n500 & n516;
  assign n518 = n487 & n517;
  assign n519 = n40 & n46;
  assign n520 = ~n427 & ~n519;
  assign n521 = ~n305 & n520;
  assign n522 = ~n400 & n521;
  assign n523 = n89 & ~n522;
  assign n524 = n117 & n141;
  assign n525 = n54 & n184;
  assign n526 = ~n524 & ~n525;
  assign n527 = n65 & n199;
  assign n528 = n56 & n122;
  assign n529 = ~n527 & ~n528;
  assign n530 = n72 & n411;
  assign n531 = n27 & n42;
  assign n532 = n58 & n531;
  assign n533 = ~n530 & ~n532;
  assign n534 = n529 & n533;
  assign n535 = n526 & n534;
  assign n536 = ~n523 & n535;
  assign n537 = n203 & n246;
  assign n538 = n203 & n411;
  assign n539 = n23 & n184;
  assign n540 = ~n538 & ~n539;
  assign n541 = n41 & n438;
  assign n542 = ~n236 & ~n541;
  assign n543 = n540 & n542;
  assign n544 = ~n537 & n543;
  assign n545 = n23 & n260;
  assign n546 = n41 & n242;
  assign n547 = n102 & n328;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n545 & n548;
  assign n550 = n114 & n340;
  assign n551 = n54 & n155;
  assign n552 = ~n550 & ~n551;
  assign n553 = n549 & n552;
  assign n554 = n23 & n438;
  assign n555 = n117 & n314;
  assign n556 = ~n554 & ~n555;
  assign n557 = n58 & n504;
  assign n558 = n203 & n326;
  assign n559 = ~n557 & ~n558;
  assign n560 = n58 & n242;
  assign n561 = n95 & n147;
  assign n562 = ~n560 & ~n561;
  assign n563 = n559 & n562;
  assign n564 = n556 & n563;
  assign n565 = n553 & n564;
  assign n566 = n544 & n565;
  assign n567 = n536 & n566;
  assign n568 = n518 & n567;
  assign n569 = ~n180 & ~n211;
  assign n570 = n102 & ~n569;
  assign n571 = ~n242 & ~n496;
  assign n572 = n54 & ~n571;
  assign n573 = ~n570 & ~n572;
  assign n574 = ~n260 & ~n350;
  assign n575 = n117 & ~n574;
  assign n576 = n573 & ~n575;
  assign n577 = n31 & n36;
  assign n578 = n66 & n577;
  assign n579 = n95 & n424;
  assign n580 = n42 & n125;
  assign n581 = n23 & n580;
  assign n582 = ~n579 & ~n581;
  assign n583 = n79 & n411;
  assign n584 = n114 & n354;
  assign n585 = n122 & n453;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n583 & n586;
  assign n588 = n582 & n587;
  assign n589 = ~n578 & n588;
  assign n590 = n576 & n589;
  assign n591 = n114 & n356;
  assign n592 = n133 & ~n591;
  assign n593 = n102 & n501;
  assign n594 = n54 & n378;
  assign n595 = ~n593 & ~n594;
  assign n596 = n122 & n184;
  assign n597 = n27 & n86;
  assign n598 = n95 & n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = n595 & n599;
  assign n601 = n117 & n577;
  assign n602 = n203 & n399;
  assign n603 = ~n601 & ~n602;
  assign n604 = n27 & n48;
  assign n605 = n41 & n604;
  assign n606 = n72 & n211;
  assign n607 = ~n605 & ~n606;
  assign n608 = n603 & n607;
  assign n609 = n600 & n608;
  assign n610 = n117 & n155;
  assign n611 = n145 & n249;
  assign n612 = n203 & n611;
  assign n613 = n102 & n318;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n610 & n614;
  assign n616 = ~n75 & ~n80;
  assign n617 = n79 & ~n616;
  assign n618 = n615 & ~n617;
  assign n619 = n609 & n618;
  assign n620 = n592 & n619;
  assign n621 = n66 & n260;
  assign n622 = n203 & n481;
  assign n623 = n147 & n203;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~n621 & n624;
  assign n626 = ~n306 & ~n411;
  assign n627 = n32 & ~n626;
  assign n628 = n114 & n243;
  assign n629 = n203 & n427;
  assign n630 = n60 & n114;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n628 & n631;
  assign n633 = ~n627 & n632;
  assign n634 = n54 & n225;
  assign n635 = n114 & n376;
  assign n636 = ~n634 & ~n635;
  assign n637 = n633 & n636;
  assign n638 = n625 & n637;
  assign n639 = n620 & n638;
  assign n640 = n590 & n639;
  assign n641 = n568 & n640;
  assign n642 = n34 & n35;
  assign n643 = n22 & n125;
  assign n644 = ~n642 & ~n643;
  assign n645 = n79 & ~n644;
  assign n646 = ~n80 & ~n165;
  assign n647 = n72 & ~n646;
  assign n648 = ~n196 & ~n647;
  assign n649 = ~n645 & n648;
  assign n650 = ~n49 & ~n580;
  assign n651 = n58 & ~n650;
  assign n652 = ~n421 & ~n651;
  assign n653 = n649 & n652;
  assign n654 = n62 & n653;
  assign n655 = ~n199 & ~n356;
  assign n656 = n54 & ~n655;
  assign n657 = ~n134 & ~n166;
  assign n658 = ~n329 & n657;
  assign n659 = n32 & ~n658;
  assign n660 = ~n153 & ~n306;
  assign n661 = ~n235 & n660;
  assign n662 = n102 & ~n661;
  assign n663 = n99 & n103;
  assign n664 = n59 & n74;
  assign n665 = ~n492 & ~n664;
  assign n666 = n66 & ~n665;
  assign n667 = ~n663 & ~n666;
  assign n668 = ~n662 & n667;
  assign n669 = ~n659 & n668;
  assign n670 = ~n656 & n669;
  assign n671 = n37 & n99;
  assign n672 = n46 & n98;
  assign n673 = n117 & n672;
  assign n674 = ~n671 & ~n673;
  assign n675 = n58 & n453;
  assign n676 = n41 & n577;
  assign n677 = ~n675 & ~n676;
  assign n678 = n674 & n677;
  assign n679 = n46 & n93;
  assign n680 = ~n519 & ~n679;
  assign n681 = ~n329 & n680;
  assign n682 = ~n265 & n681;
  assign n683 = n203 & ~n682;
  assign n684 = ~n223 & ~n230;
  assign n685 = ~n604 & n684;
  assign n686 = n23 & ~n685;
  assign n687 = ~n683 & ~n686;
  assign n688 = n678 & n687;
  assign n689 = n670 & n688;
  assign n690 = n95 & n306;
  assign n691 = n99 & n420;
  assign n692 = ~n219 & ~n691;
  assign n693 = ~n690 & n692;
  assign n694 = ~n208 & ~n418;
  assign n695 = n41 & ~n694;
  assign n696 = n693 & ~n695;
  assign n697 = n114 & n456;
  assign n698 = ~n195 & ~n218;
  assign n699 = n114 & ~n698;
  assign n700 = ~n697 & ~n699;
  assign n701 = n696 & n700;
  assign n702 = n174 & n701;
  assign n703 = n689 & n702;
  assign n704 = n654 & n703;
  assign o_1_ = ~n641 | ~n704;
  assign n706 = n31 & n125;
  assign n707 = ~n580 & ~n706;
  assign n708 = n117 & ~n707;
  assign n709 = n122 & n394;
  assign n710 = ~n326 & ~n474;
  assign n711 = n79 & ~n710;
  assign n712 = ~n709 & ~n711;
  assign n713 = ~n708 & n712;
  assign n714 = n633 & n713;
  assign n715 = ~n139 & ~n456;
  assign n716 = n58 & ~n715;
  assign n717 = ~n90 & ~n235;
  assign n718 = ~n481 & n717;
  assign n719 = n99 & ~n718;
  assign n720 = ~n716 & ~n719;
  assign n721 = n41 & n169;
  assign n722 = ~n376 & ~n604;
  assign n723 = ~n208 & n722;
  assign n724 = n54 & ~n723;
  assign n725 = ~n134 & ~n611;
  assign n726 = n102 & ~n725;
  assign n727 = n117 & n340;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n724 & n728;
  assign n730 = ~n721 & n729;
  assign n731 = n720 & n730;
  assign n732 = n714 & n731;
  assign n733 = n58 & n388;
  assign n734 = ~n359 & ~n733;
  assign n735 = n25 & n125;
  assign n736 = n122 & n735;
  assign n737 = n559 & ~n736;
  assign n738 = n734 & n737;
  assign n739 = ~n329 & ~n611;
  assign n740 = n89 & ~n739;
  assign n741 = n23 & n394;
  assign n742 = ~n445 & ~n538;
  assign n743 = ~n741 & n742;
  assign n744 = ~n740 & n743;
  assign n745 = n738 & n744;
  assign n746 = n66 & n531;
  assign n747 = ~n466 & ~n511;
  assign n748 = n95 & ~n747;
  assign n749 = ~n746 & ~n748;
  assign n750 = n23 & n208;
  assign n751 = n203 & n597;
  assign n752 = ~n750 & ~n751;
  assign n753 = n72 & n175;
  assign n754 = n54 & n220;
  assign n755 = ~n753 & ~n754;
  assign n756 = n752 & n755;
  assign n757 = n749 & n756;
  assign n758 = n45 & n66;
  assign n759 = n99 & n643;
  assign n760 = n32 & n427;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~n758 & n761;
  assign n763 = n66 & n195;
  assign n764 = ~n593 & ~n763;
  assign n765 = n762 & n764;
  assign n766 = n757 & n765;
  assign n767 = n745 & n766;
  assign n768 = n437 & n767;
  assign n769 = n58 & n418;
  assign n770 = n36 & n48;
  assign n771 = n41 & n770;
  assign n772 = ~n769 & ~n771;
  assign n773 = n352 & n772;
  assign n774 = n75 & n102;
  assign n775 = n122 & n531;
  assign n776 = ~n774 & ~n775;
  assign n777 = n32 & n147;
  assign n778 = n79 & n150;
  assign n779 = ~n777 & ~n778;
  assign n780 = n89 & n328;
  assign n781 = n102 & n597;
  assign n782 = ~n780 & ~n781;
  assign n783 = n779 & n782;
  assign n784 = n776 & n783;
  assign n785 = ~n56 & ~n207;
  assign n786 = n66 & ~n785;
  assign n787 = n93 & n126;
  assign n788 = n89 & n175;
  assign n789 = n79 & n331;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n787 & n790;
  assign n792 = ~n786 & n791;
  assign n793 = n784 & n792;
  assign n794 = n773 & n793;
  assign n795 = n44 & n98;
  assign n796 = ~n664 & ~n795;
  assign n797 = n114 & ~n796;
  assign n798 = n72 & n93;
  assign n799 = n35 & n798;
  assign n800 = ~n797 & ~n799;
  assign n801 = n99 & n246;
  assign n802 = n66 & n155;
  assign n803 = n102 & n511;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n801 & n804;
  assign n806 = n36 & n86;
  assign n807 = ~n87 & ~n806;
  assign n808 = ~n250 & n807;
  assign n809 = n203 & ~n808;
  assign n810 = n89 & n299;
  assign n811 = n32 & n466;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n809 & n812;
  assign n814 = n805 & n813;
  assign n815 = n800 & n814;
  assign n816 = n794 & n815;
  assign n817 = n768 & n816;
  assign n818 = n732 & n817;
  assign n819 = n66 & n388;
  assign n820 = n102 & n299;
  assign n821 = ~n819 & ~n820;
  assign n822 = n99 & n150;
  assign n823 = n23 & n440;
  assign n824 = n95 & n177;
  assign n825 = ~n823 & ~n824;
  assign n826 = n102 & n162;
  assign n827 = n825 & ~n826;
  assign n828 = ~n822 & n827;
  assign n829 = n58 & n672;
  assign n830 = n102 & n150;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n368 & n831;
  assign n833 = n828 & n832;
  assign n834 = n821 & n833;
  assign n835 = n66 & n213;
  assign n836 = n79 & n162;
  assign n837 = ~n835 & ~n836;
  assign n838 = n54 & n440;
  assign n839 = n837 & ~n838;
  assign n840 = n58 & n386;
  assign n841 = n99 & n306;
  assign n842 = n72 & n318;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n840 & n843;
  assign n845 = n839 & n844;
  assign n846 = ~n162 & ~n511;
  assign n847 = n203 & ~n846;
  assign n848 = n32 & n424;
  assign n849 = n95 & n448;
  assign n850 = ~n848 & ~n849;
  assign n851 = n23 & n388;
  assign n852 = n850 & ~n851;
  assign n853 = ~n847 & n852;
  assign n854 = n845 & n853;
  assign n855 = ~n184 & ~n354;
  assign n856 = n66 & ~n855;
  assign n857 = n28 & n58;
  assign n858 = n95 & n299;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n361 & n859;
  assign n861 = ~n856 & n860;
  assign n862 = n73 & n124;
  assign n863 = ~i_5_ & n862;
  assign n864 = ~n130 & ~n643;
  assign n865 = ~n863 & n864;
  assign n866 = ~n37 & n865;
  assign n867 = n95 & ~n866;
  assign n868 = n861 & ~n867;
  assign n869 = n854 & n868;
  assign n870 = n117 & n354;
  assign n871 = ~n613 & ~n870;
  assign n872 = ~n447 & ~n643;
  assign n873 = n102 & ~n872;
  assign n874 = n58 & n350;
  assign n875 = n41 & n580;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n873 & n876;
  assign n878 = n871 & n877;
  assign n879 = n517 & n878;
  assign n880 = n869 & n879;
  assign n881 = n834 & n880;
  assign o_2_ = ~n818 | ~n881;
  assign n883 = ~n119 & n387;
  assign n884 = n23 & ~n883;
  assign n885 = n286 & ~n884;
  assign n886 = n590 & n885;
  assign n887 = n119 & n122;
  assign n888 = n80 & n203;
  assign n889 = ~n887 & ~n888;
  assign n890 = n99 & n146;
  assign n891 = n889 & ~n890;
  assign n892 = ~n69 & ~n664;
  assign n893 = n41 & ~n892;
  assign n894 = n89 & n424;
  assign n895 = ~n357 & ~n894;
  assign n896 = ~n893 & n895;
  assign n897 = n891 & n896;
  assign n898 = ~n177 & ~n447;
  assign n899 = ~n103 & n898;
  assign n900 = ~n87 & n899;
  assign n901 = n32 & ~n900;
  assign n902 = n80 & n102;
  assign n903 = n117 & n278;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n901 & n904;
  assign n906 = ~n735 & ~n795;
  assign n907 = ~n243 & n906;
  assign n908 = ~n223 & n907;
  assign n909 = n41 & ~n908;
  assign n910 = n99 & n204;
  assign n911 = ~n909 & ~n910;
  assign n912 = n905 & n911;
  assign n913 = n897 & n912;
  assign n914 = n886 & n913;
  assign n915 = ~n453 & ~n496;
  assign n916 = n117 & ~n915;
  assign n917 = n58 & n604;
  assign n918 = ~n916 & ~n917;
  assign n919 = n58 & n440;
  assign n920 = ~n466 & ~n863;
  assign n921 = n79 & ~n920;
  assign n922 = ~n919 & ~n921;
  assign n923 = n918 & n922;
  assign n924 = n23 & n45;
  assign n925 = n122 & n207;
  assign n926 = n99 & n318;
  assign n927 = ~n925 & ~n926;
  assign n928 = ~n924 & n927;
  assign n929 = n36 & n93;
  assign n930 = ~n320 & ~n929;
  assign n931 = n89 & ~n930;
  assign n932 = n72 & n246;
  assign n933 = ~n622 & ~n932;
  assign n934 = ~n697 & n933;
  assign n935 = ~n931 & n934;
  assign n936 = n928 & n935;
  assign n937 = n923 & n936;
  assign n938 = n767 & n937;
  assign n939 = n122 & n496;
  assign n940 = n54 & n110;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n400 & ~n806;
  assign n943 = n102 & ~n942;
  assign n944 = ~n602 & ~n943;
  assign n945 = ~n291 & ~n360;
  assign n946 = ~n163 & ~n945;
  assign n947 = ~n130 & ~n150;
  assign n948 = n89 & ~n947;
  assign n949 = ~n293 & ~n377;
  assign n950 = n66 & ~n949;
  assign n951 = ~n948 & ~n950;
  assign n952 = ~n946 & n951;
  assign n953 = n944 & n952;
  assign n954 = n941 & n953;
  assign n955 = n938 & n954;
  assign n956 = n914 & n955;
  assign n957 = n23 & n492;
  assign n958 = ~n180 & ~n246;
  assign n959 = ~n511 & n958;
  assign n960 = ~n597 & n959;
  assign n961 = n32 & ~n960;
  assign n962 = ~n957 & ~n961;
  assign n963 = ~n260 & n441;
  assign n964 = n41 & ~n963;
  assign n965 = n117 & n456;
  assign n966 = n60 & n66;
  assign n967 = ~n530 & ~n966;
  assign n968 = ~n965 & n967;
  assign n969 = ~n153 & ~n328;
  assign n970 = ~n611 & n969;
  assign n971 = n95 & ~n970;
  assign n972 = n968 & ~n971;
  assign n973 = ~n964 & n972;
  assign n974 = ~n169 & ~n230;
  assign n975 = n54 & ~n974;
  assign n976 = n203 & n466;
  assign n977 = n130 & n203;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n478 & n978;
  assign n980 = ~n975 & n979;
  assign n981 = n72 & n265;
  assign n982 = n122 & n664;
  assign n983 = ~n981 & ~n982;
  assign n984 = n79 & n400;
  assign n985 = n983 & ~n984;
  assign n986 = n980 & n985;
  assign n987 = n973 & n986;
  assign n988 = n962 & n987;
  assign n989 = ~n134 & ~n211;
  assign n990 = n95 & ~n989;
  assign n991 = ~n264 & ~n328;
  assign n992 = n32 & ~n991;
  assign n993 = ~n990 & ~n992;
  assign n994 = ~n293 & ~n453;
  assign n995 = n58 & ~n994;
  assign n996 = n993 & ~n995;
  assign n997 = ~n171 & ~n350;
  assign n998 = n114 & ~n997;
  assign n999 = n41 & n199;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = n996 & n1000;
  assign n1002 = n54 & n377;
  assign n1003 = ~n355 & ~n1002;
  assign n1004 = ~n87 & ~n204;
  assign n1005 = n102 & ~n1004;
  assign n1006 = ~n88 & ~n1005;
  assign n1007 = n72 & n103;
  assign n1008 = n66 & n439;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = n1006 & n1009;
  assign n1011 = n1003 & n1010;
  assign n1012 = n1001 & n1011;
  assign n1013 = ~n501 & ~n863;
  assign n1014 = n99 & ~n1013;
  assign n1015 = n1012 & ~n1014;
  assign n1016 = n72 & n400;
  assign n1017 = n114 & n377;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = n41 & n531;
  assign n1020 = n79 & n187;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = n203 & n365;
  assign n1023 = n1021 & ~n1022;
  assign n1024 = n1018 & n1023;
  assign n1025 = n95 & n479;
  assign n1026 = n54 & n531;
  assign n1027 = ~n610 & ~n1026;
  assign n1028 = ~n1025 & n1027;
  assign n1029 = ~n37 & n660;
  assign n1030 = n203 & ~n1029;
  assign n1031 = n1028 & ~n1030;
  assign n1032 = n1024 & n1031;
  assign n1033 = ~n340 & ~n735;
  assign n1034 = ~n255 & n1033;
  assign n1035 = n58 & ~n1034;
  assign n1036 = ~n171 & ~n388;
  assign n1037 = n122 & ~n1036;
  assign n1038 = ~n1035 & ~n1037;
  assign n1039 = n95 & n420;
  assign n1040 = n41 & n60;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = n348 & n1041;
  assign n1043 = n148 & ~n150;
  assign n1044 = n72 & ~n1043;
  assign n1045 = n79 & n211;
  assign n1046 = n69 & n117;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n1044 & n1047;
  assign n1049 = n1042 & n1048;
  assign n1050 = n1038 & n1049;
  assign n1051 = n1032 & n1050;
  assign n1052 = n1015 & n1051;
  assign n1053 = n988 & n1052;
  assign o_3_ = ~n956 | ~n1053;
  assign n1055 = ~n225 & ~n293;
  assign n1056 = n117 & ~n1055;
  assign n1057 = n54 & n260;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~n447 & ~n806;
  assign n1060 = ~n235 & n1059;
  assign n1061 = n32 & ~n1060;
  assign n1062 = n66 & n141;
  assign n1063 = n102 & n466;
  assign n1064 = n23 & n418;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = ~n1062 & n1065;
  assign n1067 = ~n1061 & n1066;
  assign n1068 = n1058 & n1067;
  assign n1069 = n175 & n203;
  assign n1070 = n58 & n376;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = n32 & n501;
  assign n1073 = n95 & n153;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n741 & n1074;
  assign n1076 = n1071 & n1075;
  assign n1077 = n1068 & n1076;
  assign n1078 = ~n223 & ~n672;
  assign n1079 = n66 & ~n1078;
  assign n1080 = ~n114 & ~n122;
  assign n1081 = n604 & ~n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign n1083 = n203 & n420;
  assign n1084 = n122 & n770;
  assign n1085 = ~n1083 & ~n1084;
  assign n1086 = ~n200 & ~n366;
  assign n1087 = n1085 & n1086;
  assign n1088 = n1082 & n1087;
  assign n1089 = n41 & n706;
  assign n1090 = n58 & n795;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = n203 & n424;
  assign n1093 = n32 & n679;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = n99 & n597;
  assign n1096 = n95 & n326;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = n1094 & n1097;
  assign n1099 = n1091 & n1098;
  assign n1100 = n1088 & n1099;
  assign n1101 = n1077 & n1100;
  assign n1102 = n854 & n1101;
  assign n1103 = ~n119 & ~n225;
  assign n1104 = n114 & ~n1103;
  assign n1105 = ~n305 & ~n329;
  assign n1106 = n99 & ~n1105;
  assign n1107 = ~n1104 & ~n1106;
  assign n1108 = n117 & n213;
  assign n1109 = n102 & n265;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = n95 & n447;
  assign n1112 = n79 & n447;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n1110 & n1113;
  assign n1115 = n1107 & n1114;
  assign n1116 = ~n439 & ~n770;
  assign n1117 = ~n139 & n1116;
  assign n1118 = n23 & ~n1117;
  assign n1119 = ~n87 & ~n175;
  assign n1120 = n102 & ~n1119;
  assign n1121 = ~n939 & ~n1120;
  assign n1122 = ~n1118 & n1121;
  assign n1123 = n1115 & n1122;
  assign n1124 = n1102 & n1123;
  assign n1125 = n271 & n639;
  assign n1126 = n95 & n305;
  assign n1127 = n79 & n177;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n41 & n356;
  assign n1130 = n66 & n735;
  assign n1131 = n114 & n706;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1129 & n1132;
  assign n1134 = n1128 & n1133;
  assign n1135 = ~n340 & ~n456;
  assign n1136 = ~n230 & n1135;
  assign n1137 = n54 & ~n1136;
  assign n1138 = n203 & n479;
  assign n1139 = n58 & n438;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = i_5_ & n862;
  assign n1142 = n102 & n1141;
  assign n1143 = ~n763 & ~n1142;
  assign n1144 = n1140 & n1143;
  assign n1145 = ~n1137 & n1144;
  assign n1146 = n1134 & n1145;
  assign n1147 = ~n377 & ~n453;
  assign n1148 = n41 & ~n1147;
  assign n1149 = ~n28 & ~n293;
  assign n1150 = n54 & ~n1149;
  assign n1151 = n72 & ~n864;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n426 & n1152;
  assign n1154 = ~n1148 & n1153;
  assign n1155 = ~n187 & ~n204;
  assign n1156 = n89 & ~n1155;
  assign n1157 = ~n976 & ~n1156;
  assign n1158 = n297 & n1157;
  assign n1159 = n1154 & n1158;
  assign n1160 = n1146 & n1159;
  assign n1161 = ~n220 & n722;
  assign n1162 = n117 & ~n1161;
  assign n1163 = ~n166 & ~n318;
  assign n1164 = n203 & ~n1163;
  assign n1165 = n749 & ~n1164;
  assign n1166 = ~n1162 & n1165;
  assign n1167 = n36 & n64;
  assign n1168 = ~n305 & ~n474;
  assign n1169 = ~n1167 & n1168;
  assign n1170 = n32 & ~n1169;
  assign n1171 = ~n706 & ~n795;
  assign n1172 = ~n293 & n1171;
  assign n1173 = n122 & ~n1172;
  assign n1174 = ~n1170 & ~n1173;
  assign n1175 = ~n184 & ~n278;
  assign n1176 = n58 & ~n1175;
  assign n1177 = ~n163 & n1141;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = n66 & n278;
  assign n1180 = ~n224 & ~n1179;
  assign n1181 = ~n225 & ~n377;
  assign n1182 = n122 & ~n1181;
  assign n1183 = n1180 & ~n1182;
  assign n1184 = n1178 & n1183;
  assign n1185 = ~n121 & ~n340;
  assign n1186 = ~n28 & n1185;
  assign n1187 = n66 & ~n1186;
  assign n1188 = ~n78 & ~n98;
  assign n1189 = n806 & ~n1188;
  assign n1190 = ~n1187 & ~n1189;
  assign n1191 = n1184 & n1190;
  assign n1192 = n1174 & n1191;
  assign n1193 = n1166 & n1192;
  assign n1194 = n1160 & n1193;
  assign n1195 = n1125 & n1194;
  assign o_4_ = ~n1124 | ~n1195;
  assign n1197 = ~n195 & ~n243;
  assign n1198 = ~n45 & n1197;
  assign n1199 = ~n110 & n1198;
  assign n1200 = n58 & ~n1199;
  assign n1201 = ~n492 & ~n580;
  assign n1202 = ~n496 & n1201;
  assign n1203 = ~n672 & n1202;
  assign n1204 = n114 & ~n1203;
  assign n1205 = ~n1200 & ~n1204;
  assign n1206 = n53 & n394;
  assign n1207 = n95 & n365;
  assign n1208 = n102 & n264;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n412 & n1209;
  assign n1211 = ~n1206 & n1210;
  assign n1212 = ~n448 & ~n929;
  assign n1213 = ~n424 & n710;
  assign n1214 = n1212 & n1213;
  assign n1215 = ~n147 & n1214;
  assign n1216 = n99 & ~n1215;
  assign n1217 = n1211 & ~n1216;
  assign n1218 = n1205 & n1217;
  assign n1219 = n861 & n1076;
  assign n1220 = n86 & n171;
  assign n1221 = n190 & ~n1220;
  assign n1222 = n1219 & n1221;
  assign n1223 = ~n306 & n330;
  assign n1224 = n79 & ~n1223;
  assign n1225 = ~n208 & ~n293;
  assign n1226 = n117 & ~n1225;
  assign n1227 = ~n1224 & ~n1226;
  assign n1228 = n1222 & n1227;
  assign n1229 = n1218 & n1228;
  assign n1230 = n348 & ~n820;
  assign n1231 = n41 & n418;
  assign n1232 = ~n327 & ~n1231;
  assign n1233 = ~n104 & ~n903;
  assign n1234 = n1232 & n1233;
  assign n1235 = ~n221 & ~n532;
  assign n1236 = n1234 & n1235;
  assign n1237 = n1230 & n1236;
  assign n1238 = ~n593 & ~n746;
  assign n1239 = ~n1179 & n1238;
  assign n1240 = n95 & n611;
  assign n1241 = ~n1127 & ~n1240;
  assign n1242 = n263 & n1241;
  assign n1243 = n1239 & n1242;
  assign n1244 = n1237 & n1243;
  assign n1245 = n110 & n114;
  assign n1246 = n89 & n481;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = n32 & n1141;
  assign n1249 = n89 & n447;
  assign n1250 = n49 & n54;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1248 & n1251;
  assign n1253 = n66 & n112;
  assign n1254 = n122 & n139;
  assign n1255 = n72 & n197;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n1253 & n1256;
  assign n1258 = n114 & n141;
  assign n1259 = n58 & n354;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n180 & n203;
  assign n1262 = n89 & n399;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n1260 & n1263;
  assign n1265 = n1257 & n1264;
  assign n1266 = n1252 & n1265;
  assign n1267 = n1247 & n1266;
  assign n1268 = n1244 & n1267;
  assign n1269 = ~n80 & ~n320;
  assign n1270 = ~n420 & n1269;
  assign n1271 = n32 & ~n1270;
  assign n1272 = n487 & ~n1271;
  assign n1273 = n1268 & n1272;
  assign n1274 = n1229 & n1273;
  assign n1275 = n23 & n453;
  assign n1276 = n1012 & ~n1275;
  assign n1277 = n122 & n155;
  assign n1278 = n66 & n378;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n100 & ~n365;
  assign n1281 = n72 & ~n1280;
  assign n1282 = ~n493 & ~n613;
  assign n1283 = n752 & n1282;
  assign n1284 = ~n1281 & n1283;
  assign n1285 = n1279 & n1284;
  assign n1286 = ~n146 & ~n197;
  assign n1287 = n203 & ~n1286;
  assign n1288 = n102 & n863;
  assign n1289 = ~n254 & ~n401;
  assign n1290 = ~n1288 & n1289;
  assign n1291 = ~n1287 & n1290;
  assign n1292 = i_8_ & i_9_;
  assign n1293 = ~n24 & n1292;
  assign n1294 = n94 & n1293;
  assign n1295 = n317 & ~n1294;
  assign n1296 = n1291 & n1295;
  assign n1297 = n1285 & n1296;
  assign n1298 = ~n770 & ~n795;
  assign n1299 = ~n350 & n1298;
  assign n1300 = ~n386 & n1299;
  assign n1301 = n54 & ~n1300;
  assign n1302 = n43 & n183;
  assign n1303 = ~n431 & ~n1302;
  assign n1304 = n122 & ~n1303;
  assign n1305 = n95 & n250;
  assign n1306 = ~n1131 & ~n1305;
  assign n1307 = ~n1304 & n1306;
  assign n1308 = ~n1301 & n1307;
  assign n1309 = n1297 & n1308;
  assign n1310 = n1276 & n1309;
  assign n1311 = ~n420 & ~n863;
  assign n1312 = n89 & ~n1311;
  assign n1313 = ~n208 & ~n456;
  assign n1314 = n66 & ~n1313;
  assign n1315 = ~n1312 & ~n1314;
  assign n1316 = n87 & n89;
  assign n1317 = n95 & n166;
  assign n1318 = n117 & n440;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~n1316 & n1319;
  assign n1321 = n99 & n328;
  assign n1322 = n79 & n1141;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~n498 & ~n628;
  assign n1325 = n1323 & n1324;
  assign n1326 = n1320 & n1325;
  assign n1327 = n54 & n439;
  assign n1328 = n95 & n175;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = n99 & n166;
  assign n1331 = n1329 & ~n1330;
  assign n1332 = ~n112 & ~n386;
  assign n1333 = n41 & ~n1332;
  assign n1334 = n28 & n122;
  assign n1335 = n636 & ~n1334;
  assign n1336 = ~n1333 & n1335;
  assign n1337 = n1331 & n1336;
  assign n1338 = n1326 & n1337;
  assign n1339 = n1315 & n1338;
  assign n1340 = n1310 & n1339;
  assign o_5_ = ~n1274 | ~n1340;
  assign n1342 = ~n230 & ~n376;
  assign n1343 = ~n580 & n1342;
  assign n1344 = n66 & ~n1343;
  assign n1345 = ~n147 & ~n479;
  assign n1346 = n102 & ~n1345;
  assign n1347 = ~n56 & ~n504;
  assign n1348 = ~n229 & n1347;
  assign n1349 = n41 & ~n1348;
  assign n1350 = ~n1346 & ~n1349;
  assign n1351 = ~n1344 & n1350;
  assign n1352 = ~n199 & ~n260;
  assign n1353 = n58 & ~n1352;
  assign n1354 = ~n643 & ~n863;
  assign n1355 = n32 & ~n1354;
  assign n1356 = ~n1353 & ~n1355;
  assign n1357 = n23 & n456;
  assign n1358 = n89 & n448;
  assign n1359 = n72 & n326;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1357 & n1360;
  assign n1362 = n678 & n1361;
  assign n1363 = n1356 & n1362;
  assign n1364 = n1351 & n1363;
  assign n1365 = ~n194 & ~n439;
  assign n1366 = n117 & ~n1365;
  assign n1367 = n1257 & ~n1366;
  assign n1368 = n470 & n1367;
  assign n1369 = n1326 & n1368;
  assign n1370 = n1364 & n1369;
  assign n1371 = n375 & n1370;
  assign n1372 = i_6_ & n1141;
  assign n1373 = ~n100 & ~n1372;
  assign n1374 = ~n77 & n1292;
  assign n1375 = ~n1373 & n1374;
  assign n1376 = n30 & n36;
  assign n1377 = ~n706 & ~n1376;
  assign n1378 = n54 & ~n1377;
  assign n1379 = ~n601 & ~n781;
  assign n1380 = ~n1378 & n1379;
  assign n1381 = ~n1375 & n1380;
  assign n1382 = ~n162 & ~n177;
  assign n1383 = n72 & ~n1382;
  assign n1384 = ~n513 & ~n558;
  assign n1385 = ~n1383 & n1384;
  assign n1386 = n805 & n1385;
  assign n1387 = n1381 & n1386;
  assign n1388 = ~n386 & ~n418;
  assign n1389 = ~n171 & n1388;
  assign n1390 = ~n184 & n1389;
  assign n1391 = n114 & ~n1390;
  assign n1392 = n37 & n89;
  assign n1393 = ~n982 & ~n1392;
  assign n1394 = ~n1391 & n1393;
  assign n1395 = n95 & ~n717;
  assign n1396 = ~n163 & n304;
  assign n1397 = n831 & ~n1396;
  assign n1398 = ~n1395 & n1397;
  assign n1399 = ~n197 & ~n320;
  assign n1400 = n99 & ~n1399;
  assign n1401 = ~n331 & ~n400;
  assign n1402 = n203 & ~n1401;
  assign n1403 = ~n1400 & ~n1402;
  assign n1404 = n1398 & n1403;
  assign n1405 = n1394 & n1404;
  assign n1406 = n1387 & n1405;
  assign n1407 = ~n598 & ~n1111;
  assign n1408 = ~n1277 & n1407;
  assign n1409 = n203 & n360;
  assign n1410 = n102 & n320;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~n691 & n1411;
  assign n1413 = n1408 & n1412;
  assign n1414 = n49 & n114;
  assign n1415 = n72 & n399;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = n89 & n511;
  assign n1418 = n1416 & ~n1417;
  assign n1419 = n58 & n664;
  assign n1420 = n79 & n679;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1418 & n1421;
  assign n1423 = n1413 & n1422;
  assign n1424 = ~n68 & ~n604;
  assign n1425 = ~n139 & n1424;
  assign n1426 = ~n110 & n1425;
  assign n1427 = n23 & ~n1426;
  assign n1428 = ~n126 & ~n218;
  assign n1429 = n66 & ~n1428;
  assign n1430 = ~n778 & ~n1429;
  assign n1431 = ~n1427 & n1430;
  assign n1432 = n1423 & n1431;
  assign n1433 = n937 & n1432;
  assign n1434 = n79 & n365;
  assign n1435 = n58 & n218;
  assign n1436 = n122 & n580;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = n89 & n180;
  assign n1439 = n1437 & ~n1438;
  assign n1440 = ~n1434 & n1439;
  assign n1441 = n122 & n378;
  assign n1442 = n23 & n354;
  assign n1443 = ~n1441 & ~n1442;
  assign n1444 = n75 & n95;
  assign n1445 = n79 & n265;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = n1443 & n1446;
  assign n1448 = n1440 & n1447;
  assign n1449 = n1146 & n1448;
  assign n1450 = n1433 & n1449;
  assign n1451 = n1406 & n1450;
  assign o_6_ = ~n1371 | ~n1451;
  assign n1453 = n32 & n360;
  assign n1454 = ~n250 & ~n448;
  assign n1455 = n102 & ~n1454;
  assign n1456 = ~n1453 & ~n1455;
  assign n1457 = ~n156 & ~n981;
  assign n1458 = n1456 & n1457;
  assign n1459 = n68 & n122;
  assign n1460 = ~n432 & ~n1459;
  assign n1461 = n23 & n126;
  assign n1462 = n95 & n329;
  assign n1463 = n89 & n466;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = ~n1461 & n1464;
  assign n1466 = n1460 & n1465;
  assign n1467 = n1458 & n1466;
  assign n1468 = ~n1093 & ~n1444;
  assign n1469 = ~n788 & n1468;
  assign n1470 = n1028 & n1469;
  assign n1471 = n1467 & n1470;
  assign n1472 = ~n162 & ~n204;
  assign n1473 = n32 & ~n1472;
  assign n1474 = n79 & n180;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n23 & n243;
  assign n1477 = n1475 & ~n1476;
  assign n1478 = n1440 & n1477;
  assign n1479 = ~n278 & ~n453;
  assign n1480 = n114 & ~n1479;
  assign n1481 = n41 & n496;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n447 & ~n511;
  assign n1484 = n99 & ~n1483;
  assign n1485 = n89 & n318;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n1247 & n1486;
  assign n1488 = n1482 & n1487;
  assign n1489 = n1478 & n1488;
  assign n1490 = ~n69 & ~n350;
  assign n1491 = ~n242 & n1490;
  assign n1492 = n122 & ~n1491;
  assign n1493 = ~n359 & ~n583;
  assign n1494 = ~n198 & ~n917;
  assign n1495 = n1493 & n1494;
  assign n1496 = n624 & n1495;
  assign n1497 = ~n480 & n1496;
  assign n1498 = ~n1492 & n1497;
  assign n1499 = n1489 & n1498;
  assign n1500 = n1471 & n1499;
  assign n1501 = ~n377 & ~n492;
  assign n1502 = ~n208 & n1501;
  assign n1503 = n58 & ~n1502;
  assign n1504 = ~n331 & ~n929;
  assign n1505 = ~n90 & n1504;
  assign n1506 = ~n232 & n1505;
  assign n1507 = n102 & ~n1506;
  assign n1508 = ~n1503 & ~n1507;
  assign n1509 = n58 & n770;
  assign n1510 = n102 & n326;
  assign n1511 = n32 & n146;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = ~n1509 & n1512;
  assign n1514 = n122 & n169;
  assign n1515 = n490 & ~n1514;
  assign n1516 = n1513 & n1515;
  assign n1517 = n117 & n208;
  assign n1518 = n68 & n114;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = n23 & n56;
  assign n1521 = n203 & n211;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = n1519 & n1522;
  assign n1524 = n1110 & n1523;
  assign n1525 = n1516 & n1524;
  assign n1526 = ~n597 & n1059;
  assign n1527 = n72 & ~n1526;
  assign n1528 = ~n264 & ~n863;
  assign n1529 = n203 & ~n1528;
  assign n1530 = ~n1527 & ~n1529;
  assign n1531 = n1525 & n1530;
  assign n1532 = n1508 & n1531;
  assign n1533 = n1068 & n1337;
  assign n1534 = n85 & n1533;
  assign n1535 = n1532 & n1534;
  assign n1536 = ~n243 & n379;
  assign n1537 = ~n169 & n1536;
  assign n1538 = n117 & ~n1537;
  assign n1539 = n564 & ~n1538;
  assign n1540 = n1024 & n1539;
  assign n1541 = ~n187 & ~n320;
  assign n1542 = ~n328 & n1541;
  assign n1543 = n95 & ~n1542;
  assign n1544 = ~n314 & ~n795;
  assign n1545 = ~n155 & n1544;
  assign n1546 = n23 & ~n1545;
  assign n1547 = ~n1543 & ~n1546;
  assign n1548 = ~n68 & ~n453;
  assign n1549 = ~n213 & n1548;
  assign n1550 = n54 & ~n1549;
  assign n1551 = ~n110 & ~n119;
  assign n1552 = ~n314 & n1551;
  assign n1553 = n66 & ~n1552;
  assign n1554 = ~n1550 & ~n1553;
  assign n1555 = n1547 & n1554;
  assign n1556 = n1540 & n1555;
  assign n1557 = n834 & n1556;
  assign n1558 = n1535 & n1557;
  assign o_7_ = ~n1500 | ~n1558;
  assign n1560 = n616 & n1286;
  assign n1561 = ~n232 & n1560;
  assign n1562 = n89 & ~n1561;
  assign n1563 = n241 & ~n1562;
  assign n1564 = ~n169 & ~n735;
  assign n1565 = ~n121 & n1564;
  assign n1566 = n114 & ~n1565;
  assign n1567 = n1211 & ~n1566;
  assign n1568 = n1563 & n1567;
  assign n1569 = n725 & ~n862;
  assign n1570 = n72 & ~n1569;
  assign n1571 = ~n386 & ~n577;
  assign n1572 = ~n314 & n1571;
  assign n1573 = n122 & ~n1572;
  assign n1574 = ~n1570 & ~n1573;
  assign n1575 = n1525 & n1574;
  assign n1576 = n1432 & n1575;
  assign n1577 = n89 & n501;
  assign n1578 = n79 & n100;
  assign n1579 = n66 & n438;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1577 & n1580;
  assign n1582 = ~n306 & ~n481;
  assign n1583 = n72 & ~n1582;
  assign n1584 = ~n811 & ~n1583;
  assign n1585 = n1581 & n1584;
  assign n1586 = ~n119 & ~n440;
  assign n1587 = ~n735 & n1586;
  assign n1588 = n54 & ~n1587;
  assign n1589 = n95 & n1141;
  assign n1590 = n114 & n139;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = ~n1588 & n1591;
  assign n1593 = n1585 & n1592;
  assign n1594 = n1576 & n1593;
  assign n1595 = n1568 & n1594;
  assign n1596 = ~n28 & ~n171;
  assign n1597 = n41 & ~n1596;
  assign n1598 = n32 & ~n1454;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = n43 & n59;
  assign n1601 = ~n492 & ~n1600;
  assign n1602 = n54 & ~n1601;
  assign n1603 = ~n75 & ~n611;
  assign n1604 = n203 & ~n1603;
  assign n1605 = ~n1602 & ~n1604;
  assign n1606 = n1599 & n1605;
  assign n1607 = n553 & n1606;
  assign n1608 = n95 & n331;
  assign n1609 = n117 & n377;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = n510 & n1610;
  assign n1612 = n343 & n1611;
  assign n1613 = ~n49 & n906;
  assign n1614 = n117 & ~n1613;
  assign n1615 = n65 & n356;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = n1612 & n1616;
  assign n1618 = n1607 & n1617;
  assign n1619 = ~n519 & ~n611;
  assign n1620 = ~n265 & n1619;
  assign n1621 = n99 & ~n1620;
  assign n1622 = n25 & n35;
  assign n1623 = ~n230 & ~n1622;
  assign n1624 = n58 & ~n1623;
  assign n1625 = ~n1621 & ~n1624;
  assign n1626 = ~n166 & ~n481;
  assign n1627 = n102 & ~n1626;
  assign n1628 = n66 & n770;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = n1625 & n1629;
  assign n1631 = n878 & n1099;
  assign n1632 = n1630 & n1631;
  assign n1633 = n1618 & n1632;
  assign n1634 = ~n220 & ~n496;
  assign n1635 = ~n69 & n1634;
  assign n1636 = n23 & ~n1635;
  assign n1637 = n1252 & ~n1636;
  assign n1638 = n477 & n1637;
  assign n1639 = n988 & n1638;
  assign n1640 = n1633 & n1639;
  assign o_8_ = ~n1595 | ~n1640;
  assign n1642 = ~n232 & ~n679;
  assign n1643 = n99 & ~n1642;
  assign n1644 = n544 & ~n1643;
  assign n1645 = ~n438 & ~n664;
  assign n1646 = n117 & ~n1645;
  assign n1647 = n32 & ~n1619;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = n1088 & n1648;
  assign n1650 = n784 & n1649;
  assign n1651 = n1644 & n1650;
  assign n1652 = n102 & n329;
  assign n1653 = ~n344 & ~n1652;
  assign n1654 = ~n733 & n1653;
  assign n1655 = n177 & n203;
  assign n1656 = ~n126 & ~n378;
  assign n1657 = n114 & ~n1656;
  assign n1658 = ~n1655 & ~n1657;
  assign n1659 = ~n207 & ~n504;
  assign n1660 = n54 & ~n1659;
  assign n1661 = i_6_ & n1292;
  assign n1662 = n153 & n1661;
  assign n1663 = n95 & n427;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1660 & n1664;
  assign n1666 = n1658 & n1665;
  assign n1667 = ~n213 & ~n378;
  assign n1668 = ~n604 & n1667;
  assign n1669 = n41 & ~n1668;
  assign n1670 = ~n1419 & ~n1669;
  assign n1671 = n1666 & n1670;
  assign n1672 = n897 & n1671;
  assign n1673 = n1654 & n1672;
  assign n1674 = n1651 & n1673;
  assign n1675 = n1471 & n1674;
  assign n1676 = ~n643 & ~n806;
  assign n1677 = n1504 & n1676;
  assign n1678 = n89 & ~n1677;
  assign n1679 = ~n195 & ~n418;
  assign n1680 = ~n504 & n1679;
  assign n1681 = n122 & ~n1680;
  assign n1682 = ~n479 & ~n929;
  assign n1683 = n79 & ~n1682;
  assign n1684 = ~n56 & ~n118;
  assign n1685 = n58 & ~n1684;
  assign n1686 = ~n1683 & ~n1685;
  assign n1687 = ~n1681 & n1686;
  assign n1688 = ~n1678 & n1687;
  assign n1689 = n138 & n1688;
  assign n1690 = ~n168 & ~n531;
  assign n1691 = ~n49 & n1690;
  assign n1692 = n23 & ~n1691;
  assign n1693 = n1361 & ~n1692;
  assign n1694 = ~n420 & ~n424;
  assign n1695 = ~n90 & n1694;
  assign n1696 = n72 & ~n1695;
  assign n1697 = n507 & ~n1696;
  assign n1698 = n1693 & n1697;
  assign n1699 = n1593 & n1698;
  assign n1700 = n1689 & n1699;
  assign n1701 = n1268 & n1700;
  assign o_9_ = ~n1675 | ~n1701;
endmodule


