// Benchmark "x4" written by ABC on Tue May 16 16:07:54 2017

module x4 ( 
    z0, z1, a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z,
    a0, a1, a2, b0, b1, b2, c0, c1, c2, d0, d1, d2, e0, e1, e2, f0, f1, f2,
    g0, g1, g2, h0, h1, h2, i0, i1, i2, j1, j2, k0, k1, k2, l0, l1, l2, m0,
    m1, m2, n0, n1, n2, o0, o1, o2, p0, p1, p2, q0, q1, q2, r0, r1, r2, s0,
    s1, s2, t0, t1, t2, u0, u1, u2, v0, v1, v2, w0, w1, x0, x1, y0, y1,
    z2, z3, z4, a3, a4, a5, b3, b4, b5, c3, c4, c5, d3, d4, d5, e3, e4, e5,
    f3, f4, f5, g3, g4, g5, h3, h4, h5, i3, i4, i5, j3, j4, j5, k3, k4, k5,
    l3, l4, l5, m3, m4, m5, n3, n4, n5, o3, o4, o5, p3, p4, q3, q4, r3, r4,
    s3, s4, t3, t4, u3, u4, v3, v4, w2, w3, w4, x2, x3, x4, y2, y3, y4  );
  input  z0, z1, a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, a1, a2, b0, b1, b2, c0, c1, c2, d0, d1, d2, e0, e1, e2, f0,
    f1, f2, g0, g1, g2, h0, h1, h2, i0, i1, i2, j1, j2, k0, k1, k2, l0, l1,
    l2, m0, m1, m2, n0, n1, n2, o0, o1, o2, p0, p1, p2, q0, q1, q2, r0, r1,
    r2, s0, s1, s2, t0, t1, t2, u0, u1, u2, v0, v1, v2, w0, w1, x0, x1, y0,
    y1;
  output z2, z3, z4, a3, a4, a5, b3, b4, b5, c3, c4, c5, d3, d4, d5, e3, e4,
    e5, f3, f4, f5, g3, g4, g5, h3, h4, h5, i3, i4, i5, j3, j4, j5, k3, k4,
    k5, l3, l4, l5, m3, m4, m5, n3, n4, n5, o3, o4, o5, p3, p4, q3, q4, r3,
    r4, s3, s4, t3, t4, u3, u4, v3, v4, w2, w3, w4, x2, x3, x4, y2, y3, y4;
  wire n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250, n251,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n270, n271, n272, n273, n274, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n311, n312, n313, n314, n315, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n359, n360, n361, n362, n363, n365, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n395,
    n396, n397, n398, n399, n401, n402, n403, n404, n405, n406, n407, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n433, n434,
    n435, n436, n437, n438, n439, n440, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n478, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n492, n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n528, n530, n531, n532, n533, n534, n535, n536, n537,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n578, n580, n581, n582, n583, n584, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n631, n633, n634, n635, n636, n637, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n693, n695, n696, n697, n698, n699, n701, n702, n703,
    n704, n705, n706, n707, n709, n711, n712, n713, n714, n715, n717, n718,
    n719, n720, n721, n722, n723, n726, n727, n728, n729, n730, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n744, n745, n746, n747,
    n748, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n763, n764, n765, n766, n767, n770, n771, n772, n773, n774, n777, n778,
    n779, n780, n781, n784, n785, n786, n787, n788, n791, n792, n793, n794,
    n795, n798, n799, n800, n801, n802, n804, n805, n806, n807, n808, n809,
    n811, n812, n813, n814, n815, n817, n818, n819, n820, n821, n822, n824,
    n825, n826, n827, n828, n830, n831, n832, n833, n834, n836, n837, n838,
    n839, n840, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n859, n860, n861, n862, n863;
  assign n166 = ~q2 & ~r2;
  assign n167 = ~p2 & n166;
  assign n168 = ~n2 & o2;
  assign n169 = e1 & n168;
  assign n170 = n167 & n169;
  assign n171 = o2 & n167;
  assign n172 = n170 & ~n171;
  assign n173 = ~c1 & n172;
  assign n174 = p0 & n170;
  assign n175 = ~c1 & n174;
  assign n176 = ~e1 & n170;
  assign n177 = ~c1 & n176;
  assign n178 = n2 & n170;
  assign n179 = ~c1 & n178;
  assign n180 = g1 & ~n171;
  assign n181 = ~c1 & n180;
  assign n182 = g1 & p0;
  assign n183 = ~c1 & n182;
  assign n184 = ~e1 & g1;
  assign n185 = ~c1 & n184;
  assign n186 = g1 & n2;
  assign n187 = ~c1 & n186;
  assign n188 = ~n185 & ~n187;
  assign n189 = ~n183 & n188;
  assign n190 = ~n181 & n189;
  assign n191 = ~n179 & n190;
  assign n192 = ~n177 & n191;
  assign n193 = ~n175 & n192;
  assign z3 = n173 | ~n193;
  assign n195 = e1 & h2;
  assign n196 = g0 & ~h0;
  assign n197 = v2 & n196;
  assign n198 = m1 & n197;
  assign n199 = i & g0;
  assign n200 = v2 & n199;
  assign n201 = m1 & n200;
  assign n202 = h & g0;
  assign n203 = v2 & n202;
  assign n204 = m1 & n203;
  assign n205 = g & g0;
  assign n206 = v2 & n205;
  assign n207 = m1 & n206;
  assign n208 = ~n204 & ~n207;
  assign n209 = ~n201 & n208;
  assign n210 = ~n198 & n209;
  assign n211 = m1 & v2;
  assign n212 = ~i0 & n211;
  assign n213 = ~i & h0;
  assign n214 = ~h & n213;
  assign n215 = ~g & n214;
  assign n216 = g0 & n211;
  assign n217 = ~n215 & n216;
  assign n218 = e1 & ~m0;
  assign n219 = ~n217 & ~n218;
  assign n220 = ~i0 & ~m0;
  assign n221 = n210 & n220;
  assign n222 = n195 & n221;
  assign n223 = g0 & ~n215;
  assign n224 = n212 & n223;
  assign n225 = b0 & n224;
  assign n226 = ~i0 & n219;
  assign n227 = g2 & n226;
  assign n228 = ~n225 & ~n227;
  assign z4 = n222 | ~n228;
  assign n230 = q0 & n170;
  assign n231 = ~c1 & n230;
  assign n232 = h1 & ~n171;
  assign n233 = ~c1 & n232;
  assign n234 = h1 & q0;
  assign n235 = ~c1 & n234;
  assign n236 = ~e1 & h1;
  assign n237 = ~c1 & n236;
  assign n238 = h1 & n2;
  assign n239 = ~c1 & n238;
  assign n240 = ~n237 & ~n239;
  assign n241 = ~n235 & n240;
  assign n242 = ~n233 & n241;
  assign n243 = ~n179 & n242;
  assign n244 = ~n177 & n243;
  assign n245 = ~n231 & n244;
  assign a4 = n173 | ~n245;
  assign n247 = e1 & i2;
  assign n248 = n221 & n247;
  assign n249 = c0 & n224;
  assign n250 = h2 & n226;
  assign n251 = ~n249 & ~n250;
  assign a5 = n248 | ~n251;
  assign n253 = r0 & n170;
  assign n254 = ~c1 & n253;
  assign n255 = i1 & ~n171;
  assign n256 = ~c1 & n255;
  assign n257 = i1 & r0;
  assign n258 = ~c1 & n257;
  assign n259 = ~e1 & i1;
  assign n260 = ~c1 & n259;
  assign n261 = i1 & n2;
  assign n262 = ~c1 & n261;
  assign n263 = ~n260 & ~n262;
  assign n264 = ~n258 & n263;
  assign n265 = ~n256 & n264;
  assign n266 = ~n179 & n265;
  assign n267 = ~n177 & n266;
  assign n268 = ~n254 & n267;
  assign b4 = n173 | ~n268;
  assign n270 = e1 & j2;
  assign n271 = n221 & n270;
  assign n272 = d0 & n224;
  assign n273 = i2 & n226;
  assign n274 = ~n272 & ~n273;
  assign b5 = n271 | ~n274;
  assign n276 = h0 & ~t2;
  assign n277 = ~h0 & t2;
  assign n278 = ~i & ~q2;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~n276 & n279;
  assign n281 = ~p2 & r2;
  assign n282 = ~o2 & n281;
  assign n283 = n2 & n282;
  assign n284 = e1 & n2;
  assign n285 = ~o2 & n284;
  assign n286 = ~n278 & n285;
  assign n287 = n281 & n286;
  assign n288 = e1 & ~i0;
  assign n289 = n283 & n288;
  assign n290 = n280 & n289;
  assign n291 = ~i0 & s2;
  assign n292 = ~n287 & n291;
  assign c3 = n290 | n292;
  assign n294 = s0 & n170;
  assign n295 = ~c1 & n294;
  assign n296 = j1 & ~n171;
  assign n297 = ~c1 & n296;
  assign n298 = j1 & s0;
  assign n299 = ~c1 & n298;
  assign n300 = ~e1 & j1;
  assign n301 = ~c1 & n300;
  assign n302 = j1 & n2;
  assign n303 = ~c1 & n302;
  assign n304 = ~n301 & ~n303;
  assign n305 = ~n299 & n304;
  assign n306 = ~n297 & n305;
  assign n307 = ~n179 & n306;
  assign n308 = ~n177 & n307;
  assign n309 = ~n295 & n308;
  assign c4 = n173 | ~n309;
  assign n311 = e0 & g0;
  assign n312 = n212 & n311;
  assign n313 = ~n215 & n312;
  assign n314 = ~i0 & j2;
  assign n315 = n219 & n314;
  assign c5 = n313 | n315;
  assign n317 = ~h0 & m1;
  assign n318 = i & m1;
  assign n319 = h & m1;
  assign n320 = g & m1;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~n318 & n321;
  assign n323 = ~n317 & n322;
  assign n324 = ~f0 & ~k0;
  assign n325 = ~c1 & ~n324;
  assign n326 = ~k0 & ~v2;
  assign n327 = n325 & ~n326;
  assign n328 = ~c1 & v2;
  assign n329 = g0 & n328;
  assign n330 = n323 & n329;
  assign d3 = n327 | n330;
  assign n332 = t0 & n170;
  assign n333 = ~c1 & n332;
  assign n334 = k1 & ~n171;
  assign n335 = ~c1 & n334;
  assign n336 = k1 & t0;
  assign n337 = ~c1 & n336;
  assign n338 = ~e1 & k1;
  assign n339 = ~c1 & n338;
  assign n340 = k1 & n2;
  assign n341 = ~c1 & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = ~n337 & n342;
  assign n344 = ~n335 & n343;
  assign n345 = ~n179 & n344;
  assign n346 = ~n177 & n345;
  assign n347 = ~n333 & n346;
  assign d4 = n173 | ~n347;
  assign n349 = b & ~u0;
  assign n350 = k2 & n349;
  assign n351 = k2 & u2;
  assign n352 = ~c1 & ~n351;
  assign n353 = ~n350 & n352;
  assign n354 = n349 & n353;
  assign n355 = k2 & n353;
  assign n356 = u2 & n353;
  assign n357 = ~n355 & ~n356;
  assign d5 = n354 | ~n357;
  assign n359 = ~o2 & n167;
  assign n360 = ~c1 & l0;
  assign n361 = ~c1 & e1;
  assign n362 = n2 & n361;
  assign n363 = n359 & n362;
  assign e3 = n360 | n363;
  assign n365 = ~c1 & l1;
  assign e4 = n363 | n365;
  assign n367 = ~k2 & m2;
  assign n368 = ~k2 & ~l2;
  assign n369 = ~c1 & ~n368;
  assign n370 = ~n367 & n369;
  assign n371 = ~u2 & ~n349;
  assign n372 = n349 & n371;
  assign n373 = n370 & n372;
  assign n374 = u2 & n371;
  assign n375 = n370 & n374;
  assign n376 = l2 & n371;
  assign n377 = n370 & n376;
  assign n378 = ~l2 & n349;
  assign n379 = n370 & n378;
  assign n380 = ~k2 & n349;
  assign n381 = n370 & n380;
  assign n382 = ~l2 & u2;
  assign n383 = n370 & n382;
  assign n384 = ~k2 & u2;
  assign n385 = n370 & n384;
  assign n386 = ~k2 & l2;
  assign n387 = n370 & n386;
  assign n388 = ~n385 & ~n387;
  assign n389 = ~n383 & n388;
  assign n390 = ~n381 & n389;
  assign n391 = ~n379 & n390;
  assign n392 = ~n377 & n391;
  assign n393 = ~n375 & n392;
  assign e5 = n373 | ~n393;
  assign n395 = ~i0 & v2;
  assign n396 = g0 & n395;
  assign n397 = ~n220 & ~n396;
  assign n398 = g0 & v2;
  assign n399 = n323 & n398;
  assign f3 = n397 | n399;
  assign n401 = ~i0 & ~n398;
  assign n402 = l2 & m2;
  assign n403 = ~h & ~k2;
  assign n404 = ~g & n403;
  assign n405 = n402 & n404;
  assign n406 = n401 & n405;
  assign n407 = m1 & n401;
  assign f4 = n406 | n407;
  assign n409 = ~l2 & ~m2;
  assign n410 = ~k2 & ~m2;
  assign n411 = ~c1 & ~n386;
  assign n412 = ~n410 & n411;
  assign n413 = ~n409 & n412;
  assign n414 = n372 & n413;
  assign n415 = n374 & n413;
  assign n416 = m2 & n371;
  assign n417 = n413 & n416;
  assign n418 = ~m2 & n349;
  assign n419 = n413 & n418;
  assign n420 = n378 & n413;
  assign n421 = ~m2 & u2;
  assign n422 = n413 & n421;
  assign n423 = n382 & n413;
  assign n424 = ~l2 & m2;
  assign n425 = n413 & n424;
  assign n426 = ~n423 & ~n425;
  assign n427 = ~n422 & n426;
  assign n428 = ~n420 & n427;
  assign n429 = ~n419 & n428;
  assign n430 = ~n417 & n429;
  assign n431 = ~n415 & n430;
  assign f5 = n414 | ~n431;
  assign n433 = ~n0 & ~n167;
  assign n434 = ~e1 & ~n0;
  assign n435 = ~n0 & o2;
  assign n436 = ~n0 & ~n2;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n434 & n437;
  assign n439 = ~n433 & n438;
  assign n440 = ~c1 & ~i0;
  assign g3 = n439 & n440;
  assign n442 = ~n198 & n208;
  assign n443 = e1 & ~o1;
  assign n444 = h & n398;
  assign n445 = m1 & n444;
  assign n446 = g & n398;
  assign n447 = m1 & n446;
  assign n448 = ~h0 & v2;
  assign n449 = g0 & n448;
  assign n450 = m1 & n449;
  assign n451 = ~n218 & ~n450;
  assign n452 = ~n447 & n451;
  assign n453 = ~n445 & n452;
  assign n454 = g0 & ~i0;
  assign n455 = i & n454;
  assign n456 = n211 & n455;
  assign n457 = n220 & n443;
  assign n458 = n442 & n457;
  assign n459 = ~i0 & n1;
  assign n460 = n453 & n459;
  assign n461 = ~n458 & ~n460;
  assign g4 = n456 | ~n461;
  assign n463 = ~k2 & n2;
  assign n464 = l2 & n463;
  assign n465 = m2 & n464;
  assign n466 = d1 & n2;
  assign n467 = ~c1 & ~n284;
  assign n468 = ~n466 & n467;
  assign n469 = ~n465 & n468;
  assign n470 = ~k2 & n402;
  assign n471 = n469 & n470;
  assign n472 = d1 & n469;
  assign n473 = e1 & n469;
  assign n474 = n2 & n469;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n472 & n475;
  assign g5 = n471 | ~n476;
  assign n478 = ~c1 & o0;
  assign h3 = ~i0 & n478;
  assign n480 = e1 & n220;
  assign n481 = p1 & n480;
  assign n482 = ~i0 & ~o1;
  assign n483 = p1 & n482;
  assign n484 = ~e1 & ~i0;
  assign n485 = ~o1 & n484;
  assign n486 = ~i0 & m0;
  assign n487 = ~o1 & n486;
  assign n488 = ~n485 & ~n487;
  assign n489 = ~n483 & n488;
  assign n490 = ~n481 & n489;
  assign h4 = n217 | n490;
  assign n492 = ~n2 & ~o2;
  assign n493 = ~c1 & ~n492;
  assign n494 = ~d1 & ~e1;
  assign n495 = m2 & n386;
  assign n496 = n494 & ~n495;
  assign n497 = n470 & n496;
  assign n498 = n493 & n497;
  assign n499 = d1 & n496;
  assign n500 = n493 & n499;
  assign n501 = e1 & n496;
  assign n502 = n493 & n501;
  assign n503 = o2 & n496;
  assign n504 = n493 & n503;
  assign n505 = ~o2 & n470;
  assign n506 = n493 & n505;
  assign n507 = ~n2 & n470;
  assign n508 = n493 & n507;
  assign n509 = d1 & ~o2;
  assign n510 = n493 & n509;
  assign n511 = d1 & ~n2;
  assign n512 = n493 & n511;
  assign n513 = e1 & ~o2;
  assign n514 = n493 & n513;
  assign n515 = e1 & ~n2;
  assign n516 = n493 & n515;
  assign n517 = n168 & n493;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n514 & n518;
  assign n520 = ~n512 & n519;
  assign n521 = ~n510 & n520;
  assign n522 = ~n508 & n521;
  assign n523 = ~n506 & n522;
  assign n524 = ~n504 & n523;
  assign n525 = ~n502 & n524;
  assign n526 = ~n500 & n525;
  assign h5 = n498 | ~n526;
  assign n528 = ~c1 & p0;
  assign i3 = ~i0 & n528;
  assign n530 = e1 & q1;
  assign n531 = n220 & n530;
  assign n532 = n210 & n531;
  assign n533 = k & n223;
  assign n534 = n212 & n533;
  assign n535 = ~i0 & p1;
  assign n536 = n219 & n535;
  assign n537 = ~n534 & ~n536;
  assign i4 = n532 | ~n537;
  assign n539 = ~o2 & ~p2;
  assign n540 = ~n2 & ~p2;
  assign n541 = ~c1 & ~n540;
  assign n542 = ~n539 & n541;
  assign n543 = n497 & n542;
  assign n544 = n499 & n542;
  assign n545 = n501 & n542;
  assign n546 = p2 & n496;
  assign n547 = n542 & n546;
  assign n548 = ~p2 & n470;
  assign n549 = n542 & n548;
  assign n550 = n505 & n542;
  assign n551 = n507 & n542;
  assign n552 = d1 & ~p2;
  assign n553 = n542 & n552;
  assign n554 = n509 & n542;
  assign n555 = n511 & n542;
  assign n556 = e1 & ~p2;
  assign n557 = n542 & n556;
  assign n558 = n513 & n542;
  assign n559 = n515 & n542;
  assign n560 = ~o2 & p2;
  assign n561 = n542 & n560;
  assign n562 = ~n2 & p2;
  assign n563 = n542 & n562;
  assign n564 = ~n561 & ~n563;
  assign n565 = ~n559 & n564;
  assign n566 = ~n558 & n565;
  assign n567 = ~n557 & n566;
  assign n568 = ~n555 & n567;
  assign n569 = ~n554 & n568;
  assign n570 = ~n553 & n569;
  assign n571 = ~n551 & n570;
  assign n572 = ~n550 & n571;
  assign n573 = ~n549 & n572;
  assign n574 = ~n547 & n573;
  assign n575 = ~n545 & n574;
  assign n576 = ~n544 & n575;
  assign i5 = n543 | ~n576;
  assign n578 = ~c1 & q0;
  assign j3 = ~i0 & n578;
  assign n580 = e1 & r1;
  assign n581 = n221 & n580;
  assign n582 = l & n224;
  assign n583 = q1 & n226;
  assign n584 = ~n582 & ~n583;
  assign j4 = n581 | ~n584;
  assign n586 = ~p2 & ~q2;
  assign n587 = ~o2 & ~q2;
  assign n588 = ~n2 & ~q2;
  assign n589 = ~c1 & ~n588;
  assign n590 = ~n587 & n589;
  assign n591 = ~n586 & n590;
  assign n592 = p2 & q2;
  assign n593 = n497 & n591;
  assign n594 = n470 & ~n592;
  assign n595 = n591 & n594;
  assign n596 = n507 & n591;
  assign n597 = n505 & n591;
  assign n598 = n499 & n591;
  assign n599 = d1 & ~n592;
  assign n600 = n591 & n599;
  assign n601 = n511 & n591;
  assign n602 = n509 & n591;
  assign n603 = n501 & n591;
  assign n604 = e1 & ~n592;
  assign n605 = n591 & n604;
  assign n606 = n515 & n591;
  assign n607 = n513 & n591;
  assign n608 = q2 & n496;
  assign n609 = n591 & n608;
  assign n610 = q2 & ~n592;
  assign n611 = n591 & n610;
  assign n612 = ~n2 & q2;
  assign n613 = n591 & n612;
  assign n614 = ~o2 & q2;
  assign n615 = n591 & n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n611 & n616;
  assign n618 = ~n609 & n617;
  assign n619 = ~n607 & n618;
  assign n620 = ~n606 & n619;
  assign n621 = ~n605 & n620;
  assign n622 = ~n603 & n621;
  assign n623 = ~n602 & n622;
  assign n624 = ~n601 & n623;
  assign n625 = ~n600 & n624;
  assign n626 = ~n598 & n625;
  assign n627 = ~n597 & n626;
  assign n628 = ~n596 & n627;
  assign n629 = ~n595 & n628;
  assign j5 = n593 | ~n629;
  assign n631 = ~c1 & r0;
  assign k3 = ~i0 & n631;
  assign n633 = e1 & s1;
  assign n634 = n221 & n633;
  assign n635 = m & n224;
  assign n636 = r1 & n226;
  assign n637 = ~n635 & ~n636;
  assign k4 = n634 | ~n637;
  assign n639 = o2 & n592;
  assign n640 = n2 & n639;
  assign n641 = q2 & r2;
  assign n642 = p2 & n641;
  assign n643 = n470 & ~n642;
  assign n644 = n640 & n643;
  assign n645 = ~c1 & n644;
  assign n646 = d1 & ~n642;
  assign n647 = n640 & n646;
  assign n648 = ~c1 & n647;
  assign n649 = e1 & ~n642;
  assign n650 = n640 & n649;
  assign n651 = ~c1 & n650;
  assign n652 = n497 & n640;
  assign n653 = ~c1 & n652;
  assign n654 = n499 & n640;
  assign n655 = ~c1 & n654;
  assign n656 = n501 & n640;
  assign n657 = ~c1 & n656;
  assign n658 = n505 & n640;
  assign n659 = ~c1 & n658;
  assign n660 = n507 & n640;
  assign n661 = ~c1 & n660;
  assign n662 = n509 & n640;
  assign n663 = ~c1 & n662;
  assign n664 = n511 & n640;
  assign n665 = ~c1 & n664;
  assign n666 = n513 & n640;
  assign n667 = ~c1 & n666;
  assign n668 = n515 & n640;
  assign n669 = ~c1 & n668;
  assign n670 = r2 & ~n642;
  assign n671 = ~c1 & n670;
  assign n672 = r2 & n496;
  assign n673 = ~c1 & n672;
  assign n674 = ~o2 & r2;
  assign n675 = ~c1 & n674;
  assign n676 = ~n2 & r2;
  assign n677 = ~c1 & n676;
  assign n678 = ~n675 & ~n677;
  assign n679 = ~n673 & n678;
  assign n680 = ~n671 & n679;
  assign n681 = ~n669 & n680;
  assign n682 = ~n667 & n681;
  assign n683 = ~n665 & n682;
  assign n684 = ~n663 & n683;
  assign n685 = ~n661 & n684;
  assign n686 = ~n659 & n685;
  assign n687 = ~n657 & n686;
  assign n688 = ~n655 & n687;
  assign n689 = ~n653 & n688;
  assign n690 = ~n651 & n689;
  assign n691 = ~n648 & n690;
  assign k5 = n645 | ~n691;
  assign n693 = ~c1 & s0;
  assign l3 = ~i0 & n693;
  assign n695 = e1 & t1;
  assign n696 = n221 & n695;
  assign n697 = n & n224;
  assign n698 = s1 & n226;
  assign n699 = ~n697 & ~n698;
  assign l4 = n696 | ~n699;
  assign n701 = n1 & n480;
  assign n702 = b1 & ~i0;
  assign n703 = n1 & n702;
  assign n704 = b1 & n484;
  assign n705 = b1 & n486;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n703 & n706;
  assign l5 = n701 | ~n707;
  assign n709 = ~c1 & t0;
  assign m3 = ~i0 & n709;
  assign n711 = e1 & u1;
  assign n712 = n221 & n711;
  assign n713 = o & n224;
  assign n714 = t1 & n226;
  assign n715 = ~n713 & ~n714;
  assign m4 = n712 | ~n715;
  assign n717 = s2 & n365;
  assign n718 = ~t2 & n717;
  assign n719 = ~c1 & ~s2;
  assign n720 = t2 & n719;
  assign n721 = ~c1 & ~l1;
  assign n722 = t2 & n721;
  assign n723 = ~n720 & ~n722;
  assign m5 = n718 | ~n723;
  assign n3 = b & ~i0;
  assign n726 = e1 & v1;
  assign n727 = n221 & n726;
  assign n728 = p & n224;
  assign n729 = u1 & n226;
  assign n730 = ~n728 & ~n729;
  assign n4 = n727 | ~n730;
  assign n732 = u0 & ~u2;
  assign n733 = ~b & ~u2;
  assign n734 = ~i0 & ~n733;
  assign n735 = ~n732 & n734;
  assign n736 = n349 & n735;
  assign n737 = k2 & n735;
  assign n738 = ~l2 & n735;
  assign n739 = ~m2 & n735;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n737 & n740;
  assign n5 = n736 | ~n741;
  assign o3 = a & ~i0;
  assign n744 = e1 & w1;
  assign n745 = n221 & n744;
  assign n746 = q & n224;
  assign n747 = v1 & n226;
  assign n748 = ~n746 & ~n747;
  assign o4 = n745 | ~n748;
  assign n750 = ~p2 & q2;
  assign n751 = ~o2 & n750;
  assign n752 = r2 & n751;
  assign n753 = i & ~p2;
  assign n754 = ~o2 & n753;
  assign n755 = r2 & n754;
  assign n756 = ~n752 & ~n755;
  assign n757 = n284 & ~n756;
  assign n758 = n401 & n757;
  assign n759 = ~f0 & v2;
  assign n760 = n401 & n759;
  assign o5 = n758 | n760;
  assign p3 = ~i0 & v0;
  assign n763 = e1 & x1;
  assign n764 = n221 & n763;
  assign n765 = r & n224;
  assign n766 = w1 & n226;
  assign n767 = ~n765 & ~n766;
  assign p4 = n764 | ~n767;
  assign q3 = ~i0 & w0;
  assign n770 = e1 & y1;
  assign n771 = n221 & n770;
  assign n772 = s & n224;
  assign n773 = x1 & n226;
  assign n774 = ~n772 & ~n773;
  assign q4 = n771 | ~n774;
  assign r3 = ~i0 & x0;
  assign n777 = z1 & e1;
  assign n778 = n221 & n777;
  assign n779 = t & n224;
  assign n780 = y1 & n226;
  assign n781 = ~n779 & ~n780;
  assign r4 = n778 | ~n781;
  assign s3 = ~i0 & y0;
  assign n784 = a2 & e1;
  assign n785 = n221 & n784;
  assign n786 = u & n224;
  assign n787 = z1 & n226;
  assign n788 = ~n786 & ~n787;
  assign s4 = n785 | ~n788;
  assign t3 = z0 & ~i0;
  assign n791 = b2 & e1;
  assign n792 = n221 & n791;
  assign n793 = v & n224;
  assign n794 = a2 & n226;
  assign n795 = ~n793 & ~n794;
  assign t4 = n792 | ~n795;
  assign u3 = a1 & ~i0;
  assign n798 = c2 & e1;
  assign n799 = n221 & n798;
  assign n800 = w & n224;
  assign n801 = b2 & n226;
  assign n802 = ~n800 & ~n801;
  assign u4 = n799 | ~n802;
  assign n804 = ~f0 & ~i0;
  assign n805 = ~i0 & ~v2;
  assign n806 = ~n804 & ~n805;
  assign n807 = n282 & n284;
  assign n808 = ~n278 & n807;
  assign n809 = ~n399 & ~n806;
  assign v3 = n808 | ~n809;
  assign n811 = d2 & e1;
  assign n812 = n221 & n811;
  assign n813 = x & n224;
  assign n814 = c2 & n226;
  assign n815 = ~n813 & ~n814;
  assign v4 = n812 | ~n815;
  assign n817 = ~g & ~h;
  assign n818 = ~i & n817;
  assign n819 = h0 & n818;
  assign n820 = ~g0 & i0;
  assign n821 = ~m1 & n820;
  assign n822 = ~n819 & n821;
  assign w3 = v2 & n822;
  assign n824 = e1 & e2;
  assign n825 = n221 & n824;
  assign n826 = y & n224;
  assign n827 = d2 & n226;
  assign n828 = ~n826 & ~n827;
  assign w4 = n825 | ~n828;
  assign n830 = ~c1 & ~k2;
  assign n831 = l2 & n830;
  assign n832 = m2 & n831;
  assign n833 = ~c1 & d1;
  assign n834 = ~n361 & ~n833;
  assign x3 = n832 | ~n834;
  assign n836 = e1 & f2;
  assign n837 = n221 & n836;
  assign n838 = z & n224;
  assign n839 = e2 & n226;
  assign n840 = ~n838 & ~n839;
  assign x4 = n837 | ~n840;
  assign n842 = o0 & n170;
  assign n843 = ~c1 & n842;
  assign n844 = f1 & ~n171;
  assign n845 = ~c1 & n844;
  assign n846 = f1 & o0;
  assign n847 = ~c1 & n846;
  assign n848 = ~e1 & f1;
  assign n849 = ~c1 & n848;
  assign n850 = f1 & n2;
  assign n851 = ~c1 & n850;
  assign n852 = ~n849 & ~n851;
  assign n853 = ~n847 & n852;
  assign n854 = ~n845 & n853;
  assign n855 = ~n179 & n854;
  assign n856 = ~n177 & n855;
  assign n857 = ~n843 & n856;
  assign y3 = n173 | ~n857;
  assign n859 = e1 & g2;
  assign n860 = n221 & n859;
  assign n861 = a0 & n224;
  assign n862 = f2 & n226;
  assign n863 = ~n861 & ~n862;
  assign y4 = n860 | ~n863;
  assign z2 = ~i1;
  assign a3 = ~j1;
  assign b3 = ~k1;
  assign w2 = ~f1;
  assign x2 = ~g1;
  assign y2 = ~h1;
endmodule


