// Benchmark "TOP" written by ABC on Sun Apr 24 20:32:48 2016

module TOP ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2;
  wire n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012;
  assign n29 = ~m & ~n;
  assign n30 = ~h & i;
  assign n31 = ~j & l;
  assign n32 = ~k & ~n31;
  assign n33 = n30 & ~n32;
  assign n34 = h & k;
  assign n35 = i & j;
  assign n36 = l & n35;
  assign n37 = n34 & ~n36;
  assign n38 = i & k;
  assign n39 = h & j;
  assign n40 = ~n38 & n39;
  assign n41 = ~n37 & ~n40;
  assign n42 = ~n33 & n41;
  assign n43 = n29 & ~n42;
  assign n44 = e & ~f;
  assign n45 = c & n44;
  assign n46 = n43 & n45;
  assign n47 = d & n46;
  assign n48 = a & d;
  assign n49 = b & n48;
  assign n50 = m & ~n;
  assign n51 = ~l & ~n39;
  assign n52 = h & ~i;
  assign n53 = l & ~n52;
  assign n54 = ~h & j;
  assign n55 = ~n30 & ~n54;
  assign n56 = n53 & n55;
  assign n57 = ~n51 & ~n56;
  assign n58 = ~i & j;
  assign n59 = ~k & n58;
  assign n60 = i & ~j;
  assign n61 = k & n60;
  assign n62 = ~n59 & ~n61;
  assign n63 = k & ~l;
  assign n64 = ~n58 & n63;
  assign n65 = j & ~k;
  assign n66 = l & n65;
  assign n67 = ~n64 & ~n66;
  assign n68 = n62 & n67;
  assign n69 = ~n57 & n68;
  assign n70 = n50 & ~n69;
  assign n71 = ~e & g;
  assign n72 = n70 & n71;
  assign n73 = ~n32 & n50;
  assign n74 = ~g & h;
  assign n75 = ~e & n74;
  assign n76 = n73 & n75;
  assign n77 = ~n72 & ~n76;
  assign n78 = n49 & ~n77;
  assign n79 = b & c;
  assign n80 = e & n79;
  assign n81 = ~m & n;
  assign n82 = ~n32 & n81;
  assign n83 = ~f & n30;
  assign n84 = n82 & n83;
  assign n85 = ~j & ~k;
  assign n86 = k & n36;
  assign n87 = ~m & ~n86;
  assign n88 = ~n85 & n87;
  assign n89 = n & n88;
  assign n90 = ~f & h;
  assign n91 = n89 & n90;
  assign n92 = ~n84 & ~n91;
  assign n93 = n80 & ~n92;
  assign n94 = ~n78 & ~n93;
  assign n95 = ~n47 & n94;
  assign n96 = e & g;
  assign n97 = n70 & n96;
  assign n98 = e & n74;
  assign n99 = n73 & n98;
  assign n100 = ~n97 & ~n99;
  assign n101 = c & ~d;
  assign n102 = a & n101;
  assign n103 = ~n100 & n102;
  assign n104 = b & n103;
  assign n105 = g & n30;
  assign n106 = n82 & n105;
  assign n107 = g & h;
  assign n108 = n89 & n107;
  assign n109 = ~n106 & ~n108;
  assign n110 = ~d & ~e;
  assign n111 = n79 & n110;
  assign n112 = ~n109 & n111;
  assign n113 = f & n81;
  assign n114 = n33 & n113;
  assign n115 = f & h;
  assign n116 = n89 & n115;
  assign n117 = ~n114 & ~n116;
  assign n118 = b & d;
  assign n119 = ~e & n118;
  assign n120 = ~n117 & n119;
  assign n121 = ~n112 & ~n120;
  assign n122 = c & d;
  assign n123 = b & ~n122;
  assign n124 = g & ~n110;
  assign n125 = ~n117 & n124;
  assign n126 = n123 & n125;
  assign n127 = n121 & ~n126;
  assign n128 = ~n104 & n127;
  assign n129 = ~c & d;
  assign n130 = e & ~n129;
  assign n131 = ~g & n81;
  assign n132 = n33 & n131;
  assign n133 = n74 & n89;
  assign n134 = ~n132 & ~n133;
  assign n135 = b & f;
  assign n136 = ~n134 & n135;
  assign n137 = ~n130 & n136;
  assign n138 = ~l & n50;
  assign n139 = ~n38 & ~n39;
  assign n140 = g & ~n139;
  assign n141 = n138 & n140;
  assign n142 = k & n50;
  assign n143 = n74 & n142;
  assign n144 = g & n58;
  assign n145 = ~k & n50;
  assign n146 = n144 & n145;
  assign n147 = ~n143 & ~n146;
  assign n148 = ~n141 & n147;
  assign n149 = l & n50;
  assign n150 = g & ~n65;
  assign n151 = h & ~j;
  assign n152 = ~g & ~n151;
  assign n153 = ~n150 & ~n152;
  assign n154 = ~n105 & ~n144;
  assign n155 = ~i & n107;
  assign n156 = n154 & ~n155;
  assign n157 = ~n153 & n156;
  assign n158 = n149 & ~n157;
  assign n159 = n60 & n142;
  assign n160 = g & n159;
  assign n161 = n50 & n63;
  assign n162 = ~j & n161;
  assign n163 = g & n162;
  assign n164 = ~n160 & ~n163;
  assign n165 = ~n158 & n164;
  assign n166 = n148 & n165;
  assign n167 = ~a & b;
  assign n168 = e & n167;
  assign n169 = b & ~c;
  assign n170 = ~d & e;
  assign n171 = a & n170;
  assign n172 = n169 & n171;
  assign n173 = ~n168 & ~n172;
  assign n174 = ~n166 & ~n173;
  assign n175 = ~n34 & ~n139;
  assign n176 = n30 & n31;
  assign n177 = ~n37 & ~n176;
  assign n178 = ~n175 & n177;
  assign n179 = n29 & ~n178;
  assign n180 = c & f;
  assign n181 = d & e;
  assign n182 = n180 & ~n181;
  assign n183 = n179 & n182;
  assign n184 = ~n174 & ~n183;
  assign n185 = ~n137 & n184;
  assign n186 = n128 & n185;
  assign r2 = ~n95 | ~n186;
  assign n188 = a & c;
  assign n189 = ~b & n188;
  assign n190 = ~n166 & n181;
  assign n191 = f & n74;
  assign n192 = n73 & n191;
  assign n193 = f & g;
  assign n194 = n70 & n193;
  assign n195 = ~n192 & ~n194;
  assign n196 = ~e & ~n195;
  assign n197 = ~n190 & ~n196;
  assign n198 = n189 & ~n197;
  assign n199 = ~e & n180;
  assign n200 = ~n134 & n199;
  assign n201 = f & n129;
  assign n202 = n179 & n201;
  assign n203 = f & n43;
  assign n204 = ~e & n122;
  assign n205 = n203 & n204;
  assign n206 = ~n202 & ~n205;
  assign n207 = ~b & c;
  assign n208 = n71 & n101;
  assign n209 = ~n207 & ~n208;
  assign n210 = n113 & ~n178;
  assign n211 = ~n209 & n210;
  assign n212 = c & n120;
  assign n213 = ~n211 & ~n212;
  assign n214 = n206 & n213;
  assign n215 = ~n200 & n214;
  assign n216 = ~n198 & n215;
  assign n217 = n50 & ~n63;
  assign n218 = n58 & n217;
  assign n219 = n50 & ~n51;
  assign n220 = ~n53 & n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = n50 & ~n67;
  assign n223 = n30 & n149;
  assign n224 = ~n222 & ~n223;
  assign n225 = n221 & n224;
  assign n226 = g & ~n225;
  assign n227 = ~n160 & ~n226;
  assign n228 = e & ~n227;
  assign n229 = ~n99 & ~n228;
  assign n230 = d & n167;
  assign n231 = ~n229 & n230;
  assign n232 = ~c & n48;
  assign n233 = ~n44 & ~n227;
  assign n234 = ~n76 & ~n192;
  assign n235 = ~n233 & n234;
  assign n236 = n232 & ~n235;
  assign n237 = n95 & ~n236;
  assign n238 = ~n231 & n237;
  assign s2 = ~n216 | ~n238;
  assign n240 = f & ~n227;
  assign n241 = ~n192 & ~n240;
  assign n242 = d & ~e;
  assign n243 = ~n167 & ~n242;
  assign n244 = ~a & n242;
  assign n245 = ~n243 & ~n244;
  assign n246 = ~n241 & n245;
  assign n247 = ~n117 & n207;
  assign n248 = e & n247;
  assign n249 = ~n93 & ~n248;
  assign n250 = n92 & n109;
  assign n251 = b & n170;
  assign n252 = ~n250 & n251;
  assign n253 = e & n101;
  assign n254 = e & n129;
  assign n255 = ~n253 & ~n254;
  assign n256 = n203 & ~n255;
  assign n257 = n45 & n179;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~n252 & n258;
  assign n260 = n249 & n259;
  assign n261 = f & n103;
  assign n262 = n260 & ~n261;
  assign n263 = ~n246 & n262;
  assign n264 = a & ~n195;
  assign n265 = ~d & ~n169;
  assign n266 = ~n118 & ~n265;
  assign n267 = n264 & n266;
  assign n268 = ~f & ~n109;
  assign n269 = n129 & n268;
  assign n270 = n210 & n254;
  assign n271 = ~n269 & ~n270;
  assign n272 = b & ~n271;
  assign n273 = ~n267 & ~n272;
  assign t2 = ~n263 | ~n273;
  assign n275 = n98 & n102;
  assign n276 = ~a & d;
  assign n277 = ~n243 & ~n276;
  assign n278 = ~c & ~d;
  assign n279 = ~b & n278;
  assign n280 = a & ~n79;
  assign n281 = ~n279 & n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = f & ~n282;
  assign n284 = ~e & n129;
  assign n285 = ~n118 & ~n130;
  assign n286 = ~f & ~n285;
  assign n287 = ~n284 & ~n286;
  assign n288 = a & ~n287;
  assign n289 = ~n283 & ~n288;
  assign n290 = n74 & ~n289;
  assign n291 = ~n275 & ~n290;
  assign n292 = ~n32 & ~n291;
  assign n293 = g & ~n289;
  assign n294 = n96 & n102;
  assign n295 = ~n293 & ~n294;
  assign n296 = n63 & n293;
  assign n297 = ~n66 & ~n296;
  assign n298 = ~n295 & ~n297;
  assign n299 = ~n292 & ~n298;
  assign n300 = i & ~n;
  assign n301 = m & n300;
  assign n302 = ~n299 & n301;
  assign n303 = i & l;
  assign n304 = m & n303;
  assign n305 = ~h & n304;
  assign n306 = n293 & n305;
  assign n307 = k & ~m;
  assign n308 = n105 & n307;
  assign n309 = f & n308;
  assign n310 = g & n115;
  assign n311 = n88 & n310;
  assign n312 = ~n309 & ~n311;
  assign n313 = n253 & ~n312;
  assign n314 = b & n44;
  assign n315 = ~n168 & ~n314;
  assign n316 = n153 & n304;
  assign n317 = ~l & m;
  assign n318 = h & i;
  assign n319 = j & n318;
  assign n320 = g & n319;
  assign n321 = n317 & n320;
  assign n322 = ~n316 & ~n321;
  assign n323 = ~n315 & ~n322;
  assign n324 = ~n313 & ~n323;
  assign n325 = n317 & n319;
  assign n326 = ~n295 & n325;
  assign n327 = n324 & ~n326;
  assign n328 = ~n306 & n327;
  assign n329 = ~n & ~n328;
  assign n330 = n159 & n294;
  assign n331 = a & n284;
  assign n332 = ~n283 & n315;
  assign n333 = ~n331 & n332;
  assign n334 = n160 & ~n333;
  assign n335 = ~f & g;
  assign n336 = n159 & n335;
  assign n337 = a & ~n285;
  assign n338 = n336 & n337;
  assign n339 = ~n334 & ~n338;
  assign n340 = ~n330 & n339;
  assign n341 = ~n45 & ~n201;
  assign n342 = ~n284 & n341;
  assign n343 = ~n199 & n342;
  assign n344 = n43 & ~n343;
  assign n345 = ~n120 & ~n344;
  assign n346 = g & ~n345;
  assign n347 = l & ~m;
  assign n348 = ~n & n347;
  assign n349 = n253 & n348;
  assign n350 = ~j & n30;
  assign n351 = n193 & n350;
  assign n352 = n349 & n351;
  assign n353 = ~g & n318;
  assign n354 = ~n315 & n353;
  assign n355 = n142 & n354;
  assign n356 = ~n352 & ~n355;
  assign n357 = i & n161;
  assign n358 = ~n223 & ~n357;
  assign n359 = g & ~n315;
  assign n360 = ~n294 & ~n359;
  assign n361 = ~n358 & ~n360;
  assign n362 = f & n207;
  assign n363 = ~e & n207;
  assign n364 = b & e;
  assign n365 = ~n180 & n364;
  assign n366 = ~n363 & ~n365;
  assign n367 = ~n111 & n366;
  assign n368 = ~n362 & n367;
  assign n369 = ~n109 & ~n368;
  assign n370 = ~n361 & ~n369;
  assign n371 = n356 & n370;
  assign n372 = ~n346 & n371;
  assign n373 = n340 & n372;
  assign n374 = ~n329 & n373;
  assign u2 = n302 | ~n374;
  assign n376 = ~j & n149;
  assign n377 = ~n293 & n360;
  assign n378 = n52 & ~n377;
  assign n379 = n376 & n378;
  assign n380 = n135 & ~n170;
  assign n381 = ~n80 & ~n380;
  assign n382 = n74 & ~n381;
  assign n383 = n90 & n251;
  assign n384 = n115 & n119;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n382 & n385;
  assign n387 = n & ~n386;
  assign n388 = ~e & n278;
  assign n389 = n123 & ~n388;
  assign n390 = ~n314 & ~n389;
  assign n391 = ~n363 & n390;
  assign n392 = n & n391;
  assign n393 = ~n & ~n284;
  assign n394 = ~n392 & ~n393;
  assign n395 = n107 & n394;
  assign n396 = ~n387 & ~n395;
  assign n397 = n307 & ~n396;
  assign n398 = ~g & n180;
  assign n399 = ~n182 & ~n398;
  assign n400 = n341 & n399;
  assign n401 = n29 & ~n400;
  assign n402 = n113 & n207;
  assign n403 = ~n401 & ~n402;
  assign n404 = n34 & ~n403;
  assign n405 = ~n397 & ~n404;
  assign n406 = ~n35 & ~n405;
  assign n407 = l & n58;
  assign n408 = ~n30 & ~n407;
  assign n409 = n142 & ~n408;
  assign n410 = ~n162 & ~n409;
  assign n411 = ~n295 & ~n410;
  assign n412 = ~n406 & ~n411;
  assign n413 = ~n379 & n412;
  assign n414 = j & n145;
  assign n415 = h & ~n295;
  assign n416 = n107 & n168;
  assign n417 = ~n415 & ~n416;
  assign n418 = n414 & ~n417;
  assign n419 = n107 & ~n391;
  assign n420 = n386 & ~n419;
  assign n421 = n81 & ~n420;
  assign n422 = n107 & n284;
  assign n423 = n29 & n422;
  assign n424 = ~n421 & ~n423;
  assign n425 = n65 & ~n424;
  assign n426 = n39 & ~n403;
  assign n427 = ~k & n426;
  assign n428 = ~n425 & ~n427;
  assign n429 = i & ~n428;
  assign n430 = ~n418 & ~n429;
  assign n431 = k & n149;
  assign n432 = n144 & n431;
  assign n433 = n105 & n142;
  assign n434 = ~n163 & ~n433;
  assign n435 = ~n432 & n434;
  assign n436 = ~n315 & ~n435;
  assign n437 = n340 & ~n436;
  assign n438 = n430 & n437;
  assign n2 = ~n413 | ~n438;
  assign n440 = n142 & ~n291;
  assign n441 = n308 & n394;
  assign n442 = n83 & n251;
  assign n443 = ~e & f;
  assign n444 = ~h & n443;
  assign n445 = n118 & n444;
  assign n446 = ~g & ~h;
  assign n447 = ~n381 & n446;
  assign n448 = ~n445 & ~n447;
  assign n449 = i & ~n448;
  assign n450 = ~n442 & ~n449;
  assign n451 = n81 & ~n450;
  assign n452 = k & n451;
  assign n453 = ~n441 & ~n452;
  assign n454 = ~n440 & n453;
  assign n455 = n60 & n397;
  assign n456 = ~i & n31;
  assign n457 = n142 & n456;
  assign n458 = n50 & ~n62;
  assign n459 = ~n457 & ~n458;
  assign n460 = n415 & ~n459;
  assign n461 = a & n253;
  assign n462 = n289 & ~n461;
  assign n463 = n151 & n161;
  assign n464 = ~n462 & n463;
  assign n465 = n38 & ~n39;
  assign n466 = ~n403 & n465;
  assign n467 = ~n464 & ~n466;
  assign n468 = ~n160 & ~n162;
  assign n469 = h & ~n468;
  assign n470 = n107 & n457;
  assign n471 = ~n469 & ~n470;
  assign n472 = ~n143 & n471;
  assign n473 = ~n315 & ~n472;
  assign n474 = n467 & ~n473;
  assign n475 = ~n460 & n474;
  assign n476 = ~n455 & n475;
  assign n477 = n454 & n476;
  assign o2 = ~n430 | ~n477;
  assign n479 = n58 & n397;
  assign n480 = k & ~n144;
  assign n481 = n149 & ~n480;
  assign n482 = ~n146 & ~n481;
  assign n483 = ~n315 & ~n482;
  assign n484 = ~n154 & n483;
  assign n485 = ~n479 & ~n484;
  assign n486 = ~n418 & n485;
  assign n487 = ~n143 & ~n433;
  assign n488 = ~n315 & ~n487;
  assign n489 = ~h & ~i;
  assign n490 = k & ~n318;
  assign n491 = ~n489 & n490;
  assign n492 = ~n403 & n491;
  assign n493 = n454 & ~n492;
  assign n494 = ~n488 & n493;
  assign n495 = j & ~n494;
  assign n496 = ~k & ~l;
  assign n497 = ~h & n50;
  assign n498 = ~j & k;
  assign n499 = i & ~n498;
  assign n500 = n497 & n499;
  assign n501 = ~n496 & n500;
  assign n502 = ~n218 & ~n501;
  assign n503 = ~n295 & ~n502;
  assign n504 = n428 & ~n503;
  assign n505 = ~n495 & n504;
  assign p2 = ~n486 | ~n505;
  assign n507 = ~m & n65;
  assign n508 = ~n396 & n507;
  assign n509 = ~j & n34;
  assign n510 = ~n350 & ~n509;
  assign n511 = ~n175 & n510;
  assign n512 = ~n403 & ~n511;
  assign n513 = ~j & n451;
  assign n514 = ~n512 & ~n513;
  assign n515 = ~n508 & n514;
  assign n516 = n453 & n515;
  assign n517 = l & ~n516;
  assign n518 = k & n407;
  assign n519 = ~n424 & n518;
  assign n520 = n347 & n394;
  assign n521 = ~n510 & n520;
  assign n522 = g & n521;
  assign n523 = n65 & n149;
  assign n524 = n293 & n523;
  assign n525 = ~n522 & ~n524;
  assign n526 = ~n519 & n525;
  assign n527 = l & n307;
  assign n528 = n & n527;
  assign n529 = ~j & ~n386;
  assign n530 = n58 & n362;
  assign n531 = h & n530;
  assign n532 = ~n529 & ~n531;
  assign n533 = n528 & ~n532;
  assign n534 = n401 & n518;
  assign n535 = h & n534;
  assign n536 = n275 & n376;
  assign n537 = n294 & n523;
  assign n538 = ~n536 & ~n537;
  assign n539 = g & n149;
  assign n540 = n54 & n539;
  assign n541 = ~n315 & n540;
  assign n542 = n538 & ~n541;
  assign n543 = ~n535 & n542;
  assign n544 = ~n533 & n543;
  assign n545 = ~n379 & n544;
  assign n546 = n526 & n545;
  assign n547 = ~n54 & ~n61;
  assign n548 = ~n295 & ~n547;
  assign n549 = ~n61 & ~n65;
  assign n550 = n359 & ~n549;
  assign n551 = k & n275;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n288 & n332;
  assign n554 = ~n65 & n74;
  assign n555 = ~n553 & n554;
  assign n556 = n552 & ~n555;
  assign n557 = ~n548 & n556;
  assign n558 = n149 & ~n557;
  assign n559 = n546 & ~n558;
  assign q2 = n517 | ~n559;
  assign n561 = ~g & n90;
  assign n562 = n73 & n561;
  assign n563 = ~n336 & ~n562;
  assign n564 = ~n225 & n335;
  assign n565 = n563 & ~n564;
  assign n566 = e & n188;
  assign n567 = ~n565 & n566;
  assign n568 = n221 & n358;
  assign n569 = ~n162 & n568;
  assign n570 = n294 & ~n569;
  assign n571 = e & n278;
  assign n572 = i & n85;
  assign n573 = n348 & n572;
  assign n574 = n310 & n573;
  assign n575 = n571 & n574;
  assign n576 = n142 & n275;
  assign n577 = n538 & ~n576;
  assign n578 = ~n330 & n577;
  assign n579 = ~n575 & n578;
  assign n580 = ~n570 & n579;
  assign n581 = n29 & n518;
  assign n582 = ~h & n193;
  assign n583 = n571 & n582;
  assign n584 = n581 & n583;
  assign n585 = ~f & n278;
  assign n586 = n74 & n86;
  assign n587 = n446 & n496;
  assign n588 = ~i & n587;
  assign n589 = ~n586 & ~n588;
  assign n590 = n29 & ~n589;
  assign n591 = n585 & n590;
  assign n592 = ~n584 & ~n591;
  assign n593 = n580 & n592;
  assign n594 = ~n567 & n593;
  assign n595 = n70 & n335;
  assign n596 = ~n562 & ~n595;
  assign n597 = n49 & ~n596;
  assign n598 = c & n597;
  assign n599 = n594 & ~n598;
  assign n600 = ~d & ~n195;
  assign n601 = n229 & ~n600;
  assign n602 = ~a & n79;
  assign n603 = ~n601 & n602;
  assign n604 = n189 & ~n241;
  assign n605 = n204 & n264;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n603 & n606;
  assign h2 = ~n599 | ~n607;
  assign n609 = c & n132;
  assign n610 = ~n268 & ~n609;
  assign n611 = n181 & ~n610;
  assign n612 = b & n611;
  assign n613 = ~h & n58;
  assign n614 = n527 & n613;
  assign n615 = ~b & n44;
  assign n616 = g & n;
  assign n617 = n122 & n616;
  assign n618 = n615 & n617;
  assign n619 = n614 & n618;
  assign n620 = ~h & n335;
  assign n621 = n581 & n620;
  assign n622 = n254 & n621;
  assign n623 = ~n619 & ~n622;
  assign n624 = ~f & ~g;
  assign n625 = n34 & n36;
  assign n626 = n29 & n625;
  assign n627 = n624 & n626;
  assign n628 = n388 & n627;
  assign n629 = g & n90;
  assign n630 = n573 & n629;
  assign n631 = n204 & n630;
  assign n632 = n79 & n242;
  assign n633 = n335 & n632;
  assign n634 = n85 & n318;
  assign n635 = n347 & n634;
  assign n636 = n633 & n635;
  assign n637 = ~n631 & ~n636;
  assign n638 = ~n628 & n637;
  assign n639 = n79 & n181;
  assign n640 = n193 & n639;
  assign n641 = ~m & n496;
  assign n642 = n613 & n641;
  assign n643 = n640 & n642;
  assign n644 = n180 & n181;
  assign n645 = g & n644;
  assign n646 = ~h & n645;
  assign n647 = ~l & n29;
  assign n648 = n59 & n647;
  assign n649 = n646 & n648;
  assign n650 = ~n643 & ~n649;
  assign n651 = n638 & n650;
  assign n652 = n623 & n651;
  assign n653 = n171 & ~n565;
  assign n654 = n652 & ~n653;
  assign n655 = ~n612 & n654;
  assign n656 = ~n169 & ~n363;
  assign n657 = ~n109 & ~n656;
  assign n658 = ~n136 & ~n657;
  assign n659 = ~n247 & n658;
  assign n660 = d & ~n659;
  assign n661 = n655 & ~n660;
  assign n662 = n169 & n600;
  assign n663 = ~n201 & ~n207;
  assign n664 = ~n100 & ~n663;
  assign n665 = ~n662 & ~n664;
  assign n666 = a & ~n665;
  assign n667 = ~i & n29;
  assign n668 = n278 & n667;
  assign n669 = ~e & ~f;
  assign n670 = n587 & n669;
  assign n671 = n668 & n670;
  assign n672 = n614 & n633;
  assign n673 = n204 & n621;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n671 & n674;
  assign n676 = n133 & n639;
  assign n677 = n675 & ~n676;
  assign n678 = ~n120 & n580;
  assign n679 = n677 & n678;
  assign n680 = ~n78 & n679;
  assign n681 = ~n666 & n680;
  assign i2 = ~n661 | ~n681;
  assign n683 = n199 & n230;
  assign n684 = n353 & n683;
  assign n685 = n523 & n684;
  assign n686 = n30 & n507;
  assign n687 = l & n618;
  assign n688 = n686 & n687;
  assign n689 = ~n685 & ~n688;
  assign n690 = i & n65;
  assign n691 = n620 & n690;
  assign n692 = n348 & n691;
  assign n693 = n254 & n692;
  assign n694 = n674 & ~n693;
  assign n695 = n689 & n694;
  assign n696 = n618 & n635;
  assign n697 = n634 & n683;
  assign n698 = n539 & n697;
  assign n699 = ~n696 & ~n698;
  assign n700 = n254 & n630;
  assign n701 = ~n584 & ~n700;
  assign n702 = n637 & n701;
  assign n703 = n699 & n702;
  assign n704 = ~l & n85;
  assign n705 = ~f & n668;
  assign n706 = n704 & n705;
  assign n707 = n446 & n706;
  assign n708 = ~n628 & ~n707;
  assign n709 = n703 & n708;
  assign j2 = ~n695 | ~n709;
  assign n711 = f & n48;
  assign n712 = n80 & n711;
  assign n713 = n319 & n431;
  assign n714 = g & n713;
  assign n715 = n712 & n714;
  assign n716 = n319 & n527;
  assign n717 = n640 & n716;
  assign n718 = ~n715 & ~n717;
  assign n719 = n39 & n348;
  assign n720 = i & n645;
  assign n721 = n719 & n720;
  assign n722 = k & n721;
  assign n723 = n623 & ~n722;
  assign n724 = n703 & n723;
  assign n725 = n718 & n724;
  assign n726 = n571 & n627;
  assign n727 = ~n671 & ~n726;
  assign k2 = ~n725 | ~n727;
  assign n729 = n204 & n347;
  assign n730 = ~i & ~k;
  assign n731 = ~j & n730;
  assign n732 = b & n;
  assign n733 = n731 & ~n732;
  assign n734 = n729 & n733;
  assign n735 = n561 & n734;
  assign n736 = n602 & n620;
  assign n737 = n110 & n736;
  assign n738 = n457 & n737;
  assign n739 = ~n735 & ~n738;
  assign n740 = ~n575 & n739;
  assign n741 = n650 & n740;
  assign n742 = ~n591 & n741;
  assign n743 = n695 & n742;
  assign m2 = ~n725 | ~n743;
  assign n745 = ~n & n686;
  assign n746 = ~n626 & ~n745;
  assign n747 = ~d & ~n746;
  assign n748 = n122 & n167;
  assign n749 = n50 & n634;
  assign n750 = ~n748 & n749;
  assign n751 = n81 & n388;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~c & ~m;
  assign n754 = ~n81 & ~n753;
  assign n755 = ~e & n489;
  assign n756 = ~n754 & n755;
  assign n757 = ~n713 & ~n756;
  assign n758 = ~n79 & ~n757;
  assign n759 = ~n705 & ~n758;
  assign n760 = n752 & n759;
  assign n761 = ~n747 & n760;
  assign n762 = g & ~n761;
  assign n763 = c & ~n170;
  assign n764 = ~n180 & ~n763;
  assign n765 = ~b & n764;
  assign n766 = n314 & n489;
  assign n767 = ~n586 & ~n766;
  assign n768 = ~n765 & n767;
  assign n769 = ~m & ~n768;
  assign n770 = ~m & n730;
  assign n771 = ~n58 & n307;
  assign n772 = ~n770 & ~n771;
  assign n773 = n615 & ~n772;
  assign n774 = ~i & n496;
  assign n775 = ~m & ~n318;
  assign n776 = ~n774 & n775;
  assign n777 = ~m & n52;
  assign n778 = ~j & ~m;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~n776 & n779;
  assign n781 = n640 & ~n780;
  assign n782 = ~n773 & ~n781;
  assign n783 = ~n769 & n782;
  assign n784 = n & ~n783;
  assign n785 = g & n489;
  assign n786 = ~c & n785;
  assign n787 = c & n669;
  assign n788 = g & n278;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~n720 & n789;
  assign n791 = ~n786 & n790;
  assign n792 = n647 & ~n791;
  assign n793 = n71 & n626;
  assign n794 = ~b & n624;
  assign n795 = n81 & ~n85;
  assign n796 = ~l & n81;
  assign n797 = ~n795 & ~n796;
  assign n798 = n794 & ~n797;
  assign n799 = ~n793 & ~n798;
  assign n800 = ~n792 & n799;
  assign n801 = ~n48 & n669;
  assign n802 = ~n244 & ~n712;
  assign n803 = ~n801 & n802;
  assign n804 = n138 & ~n803;
  assign n805 = c & n667;
  assign n806 = ~n142 & ~n805;
  assign n807 = n446 & ~n806;
  assign n808 = ~n804 & ~n807;
  assign n809 = ~k & n778;
  assign n810 = ~n155 & ~n353;
  assign n811 = n809 & ~n810;
  assign n812 = n808 & ~n811;
  assign n813 = n800 & n812;
  assign n814 = ~n784 & n813;
  assign n815 = ~n762 & n814;
  assign n816 = ~a & n714;
  assign n817 = ~n278 & ~n634;
  assign n818 = n29 & ~n788;
  assign n819 = ~n817 & n818;
  assign n820 = ~n816 & ~n819;
  assign n821 = n244 & ~n318;
  assign n822 = a & n111;
  assign n823 = ~n279 & ~n822;
  assign n824 = ~n821 & n823;
  assign n825 = n50 & ~n824;
  assign n826 = n131 & n571;
  assign n827 = n142 & n244;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n732 & ~n754;
  assign n830 = n625 & n829;
  assign n831 = f & ~n830;
  assign n832 = n828 & n831;
  assign n833 = ~n825 & n832;
  assign n834 = b & n496;
  assign n835 = n81 & ~n834;
  assign n836 = ~n376 & ~n835;
  assign n837 = n489 & ~n836;
  assign n838 = n833 & ~n837;
  assign n839 = n820 & n838;
  assign n840 = c & ~n746;
  assign n841 = ~a & ~d;
  assign n842 = n376 & ~n841;
  assign n843 = ~n796 & ~n842;
  assign n844 = n489 & ~n843;
  assign n845 = n131 & ~n207;
  assign n846 = ~n130 & n845;
  assign n847 = n686 & n732;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~f & n848;
  assign n850 = ~n844 & n849;
  assign n851 = ~n58 & n795;
  assign n852 = ~n54 & n81;
  assign n853 = ~n151 & n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = n632 & ~n854;
  assign n856 = n850 & ~n855;
  assign n857 = ~n840 & n856;
  assign n858 = ~n839 & ~n857;
  assign n859 = n815 & ~n858;
  assign n860 = ~n65 & ~n803;
  assign n861 = ~g & n860;
  assign n862 = n96 & n634;
  assign n863 = n31 & n489;
  assign n864 = ~b & n129;
  assign n865 = ~n863 & ~n864;
  assign n866 = n44 & ~n865;
  assign n867 = ~n862 & ~n866;
  assign n868 = ~h & n624;
  assign n869 = ~n801 & ~n868;
  assign n870 = j & ~n869;
  assign n871 = n65 & n71;
  assign n872 = n276 & n871;
  assign n873 = ~n870 & ~n872;
  assign n874 = n867 & n873;
  assign n875 = ~n499 & n712;
  assign n876 = f & n446;
  assign n877 = ~a & ~b;
  assign n878 = ~n876 & ~n877;
  assign n879 = m & n878;
  assign n880 = ~n875 & n879;
  assign n881 = ~n704 & n880;
  assign n882 = n874 & n881;
  assign n883 = ~n861 & n882;
  assign n884 = ~n720 & ~n785;
  assign n885 = ~j & ~n884;
  assign n886 = n30 & n871;
  assign n887 = ~n278 & n586;
  assign n888 = ~g & ~n731;
  assign n889 = ~n155 & ~n888;
  assign n890 = n787 & ~n889;
  assign n891 = ~n887 & ~n890;
  assign n892 = ~c & n44;
  assign n893 = ~n787 & ~n892;
  assign n894 = ~n140 & ~n350;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~m & ~n895;
  assign n897 = n891 & n896;
  assign n898 = ~n886 & n897;
  assign n899 = ~n885 & n898;
  assign n900 = ~n883 & ~n899;
  assign n901 = ~c & n624;
  assign n902 = n776 & n901;
  assign n903 = ~n620 & ~n788;
  assign n904 = n770 & ~n903;
  assign n905 = n507 & n720;
  assign n906 = ~n904 & ~n905;
  assign n907 = n191 & n809;
  assign n908 = n193 & n304;
  assign n909 = j & n34;
  assign n910 = ~n181 & n909;
  assign n911 = n908 & n910;
  assign n912 = ~n907 & ~n911;
  assign n913 = ~n585 & ~n901;
  assign n914 = n778 & ~n913;
  assign n915 = i & n914;
  assign n916 = n912 & ~n915;
  assign n917 = ~g & n129;
  assign n918 = n341 & ~n917;
  assign n919 = ~m & n489;
  assign n920 = ~n918 & n919;
  assign n921 = n916 & ~n920;
  assign n922 = n906 & n921;
  assign n923 = ~n892 & ~n901;
  assign n924 = n777 & ~n923;
  assign n925 = n922 & ~n924;
  assign n926 = ~n902 & n925;
  assign n927 = ~n900 & n926;
  assign n928 = ~n & ~n927;
  assign n929 = ~n144 & n496;
  assign n930 = ~i & ~n122;
  assign n931 = ~j & n615;
  assign n932 = ~n794 & ~n871;
  assign n933 = ~n931 & n932;
  assign n934 = ~n930 & n933;
  assign n935 = ~n929 & n934;
  assign n936 = n81 & ~n935;
  assign n937 = n278 & n778;
  assign n938 = ~n496 & ~n937;
  assign n939 = n300 & ~n938;
  assign n940 = n101 & n667;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n936 & n941;
  assign n943 = n145 & n456;
  assign n944 = ~h & ~n943;
  assign n945 = n942 & n944;
  assign n946 = n122 & ~n364;
  assign n947 = n81 & ~n946;
  assign n948 = ~n45 & ~n101;
  assign n949 = n29 & ~n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = n85 & ~n950;
  assign n952 = j & n81;
  assign n953 = n615 & n952;
  assign n954 = n572 & n829;
  assign n955 = ~e & n954;
  assign n956 = ~n953 & ~n955;
  assign n957 = ~n951 & n956;
  assign n958 = n50 & n669;
  assign n959 = ~n48 & n958;
  assign n960 = ~n668 & ~n959;
  assign n961 = n957 & n960;
  assign n962 = h & n961;
  assign n963 = ~n945 & ~n962;
  assign n964 = ~k & n901;
  assign n965 = ~l & ~n923;
  assign n966 = ~n964 & ~n965;
  assign n967 = j & ~n789;
  assign n968 = ~n646 & ~n967;
  assign n969 = n966 & n968;
  assign n970 = n29 & ~n969;
  assign n971 = ~k & n81;
  assign n972 = ~n796 & ~n971;
  assign n973 = n640 & ~n972;
  assign n974 = n39 & n528;
  assign n975 = ~n644 & n974;
  assign n976 = n50 & ~n869;
  assign n977 = ~n & n937;
  assign n978 = k & n977;
  assign n979 = ~n976 & ~n978;
  assign n980 = ~n975 & n979;
  assign n981 = ~n973 & n980;
  assign n982 = ~n970 & n981;
  assign n983 = i & ~n982;
  assign n984 = n443 & n748;
  assign n985 = n414 & ~n984;
  assign n986 = ~g & n985;
  assign n987 = n335 & n713;
  assign n988 = ~n986 & ~n987;
  assign n989 = n161 & n613;
  assign n990 = n988 & ~n989;
  assign n991 = n151 & n971;
  assign n992 = ~n686 & ~n991;
  assign n993 = f & ~n992;
  assign n994 = ~n145 & ~n497;
  assign n995 = n712 & ~n994;
  assign n996 = n318 & n496;
  assign n997 = n778 & n996;
  assign n998 = ~n995 & ~n997;
  assign n999 = ~n993 & n998;
  assign n1000 = ~h & n496;
  assign n1001 = n645 & ~n1000;
  assign n1002 = ~n444 & ~n1001;
  assign n1003 = n667 & ~n1002;
  assign n1004 = ~a & ~c;
  assign n1005 = ~n207 & ~n1004;
  assign n1006 = n958 & ~n1005;
  assign n1007 = ~n1003 & ~n1006;
  assign n1008 = n999 & n1007;
  assign n1009 = n990 & n1008;
  assign n1010 = ~n983 & n1009;
  assign n1011 = ~n963 & n1010;
  assign n1012 = ~n928 & n1011;
  assign l2 = ~n859 | ~n1012;
endmodule


