// Benchmark "top" written by ABC on Sun Apr 24 20:33:48 2016

module top ( clock, 
    tin_pdata_8_8_, tin_pdata_0_0_, tin_pdata_7_7_, preset_0_0_,
    tin_pdata_2_2_, tin_pdata_9_9_, tin_pdata_1_1_, tin_pdata_4_4_, pclk,
    pirq_0_0_, tin_pdata_10_10_, tin_pdata_3_3_, tin_pdata_6_6_,
    tin_pdata_15_15_, tin_pdata_11_11_, tin_pdata_14_14_, tin_pdata_12_12_,
    tin_pdata_5_5_, preset, tin_pdata_13_13_,
    ppeakb_7_7_, ppeakp_12_12_, ppeakp_0_0_, ppeaka_7_7_, ppeaki_15_15_,
    ppeaki_11_11_, ppeaki_3_3_, paddress_3_3_, pdata_8_8_, pdata_0_0_,
    ppeakb_14_14_, ppeakb_10_10_, ppeakb_8_8_, ppeakp_1_1_, ppeaka_14_14_,
    ppeaka_10_10_, ppeaka_8_8_, ppeaki_4_4_, paddress_15_15_,
    paddress_11_11_, paddress_2_2_, ppeakb_9_9_, ppeakp_2_2_, ppeaka_9_9_,
    ppeaks_12_12_, ppeaks_0_0_, ppeaki_5_5_, paddress_5_5_, pdata_7_7_,
    ppeakb_15_15_, ppeakp_3_3_, pwr_0_0_, ppeaks_1_1_, ppeaki_6_6_,
    paddress_4_4_, piack_0_0_, ppeakp_13_13_, ppeakp_4_4_, ppeaka_15_15_,
    ppeaka_11_11_, ppeaks_2_2_, ppeaki_7_7_, paddress_10_10_,
    paddress_7_7_, pdata_2_2_, ppeakp_5_5_, ppeaks_13_13_, ppeaks_3_3_,
    ppeaki_14_14_, ppeaki_10_10_, ppeaki_8_8_, paddress_6_6_, ppeakp_6_6_,
    ppeaks_4_4_, ppeaki_9_9_, paddress_9_9_, pdata_9_9_, pdata_1_1_,
    ppeakb_11_11_, ppeakp_7_7_, ppeaks_5_5_, paddress_13_13_,
    paddress_8_8_, ppeakp_14_14_, ppeakp_10_10_, ppeakp_8_8_, ppeaks_6_6_,
    ppeaki_13_13_, pdata_4_4_, ppeakb_0_0_, ppeakp_9_9_, ppeaka_0_0_,
    ppeaks_7_7_, ppeakb_1_1_, ppeaka_1_1_, ppeaks_10_10_, ppeaks_8_8_,
    pdata_10_10_, pdata_3_3_, ppeakb_12_12_, ppeakb_2_2_, ppeaka_12_12_,
    ppeaka_2_2_, ppeaks_15_15_, ppeaks_9_9_, ppeakb_3_3_, ppeakp_15_15_,
    ppeakp_11_11_, ppeaka_13_13_, ppeaka_3_3_, paddress_14_14_,
    paddress_12_12_, pdata_6_6_, ppeakb_13_13_, ppeakb_4_4_, pdn,
    ppeaka_4_4_, ppeaki_0_0_, prd_0_0_, pdata_15_15_, pdata_11_11_,
    ppeakb_5_5_, ppeaka_5_5_, ppeaks_14_14_, ppeaki_1_1_, paddress_1_1_,
    pdata_14_14_, pdata_12_12_, pdata_5_5_, ppeakb_6_6_, ppeaka_6_6_,
    ppeaks_11_11_, ppeaki_12_12_, ppeaki_2_2_, paddress_0_0_, pdata_13_13_  );
  input  clock;
  input  tin_pdata_8_8_, tin_pdata_0_0_, tin_pdata_7_7_, preset_0_0_,
    tin_pdata_2_2_, tin_pdata_9_9_, tin_pdata_1_1_, tin_pdata_4_4_, pclk,
    pirq_0_0_, tin_pdata_10_10_, tin_pdata_3_3_, tin_pdata_6_6_,
    tin_pdata_15_15_, tin_pdata_11_11_, tin_pdata_14_14_, tin_pdata_12_12_,
    tin_pdata_5_5_, preset, tin_pdata_13_13_;
  output ppeakb_7_7_, ppeakp_12_12_, ppeakp_0_0_, ppeaka_7_7_, ppeaki_15_15_,
    ppeaki_11_11_, ppeaki_3_3_, paddress_3_3_, pdata_8_8_, pdata_0_0_,
    ppeakb_14_14_, ppeakb_10_10_, ppeakb_8_8_, ppeakp_1_1_, ppeaka_14_14_,
    ppeaka_10_10_, ppeaka_8_8_, ppeaki_4_4_, paddress_15_15_,
    paddress_11_11_, paddress_2_2_, ppeakb_9_9_, ppeakp_2_2_, ppeaka_9_9_,
    ppeaks_12_12_, ppeaks_0_0_, ppeaki_5_5_, paddress_5_5_, pdata_7_7_,
    ppeakb_15_15_, ppeakp_3_3_, pwr_0_0_, ppeaks_1_1_, ppeaki_6_6_,
    paddress_4_4_, piack_0_0_, ppeakp_13_13_, ppeakp_4_4_, ppeaka_15_15_,
    ppeaka_11_11_, ppeaks_2_2_, ppeaki_7_7_, paddress_10_10_,
    paddress_7_7_, pdata_2_2_, ppeakp_5_5_, ppeaks_13_13_, ppeaks_3_3_,
    ppeaki_14_14_, ppeaki_10_10_, ppeaki_8_8_, paddress_6_6_, ppeakp_6_6_,
    ppeaks_4_4_, ppeaki_9_9_, paddress_9_9_, pdata_9_9_, pdata_1_1_,
    ppeakb_11_11_, ppeakp_7_7_, ppeaks_5_5_, paddress_13_13_,
    paddress_8_8_, ppeakp_14_14_, ppeakp_10_10_, ppeakp_8_8_, ppeaks_6_6_,
    ppeaki_13_13_, pdata_4_4_, ppeakb_0_0_, ppeakp_9_9_, ppeaka_0_0_,
    ppeaks_7_7_, ppeakb_1_1_, ppeaka_1_1_, ppeaks_10_10_, ppeaks_8_8_,
    pdata_10_10_, pdata_3_3_, ppeakb_12_12_, ppeakb_2_2_, ppeaka_12_12_,
    ppeaka_2_2_, ppeaks_15_15_, ppeaks_9_9_, ppeakb_3_3_, ppeakp_15_15_,
    ppeakp_11_11_, ppeaka_13_13_, ppeaka_3_3_, paddress_14_14_,
    paddress_12_12_, pdata_6_6_, ppeakb_13_13_, ppeakb_4_4_, pdn,
    ppeaka_4_4_, ppeaki_0_0_, prd_0_0_, pdata_15_15_, pdata_11_11_,
    ppeakb_5_5_, ppeaka_5_5_, ppeaks_14_14_, ppeaki_1_1_, paddress_1_1_,
    pdata_14_14_, pdata_12_12_, pdata_5_5_, ppeakb_6_6_, ppeaka_6_6_,
    ppeaks_11_11_, ppeaki_12_12_, ppeaki_2_2_, paddress_0_0_, pdata_13_13_;
  reg ndout, ppeakb_12_12_, ppeakb_1_1_, ppeaka_6_6_, \[4295] , \[4310] ,
    ppeaks_5_5_, ppeakp_10_10_, \[4355] , \[4370] , \[4385] , \[4400] ,
    \[4415] , \[4430] , \[4445] , \[4460] , \[4475] , \[4490] , \[4505] ,
    \[4520] , \[4535] , \[4550] , \[4565] , \[4580] , \[4595] , \[4610] ,
    \[4625] , \[4640] , \[4655] , \[4670] , \[4700] , \[4715] , \[4730] ,
    \[4745] , \[4760] , \[4775] , \[4790] , \[4805] , \[4820] , \[4835] ,
    \[4850] , \[4865] , \[4880] , \[4895] , \[4910] , \[4925] , \[4940] ,
    \[4955] , \[4970] , ppeakb_0_0_, ppeaka_7_7_, \[5015] , \[5030] ,
    ppeaks_4_4_, ppeakp_11_11_, \[5075] , \[5090] , \[5105] , \[5120] ,
    \[5135] , \[5150] , \[5165] , \[5180] , \[5195] , \[5210] , \[5225] ,
    \[5240] , \[5255] , \[5270] , \[5285] , \[5300] , \[5315] , \[5330] ,
    \[5345] , \[5360] , \[5375] , \[5390] , \[5405] , \[5420] , \[5435] ,
    \[5450] , \[5465] , \[5480] , \[5495] , \[5510] , \[5525] , \[5540] ,
    \[5555] , \[5570] , \[5600] , \[5615] , \[5630] , \[5645] , \[5660] ,
    \[5675] , ppeakb_10_10_, ppeaka_8_8_, \[5720] , ppeaks_14_14_,
    ppeaks_7_7_, ppeakp_12_12_, \[5780] , \[5795] , \[5810] , \[5825] ,
    \[5840] , \[5855] , \[5870] , \[5885] , \[5900] , \[5915] , \[5930] ,
    \[5945] , \[5960] , \[5975] , \[5990] , \[6005] , \[6020] , \[6035] ,
    \[6050] , \[6065] , \[6080] , \[6095] , \[6110] , \[6125] , \[6140] ,
    \[6155] , \[6170] , \[6185] , \[6200] , \[6215] , \[6230] , \[6245] ,
    \[6260] , \[6275] , \[6290] , \[6305] , \[6320] , \[6335] , \[6350] ,
    \[6365] , ppeakb_11_11_, ppeakb_2_2_, \[6410] , ppeaks_15_15_,
    ppeaks_6_6_, ppeakp_13_13_, \[6470] , \[6485] , \[6500] , \[6515] ,
    \[6530] , \[6545] , \[6560] , \[6575] , \[6590] , \[6605] , \[6620] ,
    \[6635] , \[6650] , \[6665] , \[6680] , \[6695] , \[6710] , \[6725] ,
    \[6740] , \[6755] , \[6770] , \[6785] , \[6815] , \[6830] , \[6845] ,
    \[6860] , \[6875] , \[6890] , \[6905] , \[6920] , \[6935] , \[6950] ,
    \[6965] , \[6980] , \[6995] , \[7010] , \[7025] , \[7055] ,
    ppeaks_12_12_, ppeaks_1_1_, ppeakp_3_3_, \[7115] , \[7130] , \[7145] ,
    \[7160] , \[7175] , \[7190] , \[7205] , \[7220] , \[7235] , \[7250] ,
    \[7265] , \[7280] , \[7295] , \[7310] , \[7325] , \[7340] , \[7355] ,
    \[7370] , \[7385] , \[7400] , \[7415] , \[7430] , \[7445] , \[7460] ,
    \[7475] , \[7490] , \[7505] , \[7520] , \[7535] , \[7550] , \[7565] ,
    \[7580] , \[7595] , \[7625] , \[7640] , \[7655] , \[7670] , \[7685] ,
    ppeaks_13_13_, ppeakp_7_7_, ppeakp_2_2_, \[7745] , \[7760] , \[7775] ,
    \[7790] , \[7805] , \[7820] , \[7835] , \[7850] , \[7865] , \[7880] ,
    \[7895] , \[7910] , \[7925] , \[7940] , \[7955] , \[7970] , \[8000] ,
    \[8015] , \[8030] , \[8045] , \[8060] , \[8075] , \[8090] , \[8105] ,
    \[8120] , \[8135] , \[8150] , \[8165] , \[8180] , \[8195] , \[8210] ,
    \[8225] , \[8240] , \[8255] , \[8285] , \[8300] , \[8315] , \[8330] ,
    ppeaks_3_3_, ppeakp_8_8_, ppeakp_1_1_, \[8390] , \[8405] , \[8420] ,
    \[8435] , \[8450] , \[8465] , \[8480] , \[8495] , \[8510] , \[8525] ,
    \[8540] , \[8555] , \[8570] , \[8585] , \[8600] , \[8615] , \[8630] ,
    \[8645] , \[8660] , \[8675] , \[8690] , \[8705] , \[8720] , \[8735] ,
    \[8750] , \[8765] , \[8780] , \[8810] , \[8825] , \[8840] , \[8855] ,
    \[8870] , \[8885] , \[8900] , \[8915] , \[8930] , \[8945] , \[8960] ,
    \[8975] , ppeaks_11_11_, ppeaks_2_2_, ppeakp_9_9_, ppeakp_0_0_,
    \[9050] , \[9065] , \[9080] , \[9095] , \[9110] , \[9125] , \[9140] ,
    \[9155] , \[9170] , \[9185] , \[9200] , \[9215] , \[9230] , \[9245] ,
    \[9260] , \[9275] , \[9290] , \[9305] , \[9320] , \[9335] , \[9350] ,
    \[9365] , \[9380] , \[9395] , \[9410] , \[9440] , \[9455] , \[9470] ,
    \[9485] , \[9500] , \[9515] , \[9530] , \[9545] , \[9560] , \[9575] ,
    \[9590] , \[9605] , \[9620] , \[9635] , \[9650] , \[9665] , \[9680] ,
    ppeaki_6_6_, \[9710] , \[9725] , \[9740] , \[9770] , \[9785] ,
    \[9800] , \[9815] , \[9830] , \[9845] , \[9860] , \[9875] , \[9890] ,
    \[9905] , \[9920] , \[9935] , \[9950] , \[9980] , \[9995] , \[10010] ,
    \[10025] , \[10040] , \[10055] , \[10070] , \[10085] , \[10100] ,
    \[10115] , \[10130] , \[10145] , \[10175] , \[10190] , \[10205] ,
    \[10220] , ppeaki_15_15_, ppeaki_4_4_, \[10265] , \[10280] , \[10310] ,
    \[10325] , \[10340] , \[10355] , \[10370] , \[10400] , \[10415] ,
    \[10430] , \[10445] , \[10460] , \[10475] , \[10490] , \[10505] ,
    ppeaki_14_14_, ppeaki_5_5_, \[10550] , \[10565] , \[10580] , \[10595] ,
    \[10610] , \[10625] , \[10655] , \[10670] , \[10685] , \[10700] ,
    \[10715] , \[10730] , \[10745] , \[10760] , \[10775] , \[10790] ,
    \[10805] , \[10820] , \[10850] , \[10865] , \[10880] , \[10895] ,
    \[10925] , \[10940] , \[10955] , \[10970] , \[10985] , \[11015] ,
    \[11030] , \[11045] , \[11060] , \[11075] , \[11090] , \[11120] ,
    \[11135] , \[11150] , \[11165] , \[11180] , \[11195] , \[11210] ,
    \[11225] , \[11240] , \[11255] , \[11270] , \[11285] , \[11300] ,
    \[11315] , \[11330] , \[11345] , \[11375] , \[11390] , \[11405] ,
    \[11420] , \[11435] , \[11450] , \[11465] , \[11480] , \[11495] ,
    \[11510] , \[11525] , \[11540] , \[11555] , \[11570] , \[11585] ,
    \[11600] , \[11615] , \[11630] , \[11645] , \[11660] , \[11675] ,
    \[11690] , \[11705] , \[11720] , \[11735] , \[11750] , \[11765] ,
    \[11780] , \[11795] , \[11810] , ppeaki_9_9_, ppeakb_14_14_, \[11885] ,
    \[11900] , \[11915] , \[11930] , ppeaki_8_8_, ppeakb_15_15_, \[12005] ,
    \[12020] , \[12035] , \[12050] , \[12065] , \[12080] , ppeaki_7_7_,
    \[12125] , \[12140] , \[12155] , \[12170] , \[12185] , \[12200] ,
    ppeakb_13_13_, \[12245] , \[12260] , \[12275] , ppeaki_13_13_,
    ppeaki_2_2_, \[12335] , \[12350] , \[12365] , \[12380] , \[12395] ,
    \[12410] , \[12425] , \[12440] , \[12455] , \[12470] , \[12485] ,
    ppeaki_12_12_, ppeaki_3_3_, \[12545] , \[12560] , \[12575] , \[12590] ,
    \[12605] , \[12620] , \[12635] , \[12650] , \[12665] , \[12680] ,
    \[12695] , ppeaki_11_11_, ppeaki_0_0_, \[12770] , \[12800] , \[12815] ,
    \[12830] , \[12845] , \[12860] , \[12875] , \[12890] , \[12905] ,
    \[12920] , \[12935] , ppeaki_10_10_, ppeaki_1_1_, \[13010] , \[13025] ,
    \[13040] , \[13055] , \[13070] , \[13085] , \[13100] , \[13115] ,
    \[13130] , \[13160] , \[13175] , ppeakb_4_4_, ppeaka_9_9_, \[13220] ,
    \[13235] , \[13250] , \[13265] , \[13280] , \[13295] , \[13310] ,
    \[13325] , \[13340] , \[13355] , \[13370] , \[13385] , \[13400] ,
    \[13415] , \[13430] , \[13445] , \[13460] , \[13475] , \[13490] ,
    \[13505] , ppeakb_5_5_, \[13550] , ppeakp_6_6_, \[13580] , \[13595] ,
    \[13610] , \[13625] , \[13640] , \[13655] , \[13670] , \[13685] ,
    \[13700] , \[13715] , \[13730] , \[13745] , \[13775] , \[13790] ,
    \[13805] , \[13820] , \[13835] , \[13850] , \[13865] , \[13880] ,
    \[13895] , ppeaka_11_11_, ppeaka_0_0_, ppeakp_5_5_, \[13955] ,
    \[13970] , \[13985] , \[14000] , \[14015] , \[14030] , \[14045] ,
    \[14060] , \[14075] , \[14090] , \[14105] , \[14120] , \[14135] ,
    \[14150] , \[14165] , \[14180] , \[14210] , \[14225] , \[14240] ,
    \[14255] , \[14270] , \[14285] , ppeakb_3_3_, ppeaka_10_10_,
    ppeaka_1_1_, ppeakp_4_4_, \[14360] , \[14375] , \[14390] , \[14405] ,
    \[14420] , \[14435] , \[14450] , \[14465] , \[14480] , \[14495] ,
    \[14510] , \[14525] , \[14540] , \[14555] , \[14570] , \[14585] ,
    \[14600] , \[14615] , \[14630] , \[14660] , \[14675] , \[14690] ,
    \[14705] , ppeakb_8_8_, ppeaka_13_13_, ppeaka_2_2_, \[14765] ,
    ppeaks_9_9_, ppeakp_14_14_, \[14810] , \[14825] , \[14840] , \[14855] ,
    \[14870] , \[14885] , \[14900] , \[14915] , \[14930] , \[14960] ,
    \[14975] , \[14990] , \[15005] , \[15020] , \[15035] , \[15050] ,
    \[15065] , \[15080] , ppeakb_9_9_, ppeaka_12_12_, ppeaka_3_3_,
    \[15140] , ppeaks_8_8_, ppeakp_15_15_, \[15185] , \[15200] , \[15215] ,
    \[15230] , \[15245] , \[15260] , \[15275] , \[15290] , \[15305] ,
    \[15320] , \[15335] , \[15350] , \[15365] , \[15380] , \[15395] ,
    \[15410] , \[15425] , \[15440] , ppeakb_6_6_, ppeaka_15_15_,
    ppeaka_4_4_, \[15500] , \[15515] , ppeaks_0_0_, \[15545] , \[15560] ,
    \[15575] , \[15590] , \[15605] , \[15620] , \[15635] , \[15650] ,
    \[15665] , \[15680] , \[15695] , \[15710] , \[15725] , \[15755] ,
    \[15770] , \[15785] , ppeakb_7_7_, ppeaka_14_14_, ppeaka_5_5_,
    \[15845] , \[15860] , ppeaks_10_10_, \[15890] , \[15905] , \[15920] ,
    \[15935] , \[15950] , \[15965] , \[15980] , \[15995] , \[16010] ,
    \[16025] , \[16040] , \[16055] , \[16070] , \[16085] , \[16100] ,
    paddress_8_8_, \[16907] , \[16920] , \[16933] , paddress_9_9_,
    \[16959] , \[16972] , \[16985] , \[16998] , \[17011] , \[17024] ,
    \[17037] , \[17050] , \[17063] , \[17076] , \[17089] , \[17102] ,
    \[17115] , \[17128] , \[17141] , \[17154] , \[17167] , \[17180] ,
    \[17193] , \[17206] , \[17219] , \[17232] , \[17245] , \[17258] ,
    \[17271] , \[17284] , \[17297] , \[17310] , \[17323] , \[17336] ,
    \[17349] , \[17362] , \[17375] , \[17388] , paddress_11_11_, \[17414] ,
    \[17427] , \[17453] , paddress_10_10_, \[17479] , \[17492] , \[17505] ,
    \[17518] , \[17531] , \[17544] , paddress_13_13_, \[17570] , \[17583] ,
    \[17596] , \[17609] , paddress_12_12_, \[17635] , \[17648] , \[17661] ,
    \[17674] , paddress_15_15_, \[17700] , \[17713] , paddress_14_14_,
    \[17739] , \[17752] , \[17765] , \[17778] , \[17791] , \[17804] ,
    \[17817] , pwr_0_0_, \[17843] , \[17856] , \[17869] , \[17882] ,
    prd_0_0_, \[17908] , \[17921] , \[17934] , \[17947] , \[17960] ,
    \[17973] , \[17986] , \[17999] , \[18012] , \[18025] , \[18038] , pdn,
    \[18064] , \[18077] , \[18090] , \[18103] , \[18116] , \[18129] ,
    \[18142] , \[18155] , \[18168] , \[18181] , \[18194] , \[18207] ,
    \[18220] , \[18233] , \[18246] , paddress_0_0_, piack_0_0_, \[18285] ,
    \[18298] , \[18311] , paddress_1_1_, \[18337] , \[18350] , \[18363] ,
    \[18376] , \[18389] , paddress_2_2_, \[18415] , \[18428] , \[18441] ,
    paddress_3_3_, \[18467] , \[18480] , \[18493] , \[18506] ,
    paddress_4_4_, paddress_5_5_, \[18545] , paddress_6_6_, \[18571] ,
    \[18584] , \[18597] , \[18610] , paddress_7_7_, \[18636] ;
  wire n2795, n2796, n2798, n2799_1, n2801, n2802, n2804_1, n2805, n2807,
    n2808, n2810, n2811, n2813, n2814_1, n2816, n2817, n2819_1, n2820,
    n2822, n2823, n2825, n2826, n2828, n2829_1, n2831, n2832, n2834_1,
    n2835, n2837, n2838, n2840, n2841, n2843, n2844_1, n2845, n2846, n2848,
    n2849_1, n2850, n2851, n2852, n2853_1, n2854, n2855, n2856, n2857_1,
    n2858, n2859, n2860, n2861, n2862_1, n2863, n2864, n2865, n2866,
    n2867_1, n2868, n2869, n2870, n2871, n2872_1, n2873, n2874, n2875,
    n2876, n2877_1, n2878, n2879, n2880, n2881, n2882_1, n2883, n2884,
    n2885, n2886, n2887_1, n2888, n2889, n2890, n2891, n2892_1, n2893,
    n2894, n2895, n2896, n2897_1, n2898, n2899, n2900, n2901, n2902_1,
    n2903, n2904, n2905, n2906, n2907_1, n2908, n2909, n2910, n2911,
    n2912_1, n2913, n2914, n2915, n2916_1, n2917, n2918, n2919, n2920_1,
    n2921, n2922, n2923, n2924, n2925_1, n2926, n2927, n2928, n2929,
    n2930_1, n2931, n2932, n2933, n2934, n2935_1, n2936, n2937, n2938,
    n2939, n2940_1, n2941, n2942, n2943, n2944, n2945_1, n2946, n2947,
    n2948, n2949, n2950_1, n2951, n2952, n2953, n2954, n2955_1, n2956,
    n2957, n2958, n2959, n2960_1, n2961, n2962, n2963, n2964, n2965_1,
    n2966, n2967, n2968, n2969, n2970_1, n2971, n2972, n2973, n2974,
    n2975_1, n2976, n2977, n2978, n2979_1, n2980, n2981, n2982, n2983_1,
    n2984, n2985, n2986, n2987, n2988_1, n2989, n2990, n2991, n2993_1,
    n2994, n2995, n2996, n2997, n2998_1, n2999, n3000, n3001, n3002,
    n3003_1, n3004, n3005, n3006, n3007, n3008_1, n3009, n3010, n3011,
    n3012, n3013_1, n3014, n3015, n3016, n3018_1, n3019, n3020, n3021,
    n3022, n3023_1, n3024, n3025, n3026, n3027, n3028_1, n3029, n3030,
    n3031, n3032, n3033_1, n3034, n3035, n3036, n3037, n3038_1, n3039,
    n3040, n3041, n3042_1, n3043, n3044, n3045, n3046_1, n3047, n3048,
    n3049, n3050, n3051_1, n3052, n3053, n3054, n3055, n3056_1, n3057,
    n3058, n3059, n3061_1, n3062, n3063, n3064, n3065, n3066_1, n3067,
    n3068, n3069, n3070, n3071_1, n3072, n3074, n3075, n3076_1, n3077,
    n3078, n3079, n3081_1, n3082, n3083, n3084, n3085, n3086_1, n3087,
    n3088, n3089, n3090, n3091_1, n3092, n3093, n3094, n3095, n3096_1,
    n3097, n3098, n3099, n3100, n3101_1, n3102, n3103, n3104, n3105,
    n3106_1, n3107, n3108, n3109, n3110, n3111_1, n3112, n3113, n3114,
    n3115, n3116_1, n3117, n3118, n3119, n3120, n3121_1, n3122, n3124,
    n3125, n3126_1, n3127, n3128, n3129, n3130, n3131_1, n3132, n3133,
    n3134, n3135, n3136_1, n3137, n3138, n3139, n3140, n3141_1, n3142,
    n3143, n3144, n3145, n3146_1, n3147, n3148, n3149, n3150_1, n3151,
    n3152, n3153, n3154, n3155_1, n3156, n3157, n3158, n3159_1, n3160,
    n3162, n3163, n3164_1, n3165, n3167, n3168, n3169_1, n3171, n3172,
    n3173, n3174_1, n3175, n3176, n3177, n3178, n3179_1, n3181, n3182,
    n3183, n3184_1, n3186, n3187, n3188, n3190, n3191, n3192, n3193,
    n3194_1, n3195, n3197, n3198, n3200, n3201, n3203, n3204_1, n3205,
    n3206, n3208, n3209_1, n3210, n3211, n3213, n3214_1, n3215, n3217,
    n3218, n3219_1, n3220, n3221, n3223, n3224_1, n3225, n3226, n3228,
    n3230, n3231, n3232, n3233, n3234_1, n3236, n3237, n3238, n3239_1,
    n3240, n3241, n3243, n3244_1, n3246, n3247, n3249_1, n3250, n3251,
    n3252, n3254_1, n3255, n3256, n3257, n3259_1, n3260, n3261, n3262,
    n3263, n3264_1, n3265, n3266, n3267, n3268_1, n3269, n3270, n3271,
    n3272_1, n3273, n3274, n3275, n3276_1, n3277, n3278, n3279, n3280,
    n3281_1, n3282, n3283, n3284, n3285, n3286_1, n3287, n3288, n3289,
    n3290, n3291_1, n3292, n3293, n3294, n3295, n3296_1, n3297, n3298,
    n3299, n3300, n3301_1, n3302, n3303, n3304, n3305, n3306_1, n3307,
    n3308, n3309, n3310, n3311_1, n3312, n3313, n3315, n3316_1, n3317,
    n3318, n3319, n3320, n3321_1, n3322, n3323, n3324, n3325, n3326_1,
    n3327, n3328, n3329, n3330, n3331_1, n3332, n3333, n3334, n3335,
    n3336_1, n3337, n3338, n3339, n3340, n3341_1, n3342, n3343, n3344,
    n3345, n3346_1, n3347, n3348, n3349, n3350, n3351_1, n3352, n3353,
    n3354, n3355, n3356_1, n3357, n3358, n3359, n3360, n3361_1, n3362,
    n3363, n3364, n3365, n3366_1, n3367, n3368, n3369, n3370, n3371_1,
    n3372, n3373, n3374, n3375, n3376_1, n3377, n3378, n3379, n3380,
    n3381_1, n3382, n3383, n3384, n3385, n3386_1, n3387, n3388, n3389,
    n3390_1, n3391, n3392, n3393, n3394_1, n3395, n3396, n3397, n3398_1,
    n3399, n3400, n3401, n3402_1, n3403, n3404, n3405, n3406, n3407_1,
    n3408, n3409, n3410, n3411, n3412_1, n3413, n3414, n3415, n3416,
    n3417_1, n3418, n3419, n3420, n3421, n3422_1, n3423, n3424, n3425,
    n3426, n3427_1, n3428, n3429, n3430, n3431, n3432_1, n3433, n3434,
    n3435, n3436, n3437_1, n3438, n3439, n3440, n3441, n3442_1, n3443,
    n3444, n3445, n3446, n3447_1, n3448, n3449, n3450, n3451, n3452_1,
    n3453, n3454, n3455, n3456, n3457_1, n3458, n3459, n3460, n3461,
    n3462_1, n3463, n3464, n3465, n3466, n3467_1, n3468, n3469, n3470,
    n3471, n3472_1, n3473, n3474, n3475, n3476, n3477_1, n3478, n3479,
    n3480, n3481, n3482_1, n3483, n3484, n3485, n3486, n3487_1, n3488,
    n3489, n3490, n3491, n3492_1, n3493, n3494, n3495, n3496, n3497_1,
    n3498, n3499, n3500, n3501, n3502_1, n3503, n3504, n3505, n3506,
    n3507_1, n3508, n3509, n3510, n3511, n3512_1, n3513, n3514, n3515,
    n3516, n3517_1, n3518, n3519, n3520, n3521_1, n3522, n3523, n3524,
    n3525_1, n3526, n3527, n3528, n3529_1, n3530, n3531, n3532, n3533,
    n3534_1, n3535, n3536, n3537, n3538_1, n3539, n3540, n3541, n3542_1,
    n3543, n3545, n3546, n3547_1, n3548, n3549, n3550, n3551, n3553, n3554,
    n3555, n3556, n3557_1, n3558, n3560, n3561, n3562_1, n3563, n3564,
    n3565, n3566, n3568, n3569, n3570, n3571, n3572_1, n3573, n3574, n3575,
    n3577_1, n3578, n3579, n3580, n3581, n3582_1, n3583, n3584, n3585,
    n3586, n3587_1, n3588, n3589, n3590, n3591, n3592_1, n3593, n3594,
    n3595, n3596, n3597_1, n3598, n3599, n3600, n3601, n3602_1, n3603,
    n3604, n3605, n3606, n3607_1, n3608, n3609, n3610, n3611, n3612_1,
    n3613, n3614, n3615, n3616, n3617_1, n3618, n3619, n3620, n3621,
    n3622_1, n3623, n3624, n3625, n3626, n3627_1, n3628, n3629, n3630,
    n3631, n3632_1, n3633, n3634, n3635, n3636_1, n3637, n3638, n3639,
    n3640_1, n3641, n3642, n3643, n3644_1, n3645, n3646, n3647, n3649_1,
    n3650, n3651, n3652, n3653_1, n3654, n3655, n3657_1, n3658, n3659,
    n3660, n3661, n3662_1, n3664, n3665, n3666, n3667_1, n3668, n3669,
    n3671, n3672_1, n3673, n3674, n3675, n3676, n3677_1, n3678, n3680,
    n3681, n3682_1, n3683, n3685, n3686, n3688, n3689, n3690, n3691,
    n3692_1, n3693, n3694, n3695, n3696, n3697_1, n3698, n3699, n3700,
    n3701, n3702_1, n3703, n3704, n3705, n3706, n3707_1, n3708, n3709,
    n3710, n3711, n3712_1, n3713, n3714, n3715, n3716, n3717_1, n3718,
    n3719, n3720, n3721, n3722_1, n3723, n3724, n3725, n3726, n3727_1,
    n3728, n3729, n3730, n3731, n3732_1, n3733, n3734, n3735, n3736,
    n3737_1, n3738, n3739, n3740, n3741, n3742_1, n3743, n3744, n3745,
    n3746, n3747_1, n3748, n3749, n3750, n3751_1, n3752, n3753, n3754,
    n3755_1, n3756, n3757, n3758, n3759_1, n3760, n3761, n3762, n3763,
    n3764_1, n3765, n3766, n3767, n3768, n3769_1, n3770, n3771, n3772,
    n3773_1, n3774, n3775, n3776, n3777, n3778_1, n3779, n3780, n3781,
    n3782, n3783_1, n3784, n3785, n3786, n3787, n3788_1, n3789, n3790,
    n3791, n3792, n3793_1, n3794, n3795, n3796, n3797, n3798_1, n3799,
    n3800, n3801, n3802, n3803_1, n3804, n3805, n3806, n3807, n3808_1,
    n3809, n3810, n3811, n3812, n3813_1, n3814, n3815, n3816, n3817,
    n3818_1, n3819, n3820, n3821, n3822, n3823_1, n3824, n3825, n3826,
    n3827, n3828_1, n3829, n3830, n3831, n3832, n3833_1, n3834, n3835,
    n3836, n3837, n3838_1, n3839, n3840, n3841, n3842, n3843_1, n3844,
    n3845, n3846, n3847, n3848_1, n3849, n3850, n3851, n3852, n3853_1,
    n3854, n3855, n3856, n3857_1, n3858, n3859, n3860, n3861_1, n3862,
    n3863, n3864, n3865_1, n3866, n3867, n3868, n3870_1, n3871, n3872,
    n3873, n3874, n3875_1, n3876, n3877, n3878, n3879_1, n3880, n3881,
    n3882, n3883, n3884_1, n3885, n3886, n3887, n3888, n3889_1, n3890,
    n3891, n3892, n3893, n3894_1, n3895, n3896, n3897, n3898, n3899_1,
    n3900, n3901, n3902, n3903, n3904_1, n3905, n3906, n3907, n3908,
    n3909_1, n3910, n3911, n3912, n3913, n3914_1, n3915, n3916, n3917,
    n3918, n3919_1, n3920, n3921, n3922, n3923, n3924_1, n3925, n3926,
    n3927, n3928, n3929_1, n3930, n3931, n3932, n3933, n3934_1, n3935,
    n3936, n3937, n3938, n3939_1, n3940, n3941, n3942, n3943, n3944_1,
    n3945, n3946, n3947, n3948, n3949_1, n3950, n3951, n3952, n3953,
    n3954_1, n3955, n3956, n3957, n3958_1, n3959, n3960, n3962, n3963_1,
    n3964, n3965, n3966, n3967, n3968_1, n3969, n3971, n3972, n3973_1,
    n3974, n3975, n3976, n3977_1, n3978, n3979, n3980, n3981, n3982_1,
    n3983, n3984, n3985, n3986, n3987_1, n3988, n3989, n3990, n3991,
    n3992_1, n3993, n3994, n3995, n3996, n3997_1, n3998, n3999, n4000,
    n4001, n4002_1, n4003, n4004, n4005, n4006, n4007_1, n4008, n4009,
    n4010, n4011, n4012_1, n4013, n4014, n4015, n4016, n4017_1, n4018,
    n4019, n4020, n4021, n4022_1, n4023, n4024, n4025, n4026, n4027_1,
    n4028, n4029, n4030, n4031, n4032_1, n4033, n4034, n4035, n4036,
    n4037_1, n4038, n4039, n4040, n4041, n4042_1, n4043, n4044, n4045,
    n4046, n4047_1, n4048, n4049, n4050, n4051, n4052_1, n4053, n4054,
    n4055, n4056, n4057_1, n4058, n4059, n4060, n4061, n4062_1, n4063,
    n4064, n4065, n4066, n4067_1, n4068, n4069, n4070, n4071, n4072_1,
    n4073, n4074, n4075, n4076, n4077_1, n4078, n4079, n4080, n4081, n4083,
    n4084, n4085, n4086, n4087_1, n4088, n4089, n4091, n4092_1, n4093,
    n4094, n4095, n4096, n4097_1, n4098, n4100, n4101, n4102_1, n4103,
    n4104, n4105, n4107_1, n4108, n4109, n4110, n4111, n4112_1, n4114,
    n4115, n4116, n4117_1, n4119, n4120, n4121, n4123, n4124, n4125, n4126,
    n4127_1, n4128, n4129, n4130, n4131, n4132_1, n4133, n4134, n4135,
    n4136, n4137_1, n4138, n4139, n4140, n4141, n4142_1, n4143, n4144,
    n4145, n4146, n4147_1, n4149, n4150, n4151_1, n4152, n4153, n4154,
    n4155, n4156_1, n4157, n4158, n4159, n4160, n4161_1, n4162, n4163,
    n4164, n4165, n4166_1, n4167, n4168, n4169, n4170_1, n4171, n4172,
    n4173, n4174, n4175_1, n4177, n4178, n4179, n4180_1, n4181, n4182,
    n4184, n4185_1, n4186, n4187, n4188, n4189, n4191, n4192, n4193, n4194,
    n4195_1, n4196, n4197, n4198, n4199, n4200_1, n4201, n4202, n4203,
    n4204_1, n4205, n4206, n4207, n4208, n4209_1, n4210, n4211, n4212,
    n4213, n4214_1, n4215, n4216, n4217, n4218, n4219_1, n4220, n4221,
    n4222, n4224_1, n4225, n4226, n4227, n4228_1, n4229, n4230, n4231,
    n4232, n4233_1, n4235, n4236, n4237, n4239, n4240, n4241, n4243_1,
    n4244, n4245, n4247, n4248_1, n4249, n4251, n4252_1, n4254, n4255,
    n4257_1, n4258, n4260, n4261, n4262_1, n4264, n4265, n4266_1, n4268,
    n4269, n4270, n4272, n4273, n4274, n4276_1, n4277, n4279, n4280,
    n4281_1, n4283, n4284, n4286_1, n4287, n4289, n4290, n4292, n4293,
    n4294, n4296_1, n4297, n4298, n4299, n4301_1, n4302, n4304, n4305_1,
    n4306, n4308, n4309, n4311, n4312, n4313, n4315_1, n4316, n4317, n4319,
    n4320_1, n4322, n4323, n4324, n4325_1, n4326, n4327, n4329_1, n4330,
    n4331, n4333, n4334_1, n4335, n4337, n4338, n4340, n4341, n4342, n4343,
    n4344_1, n4345, n4347, n4348, n4350, n4351, n4353, n4354_1, n4355,
    n4356, n4357, n4358, n4359_1, n4361, n4362, n4363, n4364_1, n4365,
    n4366, n4367, n4369_1, n4370, n4372, n4373, n4374_1, n4375, n4376,
    n4377, n4378, n4380, n4381, n4384_1, n4385, n4386, n4388_1, n4389,
    n4390, n4391, n4392, n4393_1, n4395, n4396, n4397, n4398_1, n4399,
    n4400, n4402, n4403_1, n4404, n4406, n4407, n4408_1, n4409, n4410,
    n4411, n4412, n4413_1, n4414, n4415, n4416, n4417, n4418_1, n4419,
    n4420, n4421, n4422, n4423_1, n4424, n4425, n4426, n4427, n4428_1,
    n4429, n4431, n4432, n4433_1, n4434, n4435, n4436, n4437, n4438_1,
    n4439, n4440, n4441, n4442, n4443_1, n4444, n4445, n4446, n4447,
    n4448_1, n4449, n4450, n4451, n4452, n4453_1, n4454, n4455, n4456,
    n4457, n4458_1, n4459, n4461, n4462, n4463_1, n4464, n4465, n4466,
    n4468, n4469, n4470, n4471_1, n4472, n4473, n4474, n4475, n4476_1,
    n4477, n4478, n4479, n4480, n4481_1, n4482, n4483, n4484, n4485,
    n4486_1, n4487, n4488, n4489, n4490_1, n4491, n4492, n4493, n4494,
    n4495_1, n4496, n4497, n4498, n4499, n4501, n4502, n4503, n4504,
    n4505_1, n4506, n4507, n4508, n4509, n4510_1, n4511, n4512, n4513,
    n4514, n4515_1, n4516, n4517, n4518, n4519_1, n4520, n4521, n4522,
    n4523, n4524_1, n4525, n4526, n4527, n4528, n4529_1, n4530, n4531,
    n4533, n4534_1, n4535, n4536, n4537, n4538_1, n4539, n4540, n4541,
    n4542, n4544, n4545, n4546, n4548_1, n4549, n4550, n4552, n4553_1,
    n4554, n4556, n4557, n4559, n4560, n4562_1, n4563, n4565, n4566_1,
    n4567, n4569, n4570, n4571_1, n4573, n4574, n4575_1, n4577, n4578,
    n4579, n4581, n4582, n4583, n4585_1, n4586, n4587, n4589, n4590_1,
    n4592, n4593, n4595_1, n4596, n4598, n4599_1, n4600, n4602, n4603,
    n4604, n4605, n4606, n4607, n4609, n4610, n4612, n4613, n4614, n4616,
    n4617, n4619, n4620, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4630, n4631, n4633, n4634, n4635, n4637, n4638, n4639, n4641, n4642,
    n4643, n4645, n4646, n4648, n4649, n4651, n4652, n4654, n4655, n4657,
    n4658, n4659, n4661, n4662, n4663, n4665, n4666, n4667, n4669, n4670,
    n4671, n4672, n4673, n4674, n4676, n4677, n4678, n4680, n4681, n4683,
    n4684, n4685, n4686, n4688, n4689, n4690, n4691, n4692, n4693, n4695,
    n4696, n4698, n4699, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4751, n4752, n4753, n4754, n4755, n4756, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4834, n4835, n4836, n4838, n4839, n4840, n4842, n4843, n4844, n4846,
    n4847, n4849, n4850, n4852, n4853, n4855, n4856, n4857, n4859, n4860,
    n4861, n4863, n4864, n4865, n4867, n4868, n4869, n4871, n4872, n4873,
    n4875, n4876, n4878, n4879, n4881, n4882, n4884, n4885, n4886, n4888,
    n4889, n4891, n4892, n4894, n4895, n4896, n4898, n4899, n4901, n4902,
    n4904, n4905, n4906, n4908, n4909, n4911, n4912, n4913, n4915, n4916,
    n4917, n4919, n4920, n4922, n4923, n4925, n4926, n4928, n4929, n4931,
    n4932, n4933, n4935, n4936, n4937, n4939, n4940, n4941, n4943, n4944,
    n4945, n4947, n4948, n4949, n4951, n4952, n4953, n4954, n4955, n4956,
    n4958, n4959, n4961, n4962, n4964, n4965, n4967, n4968, n4969, n4970,
    n4971, n4972, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
    n5033, n5034, n5035, n5036, n5037, n5038, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5051, n5052, n5053, n5055,
    n5056, n5057, n5059, n5061, n5062, n5064, n5065, n5066, n5068, n5069,
    n5070, n5072, n5073, n5074, n5076, n5077, n5078, n5080, n5081, n5082,
    n5084, n5085, n5086, n5088, n5090, n5092, n5094, n5095, n5096, n5098,
    n5099, n5100, n5102, n5103, n5105, n5106, n5107, n5109, n5110, n5112,
    n5113, n5114, n5116, n5117, n5118, n5120, n5121, n5123, n5124, n5126,
    n5127, n5128, n5130, n5131, n5132, n5134, n5135, n5137, n5138, n5140,
    n5141, n5143, n5144, n5146, n5147, n5148, n5150, n5151, n5152, n5154,
    n5155, n5156, n5158, n5159, n5160, n5162, n5163, n5165, n5166, n5168,
    n5169, n5171, n5172, n5174, n5175, n5177, n5178, n5179, n5180, n5181,
    n5182, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5239, n5240, n5241, n5243, n5244, n5245, n5247,
    n5249, n5250, n5252, n5253, n5254, n5256, n5257, n5258, n5260, n5261,
    n5262, n5264, n5265, n5266, n5268, n5269, n5270, n5272, n5273, n5274,
    n5276, n5278, n5280, n5282, n5283, n5284, n5286, n5287, n5288, n5290,
    n5291, n5293, n5294, n5296, n5297, n5298, n5300, n5301, n5302, n5304,
    n5305, n5307, n5308, n5310, n5311, n5312, n5314, n5315, n5316, n5318,
    n5319, n5321, n5322, n5324, n5325, n5327, n5328, n5330, n5331, n5332,
    n5334, n5335, n5336, n5338, n5339, n5340, n5342, n5343, n5344, n5346,
    n5347, n5349, n5350, n5352, n5353, n5355, n5356, n5358, n5359, n5361,
    n5362, n5364, n5365, n5366, n5367, n5368, n5369, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5426,
    n5427, n5428, n5430, n5431, n5432, n5434, n5436, n5438, n5439, n5441,
    n5442, n5443, n5445, n5446, n5447, n5449, n5450, n5451, n5453, n5454,
    n5455, n5457, n5459, n5461, n5462, n5464, n5465, n5467, n5468, n5469,
    n5471, n5472, n5473, n5475, n5476, n5478, n5479, n5481, n5482, n5484,
    n5485, n5486, n5488, n5489, n5490, n5492, n5493, n5495, n5496, n5498,
    n5499, n5500, n5502, n5503, n5504, n5506, n5507, n5509, n5510, n5512,
    n5513, n5515, n5516, n5518, n5519, n5520, n5522, n5523, n5524, n5526,
    n5527, n5528, n5530, n5531, n5533, n5534, n5536, n5537, n5538, n5540,
    n5541, n5543, n5544, n5546, n5547, n5549, n5550, n5552, n5553, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
    n5639, n5640, n5641, n5643, n5644, n5645, n5647, n5648, n5649, n5651,
    n5653, n5655, n5656, n5657, n5659, n5660, n5661, n5663, n5664, n5665,
    n5667, n5668, n5669, n5671, n5672, n5673, n5675, n5677, n5679, n5680,
    n5682, n5683, n5685, n5686, n5687, n5689, n5690, n5691, n5693, n5694,
    n5696, n5697, n5699, n5700, n5702, n5703, n5704, n5706, n5707, n5708,
    n5710, n5711, n5713, n5714, n5716, n5717, n5718, n5720, n5721, n5722,
    n5724, n5725, n5727, n5728, n5730, n5731, n5733, n5734, n5736, n5737,
    n5738, n5740, n5741, n5742, n5744, n5745, n5746, n5748, n5749, n5750,
    n5752, n5753, n5755, n5756, n5758, n5759, n5760, n5762, n5763, n5765,
    n5766, n5768, n5769, n5771, n5772, n5774, n5775, n5777, n5778, n5779,
    n5780, n5782, n5783, n5784, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5795, n5797, n5798, n5800, n5801, n5803, n5804, n5806,
    n5807, n5809, n5810, n5811, n5813, n5814, n5815, n5817, n5818, n5820,
    n5821, n5823, n5824, n5826, n5827, n5829, n5830, n5832, n5833, n5835,
    n5836, n5838, n5839, n5840, n5842, n5843, n5844, n5845, n5847, n5849,
    n5850, n5852, n5853, n5855, n5856, n5858, n5859, n5861, n5862, n5864,
    n5865, n5866, n5868, n5869, n5870, n5872, n5873, n5875, n5876, n5878,
    n5879, n5881, n5882, n5884, n5885, n5887, n5888, n5890, n5891, n5892,
    n5894, n5895, n5896, n5898, n5899, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5909, n5911, n5912, n5913, n5915, n5916, n5918, n5919,
    n5921, n5922, n5924, n5925, n5926, n5928, n5929, n5930, n5932, n5933,
    n5935, n5936, n5938, n5939, n5941, n5942, n5944, n5945, n5947, n5948,
    n5949, n5951, n5952, n5953, n5955, n5956, n5957, n5959, n5960, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5971, n5972, n5973,
    n5975, n5976, n5977, n5979, n5980, n5981, n5983, n5984, n5986, n5987,
    n5989, n5990, n5992, n5993, n5994, n5996, n5997, n5999, n6000, n6002,
    n6003, n6005, n6006, n6008, n6009, n6011, n6012, n6014, n6015, n6016,
    n6018, n6019, n6020, n6022, n6023, n6024, n6026, n6027, n6028, n6029,
    n6031, n6032, n6033, n6035, n6036, n6037, n6039, n6040, n6042, n6043,
    n6044, n6046, n6047, n6049, n6050, n6051, n6053, n6054, n6055, n6057,
    n6058, n6059, n6061, n6062, n6064, n6065, n6067, n6068, n6070, n6071,
    n6072, n6074, n6075, n6076, n6078, n6079, n6080, n6082, n6083, n6084,
    n6086, n6087, n6088, n6090, n6091, n6093, n6094, n6096, n6097, n6098,
    n6100, n6101, n6103, n6104, n6106, n6107, n6108, n6110, n6111, n6112,
    n6114, n6115, n6117, n6118, n6120, n6121, n6123, n6124, n6126, n6127,
    n6128, n6130, n6131, n6132, n6134, n6135, n6136, n6138, n6139, n6140,
    n6142, n6143, n6144, n6146, n6147, n6149, n6150, n6151, n6153, n6154,
    n6156, n6157, n6158, n6160, n6161, n6162, n6164, n6165, n6166, n6168,
    n6169, n6171, n6172, n6174, n6175, n6177, n6178, n6180, n6181, n6182,
    n6184, n6185, n6186, n6188, n6189, n6190, n6192, n6193, n6194, n6196,
    n6197, n6198, n6200, n6201, n6202, n6204, n6205, n6206, n6208, n6209,
    n6210, n6212, n6213, n6214, n6216, n6217, n6218, n6220, n6221, n6222,
    n6224, n6225, n6227, n6228, n6230, n6231, n6233, n6234, n6236, n6237,
    n6238, n6240, n6241, n6242, n6244, n6245, n6246, n6248, n6249, n6250,
    n6252, n6253, n6254, n6256, n6257, n6258, n6259, n6260, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6287, n6288, n6289, n6291, n6292, n6293, n6295, n6296,
    n6297, n6299, n6300, n6301, n6303, n6304, n6305, n6306, n6307, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6333, n6334, n6335, n6336, n6338, n6339, n6340, n6342,
    n6343, n6344, n6346, n6347, n6348, n6350, n6351, n6352, n6354, n6355,
    n6356, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6367,
    n6368, n6370, n6371, n6372, n6374, n6375, n6376, n6378, n6379, n6380,
    n6382, n6383, n6384, n6386, n6387, n6388, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6414,
    n6415, n6417, n6418, n6419, n6421, n6422, n6423, n6425, n6426, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6438, n6439, n6441,
    n6442, n6444, n6445, n6447, n6448, n6449, n6451, n6452, n6453, n6455,
    n6456, n6457, n6459, n6460, n6462, n6463, n6465, n6466, n6468, n6469,
    n6470, n6472, n6473, n6474, n6476, n6477, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6487, n6488, n6490, n6491, n6493, n6494, n6496,
    n6497, n6498, n6500, n6501, n6502, n6504, n6505, n6506, n6508, n6509,
    n6510, n6512, n6513, n6515, n6516, n6518, n6519, n6521, n6522, n6523,
    n6525, n6526, n6527, n6528, n6529, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6539, n6540, n6542, n6543, n6544, n6546, n6547, n6549,
    n6550, n6551, n6553, n6554, n6555, n6557, n6558, n6559, n6561, n6562,
    n6563, n6565, n6566, n6568, n6569, n6571, n6572, n6574, n6575, n6576,
    n6578, n6579, n6580, n6581, n6582, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6592, n6593, n6594, n6596, n6597, n6598, n6600, n6601,
    n6602, n6604, n6605, n6607, n6608, n6610, n6611, n6612, n6614, n6615,
    n6616, n6618, n6619, n6620, n6622, n6623, n6624, n6626, n6627, n6629,
    n6630, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
    n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
    n6682, n6683, n6685, n6686, n6687, n6689, n6690, n6691, n6693, n6694,
    n6695, n6697, n6698, n6699, n6701, n6703, n6704, n6705, n6707, n6708,
    n6710, n6711, n6713, n6714, n6715, n6717, n6718, n6720, n6721, n6723,
    n6724, n6725, n6727, n6728, n6730, n6731, n6733, n6734, n6735, n6737,
    n6738, n6739, n6741, n6742, n6743, n6745, n6746, n6747, n6749, n6750,
    n6752, n6753, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
    n6773, n6774, n6775, n6776, n6777, n6778, n6780, n6781, n6782, n6783,
    n6784, n6785, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6798, n6799, n6800, n6802, n6803, n6804, n6806, n6807,
    n6808, n6810, n6812, n6813, n6814, n6816, n6817, n6819, n6820, n6822,
    n6823, n6824, n6826, n6827, n6829, n6830, n6832, n6833, n6835, n6836,
    n6837, n6839, n6840, n6842, n6843, n6844, n6846, n6847, n6848, n6850,
    n6851, n6852, n6854, n6855, n6856, n6858, n6859, n6861, n6862, n6864,
    n6865, n6867, n6868, n6869, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
    n6918, n6919, n6920, n6921, n6922, n6923, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934, n6936, n6937, n6938, n6940,
    n6941, n6942, n6944, n6945, n6946, n6948, n6950, n6951, n6952, n6954,
    n6955, n6956, n6958, n6959, n6961, n6962, n6964, n6965, n6966, n6968,
    n6969, n6970, n6972, n6973, n6975, n6976, n6978, n6979, n6980, n6982,
    n6983, n6985, n6986, n6988, n6989, n6990, n6992, n6993, n6994, n6996,
    n6997, n6998, n7000, n7001, n7003, n7004, n7006, n7007, n7009, n7010,
    n7011, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
    n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7037, n7038, n7039, n7040, n7041, n7042,
    n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
    n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7101, n7102, n7103, n7105, n7106,
    n7107, n7109, n7110, n7111, n7113, n7114, n7115, n7117, n7119, n7120,
    n7121, n7123, n7124, n7125, n7127, n7128, n7130, n7131, n7133, n7134,
    n7135, n7137, n7138, n7139, n7141, n7142, n7144, n7145, n7147, n7148,
    n7149, n7151, n7152, n7154, n7155, n7157, n7158, n7159, n7161, n7162,
    n7163, n7165, n7166, n7167, n7169, n7170, n7172, n7173, n7175, n7176,
    n7178, n7179, n7180, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
    n7230, n7231, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7259, n7260, n7261,
    n7262, n7263, n7264, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7309, n7310, n7311, n7313, n7314, n7315,
    n7317, n7318, n7320, n7322, n7323, n7324, n7326, n7327, n7328, n7330,
    n7331, n7333, n7334, n7335, n7337, n7339, n7340, n7342, n7343, n7344,
    n7346, n7347, n7348, n7350, n7351, n7353, n7354, n7355, n7357, n7358,
    n7359, n7361, n7362, n7363, n7365, n7366, n7368, n7369, n7370, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
    n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7449, n7450, n7451, n7452, n7453, n7454, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7499, n7500, n7501, n7503, n7504, n7505, n7507, n7508, n7509, n7511,
    n7513, n7514, n7515, n7517, n7518, n7519, n7521, n7522, n7524, n7525,
    n7526, n7528, n7530, n7531, n7533, n7534, n7536, n7537, n7538, n7540,
    n7541, n7543, n7544, n7545, n7547, n7548, n7549, n7551, n7552, n7553,
    n7555, n7556, n7558, n7559, n7560, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634, n7636, n7637, n7638, n7639,
    n7640, n7641, n7643, n7644, n7645, n7646, n7647, n7648, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7682,
    n7683, n7684, n7686, n7687, n7688, n7690, n7691, n7692, n7694, n7696,
    n7698, n7699, n7700, n7702, n7703, n7705, n7706, n7707, n7709, n7711,
    n7712, n7714, n7715, n7717, n7718, n7719, n7721, n7722, n7723, n7725,
    n7726, n7727, n7729, n7730, n7732, n7733, n7734, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7814, n7815, n7816, n7817, n7818, n7819, n7821, n7822,
    n7823, n7824, n7825, n7826, n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
    n7854, n7855, n7856, n7857, n7858, n7860, n7861, n7862, n7864, n7865,
    n7866, n7868, n7869, n7870, n7872, n7874, n7876, n7877, n7878, n7880,
    n7881, n7883, n7884, n7885, n7887, n7888, n7889, n7891, n7892, n7894,
    n7895, n7897, n7898, n7899, n7901, n7902, n7903, n7905, n7906, n7908,
    n7909, n7910, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7962, n7963, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978, n7980, n7981, n7982, n7983,
    n7985, n7986, n7988, n7989, n7990, n7991, n7992, n7993, n7996, n7997,
    n7998, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8018, n8019, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048, n8050, n8051, n8052, n8053,
    n8054, n8056, n8058, n8060, n8061, n8062, n8063, n8064, n8066, n8069,
    n8070, n8072, n8073, n8074, n8075, n8076, n8078, n8079, n8080, n8081,
    n8082, n8085, n8087, n8088, n8089, n8090, n8091, n8093, n8096, n8097,
    n8099, n8100, n8101, n8102, n8103, n8105, n8106, n8109, n8111, n8112,
    n8113, n8114, n8115, n8117, n8118, n8121, n8122, n8123, n8124, n8125,
    n8127, n8130, n8132, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8163, n8165, n8166, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8197, n8199, n8200, n8201, n8202, n8203, n8206, n8208,
    n8209, n8211, n8212, n8213, n8214, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8265, n8267, n8268, n8269, n8271, n8272, n8273, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8304, n8306, n8309,
    n8310, n8311, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8343, n8344, n8345, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
    n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8378, n8380, n8381, n8382, n8383, n8384, n8386, n8387,
    n8388, n8389, n8390, n8392, n8395, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8411, n8413,
    n8415, n8417, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8455, n8457, n8458,
    n8459, n8460, n8461, n8463, n8465, n8467, n8469, n8470, n8471, n8472,
    n8473, n8475, n8477, n8479, n8480, n8481, n8482, n8484, n8486, n8488,
    n8490, n8491, n8493, n8495, n8496, n8497, n8499, n8501, n8503, n8505,
    n8507, n8508, n8509, n8511, n8513, n8514, n8515, n8516, n8517, n8519,
    n8521, n8523, n8524, n8525, n8527, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
    n8554, n8555, n8556, n8557, n8558, n8560, n8561, n8562, n8564, n8565,
    n8567, n8569, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8602, n8603, n8604, n8605, n8606, n8608, n8610, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8641, n8644, n8645,
    n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671, n8673, n8674, n8677, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8737, n8738, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8769, n8771, n8774, n8775, n8776,
    n8777, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n274, n279, n283, n287, n291, n296, n301, n305,
    n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n359, n364,
    n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419, n424,
    n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484,
    n489, n494, n499, n504, n509, n514, n518, n522, n527, n532, n536, n540,
    n545, n550, n555, n560, n565, n570, n575, n580, n585, n590, n595, n600,
    n605, n610, n615, n620, n625, n630, n635, n640, n645, n650, n655, n660,
    n665, n670, n675, n680, n685, n690, n695, n700, n705, n710, n715, n720,
    n725, n730, n735, n740, n744, n748, n753, n757, n761, n765, n770, n775,
    n780, n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835,
    n840, n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895,
    n900, n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955,
    n960, n965, n969, n973, n978, n982, n986, n990, n995, n1000, n1005,
    n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055,
    n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1095, n1100, n1105,
    n1110, n1115, n1120, n1125, n1130, n1135, n1140, n1145, n1150, n1155,
    n1160, n1165, n1170, n1175, n1180, n1184, n1188, n1192, n1197, n1202,
    n1207, n1212, n1217, n1222, n1227, n1232, n1237, n1242, n1247, n1252,
    n1257, n1262, n1267, n1272, n1277, n1282, n1287, n1292, n1297, n1302,
    n1307, n1312, n1317, n1322, n1327, n1332, n1337, n1342, n1347, n1352,
    n1357, n1362, n1367, n1372, n1377, n1382, n1386, n1390, n1394, n1399,
    n1404, n1409, n1414, n1419, n1424, n1429, n1434, n1439, n1444, n1449,
    n1454, n1459, n1464, n1469, n1474, n1479, n1484, n1489, n1494, n1499,
    n1504, n1509, n1514, n1519, n1524, n1529, n1534, n1539, n1544, n1549,
    n1554, n1559, n1564, n1569, n1574, n1579, n1584, n1588, n1592, n1596,
    n1601, n1606, n1611, n1616, n1621, n1626, n1631, n1636, n1641, n1646,
    n1651, n1656, n1661, n1666, n1671, n1676, n1681, n1686, n1691, n1696,
    n1701, n1706, n1711, n1716, n1721, n1726, n1731, n1736, n1741, n1746,
    n1751, n1756, n1761, n1766, n1771, n1776, n1781, n1786, n1791, n1795,
    n1799, n1803, n1807, n1812, n1817, n1822, n1827, n1832, n1837, n1842,
    n1847, n1852, n1857, n1862, n1867, n1872, n1877, n1882, n1887, n1892,
    n1897, n1902, n1907, n1912, n1917, n1922, n1927, n1932, n1937, n1942,
    n1947, n1952, n1957, n1962, n1967, n1972, n1977, n1982, n1987, n1992,
    n1997, n2002, n2007, n2012, n2017, n2021, n2026, n2031, n2036, n2041,
    n2046, n2051, n2056, n2061, n2066, n2071, n2076, n2081, n2086, n2091,
    n2096, n2101, n2106, n2111, n2116, n2121, n2126, n2131, n2136, n2141,
    n2146, n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2185, n2189,
    n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2229, n2234, n2239,
    n2244, n2249, n2254, n2259, n2264, n2268, n2272, n2277, n2282, n2287,
    n2292, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337,
    n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387,
    n2392, n2397, n2402, n2407, n2412, n2417, n2422, n2427, n2432, n2437,
    n2442, n2447, n2452, n2457, n2462, n2467, n2472, n2477, n2482, n2487,
    n2492, n2497, n2502, n2507, n2512, n2517, n2522, n2527, n2532, n2537,
    n2542, n2547, n2552, n2557, n2562, n2567, n2572, n2577, n2582, n2587,
    n2592, n2597, n2602, n2607, n2612, n2617, n2622, n2627, n2632, n2637,
    n2642, n2647, n2652, n2657, n2662, n2667, n2671, n2675, n2680, n2685,
    n2690, n2695, n2699, n2703, n2708, n2713, n2718, n2723, n2728, n2733,
    n2737, n2742, n2747, n2752, n2757, n2762, n2767, n2771, n2776, n2781,
    n2786, n2790, n2794, n2799, n2804, n2809, n2814, n2819, n2824, n2829,
    n2834, n2839, n2844, n2849, n2853, n2857, n2862, n2867, n2872, n2877,
    n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2916, n2920, n2925,
    n2930, n2935, n2940, n2945, n2950, n2955, n2960, n2965, n2970, n2975,
    n2979, n2983, n2988, n2993, n2998, n3003, n3008, n3013, n3018, n3023,
    n3028, n3033, n3038, n3042, n3046, n3051, n3056, n3061, n3066, n3071,
    n3076, n3081, n3086, n3091, n3096, n3101, n3106, n3111, n3116, n3121,
    n3126, n3131, n3136, n3141, n3146, n3150, n3155, n3159, n3164, n3169,
    n3174, n3179, n3184, n3189, n3194, n3199, n3204, n3209, n3214, n3219,
    n3224, n3229, n3234, n3239, n3244, n3249, n3254, n3259, n3264, n3268,
    n3272, n3276, n3281, n3286, n3291, n3296, n3301, n3306, n3311, n3316,
    n3321, n3326, n3331, n3336, n3341, n3346, n3351, n3356, n3361, n3366,
    n3371, n3376, n3381, n3386, n3390, n3394, n3398, n3402, n3407, n3412,
    n3417, n3422, n3427, n3432, n3437, n3442, n3447, n3452, n3457, n3462,
    n3467, n3472, n3477, n3482, n3487, n3492, n3497, n3502, n3507, n3512,
    n3517, n3521, n3525, n3529, n3534, n3538, n3542, n3547, n3552, n3557,
    n3562, n3567, n3572, n3577, n3582, n3587, n3592, n3597, n3602, n3607,
    n3612, n3617, n3622, n3627, n3632, n3636, n3640, n3644, n3649, n3653,
    n3657, n3662, n3667, n3672, n3677, n3682, n3687, n3692, n3697, n3702,
    n3707, n3712, n3717, n3722, n3727, n3732, n3737, n3742, n3747, n3751,
    n3755, n3759, n3764, n3769, n3773, n3778, n3783, n3788, n3793, n3798,
    n3803, n3808, n3813, n3818, n3823, n3828, n3833, n3838, n3843, n3848,
    n3853, n3857, n3861, n3865, n3870, n3875, n3879, n3884, n3889, n3894,
    n3899, n3904, n3909, n3914, n3919, n3924, n3929, n3934, n3939, n3944,
    n3949, n3954, n3958, n3963, n3968, n3973, n3977, n3982, n3987, n3992,
    n3997, n4002, n4007, n4012, n4017, n4022, n4027, n4032, n4037, n4042,
    n4047, n4052, n4057, n4062, n4067, n4072, n4077, n4082, n4087, n4092,
    n4097, n4102, n4107, n4112, n4117, n4122, n4127, n4132, n4137, n4142,
    n4147, n4151, n4156, n4161, n4166, n4170, n4175, n4180, n4185, n4190,
    n4195, n4200, n4204, n4209, n4214, n4219, n4224, n4228, n4233, n4238,
    n4243, n4248, n4252, n4257, n4262, n4266, n4271, n4276, n4281, n4286,
    n4291, n4296, n4301, n4305, n4310, n4315, n4320, n4325, n4329, n4334,
    n4339, n4344, n4349, n4354, n4359, n4364, n4369, n4374, n4379, n4384,
    n4388, n4393, n4398, n4403, n4408, n4413, n4418, n4423, n4428, n4433,
    n4438, n4443, n4448, n4453, n4458, n4463, n4467, n4471, n4476, n4481,
    n4486, n4490, n4495, n4500, n4505, n4510, n4515, n4519, n4524, n4529,
    n4534, n4538, n4543, n4548, n4553, n4558, n4562, n4566, n4571, n4575,
    n4580, n4585, n4590, n4595, n4599;
  assign n2795 = \[16959]  & \[17882] ;
  assign n2796 = tin_pdata_8_8_ & ~\[17882] ;
  assign pdata_8_8_ = n2795 | n2796;
  assign n2798 = \[17479]  & \[18337] ;
  assign n2799_1 = tin_pdata_0_0_ & ~\[17479] ;
  assign pdata_0_0_ = n2798 | n2799_1;
  assign n2801 = \[16907]  & \[17869] ;
  assign n2802 = tin_pdata_7_7_ & ~\[17869] ;
  assign pdata_7_7_ = n2801 | n2802;
  assign n2804_1 = \[17323]  & \[18181] ;
  assign n2805 = tin_pdata_2_2_ & ~\[18181] ;
  assign pdata_2_2_ = n2804_1 | n2805;
  assign n2807 = \[17765]  & \[18571] ;
  assign n2808 = tin_pdata_9_9_ & ~\[18571] ;
  assign pdata_9_9_ = n2807 | n2808;
  assign n2810 = \[17258]  & \[18116] ;
  assign n2811 = tin_pdata_1_1_ & ~\[18116] ;
  assign pdata_1_1_ = n2810 | n2811;
  assign n2813 = \[17193]  & \[18038] ;
  assign n2814_1 = tin_pdata_4_4_ & ~\[18038] ;
  assign pdata_4_4_ = n2813 | n2814_1;
  assign n2816 = \[17011]  & \[17921] ;
  assign n2817 = tin_pdata_10_10_ & ~\[17011] ;
  assign pdata_10_10_ = n2816 | n2817;
  assign n2819_1 = \[17128]  & \[17960] ;
  assign n2820 = tin_pdata_3_3_ & ~\[17960] ;
  assign pdata_3_3_ = n2819_1 | n2820;
  assign n2822 = \[17063]  & \[17934] ;
  assign n2823 = tin_pdata_6_6_ & ~\[17934] ;
  assign pdata_6_6_ = n2822 | n2823;
  assign n2825 = \[17076]  & \[17947] ;
  assign n2826 = tin_pdata_15_15_ & ~\[17947] ;
  assign pdata_15_15_ = n2825 | n2826;
  assign n2828 = \[17336]  & \[18194] ;
  assign n2829_1 = tin_pdata_11_11_ & ~\[17336] ;
  assign pdata_11_11_ = n2828 | n2829_1;
  assign n2831 = \[17778]  & \[18584] ;
  assign n2832 = tin_pdata_14_14_ & ~\[18584] ;
  assign pdata_14_14_ = n2831 | n2832;
  assign n2834_1 = \[17141]  & \[17973] ;
  assign n2835 = tin_pdata_12_12_ & ~\[17141] ;
  assign pdata_12_12_ = n2834_1 | n2835;
  assign n2837 = \[16998]  & \[17908] ;
  assign n2838 = tin_pdata_5_5_ & ~\[17908] ;
  assign pdata_5_5_ = n2837 | n2838;
  assign n2840 = \[17492]  & \[18350] ;
  assign n2841 = tin_pdata_13_13_ & ~\[18350] ;
  assign pdata_13_13_ = n2840 | n2841;
  assign n2843 = \[17791]  & ~\[17843] ;
  assign n2844_1 = ~ndout & ~n2843;
  assign n2845 = ~pdata_2_2_ & n2843;
  assign n2846 = ~preset & ~n2845;
  assign n274 = ~n2844_1 & n2846;
  assign n2848 = \[17531]  & \[18155] ;
  assign n2849_1 = ppeaki_0_0_ & ~\[17531] ;
  assign n2850 = ~n2848 & ~n2849_1;
  assign n2851 = \[17531]  & \[18090] ;
  assign n2852 = ppeaki_3_3_ & ~\[17531] ;
  assign n2853_1 = ~n2851 & ~n2852;
  assign n2854 = \[17531]  & \[18012] ;
  assign n2855 = ppeaki_2_2_ & ~\[17531] ;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857_1 = n2853_1 & n2856;
  assign n2858 = \[17531]  & \[18233] ;
  assign n2859 = ppeaki_1_1_ & ~\[17531] ;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = n2857_1 & n2860;
  assign n2862_1 = ~n2850 & n2861;
  assign n2863 = ~\[17609]  & \[17752] ;
  assign n2864 = ~\[17544]  & n2863;
  assign n2865 = ~\[17674]  & n2864;
  assign n2866 = ~ppeaki_6_6_ & ~\[17752] ;
  assign n2867_1 = ~ppeaki_7_7_ & n2866;
  assign n2868 = ~ppeaki_5_5_ & n2867_1;
  assign n2869 = ~n2865 & ~n2868;
  assign n2870 = n2862_1 & n2869;
  assign n2871 = n2853_1 & ~n2856;
  assign n2872_1 = n2850 & n2860;
  assign n2873 = ~n2853_1 & n2856;
  assign n2874 = n2872_1 & ~n2873;
  assign n2875 = ~n2871 & n2874;
  assign n2876 = \[17596]  & ~\[18597] ;
  assign n2877_1 = ~\[17661]  & n2876;
  assign n2878 = ~\[18636]  & n2877_1;
  assign n2879 = ~n2875 & n2878;
  assign n2880 = ~n2870 & n2879;
  assign n2881 = ~\[18636]  & ~n2877_1;
  assign n2882_1 = ~n2880 & ~n2881;
  assign n2883 = ~\[17089]  & pdn;
  assign n2884 = ~\[17856]  & \[18207] ;
  assign n2885 = ~\[10805]  & ~\[18207] ;
  assign n2886 = ~\[11345]  & ~\[12695] ;
  assign n2887_1 = ~\[12080]  & n2886;
  assign n2888 = n2885 & n2887_1;
  assign n2889 = ~\[11930]  & ~\[12275] ;
  assign n2890 = ~\[10820]  & ~\[11585] ;
  assign n2891 = ~\[11090]  & n2890;
  assign n2892_1 = ~\[12185]  & ~\[12200] ;
  assign n2893 = ~\[12065]  & n2892_1;
  assign n2894 = n2891 & n2893;
  assign n2895 = ~\[11810]  & ~\[12935] ;
  assign n2896 = ~\[11600]  & n2895;
  assign n2897_1 = ~\[12485]  & n2896;
  assign n2898 = n2894 & n2897_1;
  assign n2899 = n2889 & n2898;
  assign n2900 = n2888 & n2899;
  assign n2901 = ~n2884 & ~n2900;
  assign n2902_1 = \[17986]  & n2901;
  assign n2903 = ~\[17804]  & n2902_1;
  assign n2904 = ~\[17596]  & n2903;
  assign n2905 = ~n2883 & ~n2904;
  assign n2906 = ~n2882_1 & n2905;
  assign n2907_1 = ~preset & n2882_1;
  assign n2908 = n2862_1 & n2907_1;
  assign n2909 = ~ppeaki_4_4_ & n2868;
  assign n2910 = ~\[17713]  & n2865;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912_1 = n2908 & ~n2911;
  assign n2913 = \[6470]  & n2912_1;
  assign n2914 = ~n2850 & n2860;
  assign n2915 = ~n2853_1 & ~n2856;
  assign n2916_1 = n2914 & n2915;
  assign n2917 = n2907_1 & n2916_1;
  assign n2918 = \[9230]  & n2917;
  assign n2919 = ~n2913 & ~n2918;
  assign n2920_1 = ~preset & n2904;
  assign n2921 = ~preset_0_0_ & ~\[17024] ;
  assign n2922 = \[17024]  & ~\[18545] ;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2901 & ~n2923;
  assign n2925_1 = ~preset & n2883;
  assign n2926 = n2924 & n2925_1;
  assign n2927 = ~n2920_1 & ~n2926;
  assign n2928 = \[18064]  & \[18129] ;
  assign n2929 = pirq_0_0_ & ~\[18064] ;
  assign n2930_1 = ~n2928 & ~n2929;
  assign n2931 = ~n2927 & ~n2930_1;
  assign n2932 = \[15845]  & n2931;
  assign n2933 = \[17713]  & n2865;
  assign n2934 = ppeaki_4_4_ & n2868;
  assign n2935_1 = ~n2933 & ~n2934;
  assign n2936 = n2908 & ~n2935_1;
  assign n2937 = \[15545]  & n2936;
  assign n2938 = n2850 & ~n2860;
  assign n2939 = n2873 & n2938;
  assign n2940_1 = n2907_1 & n2939;
  assign n2941 = \[5945]  & n2940_1;
  assign n2942 = ~n2937 & ~n2941;
  assign n2943 = ~n2932 & n2942;
  assign n2944 = n2919 & n2943;
  assign n2945_1 = ~n2906 & ~n2944;
  assign n2946 = n2850 & ~n2853_1;
  assign n2947 = n2856 & ~n2946;
  assign n2948 = ~n2860 & n2947;
  assign n2949 = n2871 & n2914;
  assign n2950_1 = ~n2948 & ~n2949;
  assign n2951 = ppeaka_12_12_ & ~n2950_1;
  assign n2952 = n2873 & n2914;
  assign n2953 = \[13325]  & n2952;
  assign n2954 = ~n2850 & ~n2860;
  assign n2955_1 = n2871 & n2954;
  assign n2956 = \[8495]  & n2955_1;
  assign n2957 = ~n2953 & ~n2956;
  assign n2958 = n2860 & n2946;
  assign n2959 = n2856 & n2958;
  assign n2960_1 = \[15260]  & n2959;
  assign n2961 = n2871 & n2872_1;
  assign n2962 = \[6545]  & n2961;
  assign n2963 = ~n2960_1 & ~n2962;
  assign n2964 = n2915 & n2938;
  assign n2965_1 = \[7955]  & n2964;
  assign n2966 = n2963 & ~n2965_1;
  assign n2967 = n2957 & n2966;
  assign n2968 = ~n2951 & n2967;
  assign n2969 = n2907_1 & ~n2968;
  assign n2970_1 = ppeaki_5_5_ & n2867_1;
  assign n2971 = ~ppeaki_4_4_ & n2970_1;
  assign n2972 = ~\[17713]  & n2864;
  assign n2973 = \[17674]  & n2972;
  assign n2974 = ~n2971 & ~n2973;
  assign n2975_1 = n2908 & ~n2974;
  assign n2976 = ~n2856 & n2907_1;
  assign n2977 = n2853_1 & n2938;
  assign n2978 = ~n2914 & ~n2938;
  assign n2979_1 = ~n2853_1 & n2978;
  assign n2980 = ~n2977 & ~n2979_1;
  assign n2981 = n2976 & ~n2980;
  assign n2982 = ~n2975_1 & ~n2981;
  assign n2983_1 = n2883 & ~n2924;
  assign n2984 = ~n2906 & ~n2983_1;
  assign n2985 = ~preset & ~n2984;
  assign n2986 = ~preset & n2930_1;
  assign n2987 = ~n2905 & n2986;
  assign n2988_1 = ~n2985 & ~n2987;
  assign n2989 = n2982 & n2988_1;
  assign n2990 = ppeakb_12_12_ & ~n2989;
  assign n2991 = ~n2969 & ~n2990;
  assign n279 = n2945_1 | ~n2991;
  assign n2993_1 = \[15650]  & n2940_1;
  assign n2994 = \[9065]  & n2936;
  assign n2995 = ~n2993_1 & ~n2994;
  assign n2996 = \[5030]  & n2931;
  assign n2997 = \[5285]  & n2917;
  assign n2998_1 = \[5075]  & n2912_1;
  assign n2999 = ~n2997 & ~n2998_1;
  assign n3000 = ~n2996 & n2999;
  assign n3001 = n2995 & n3000;
  assign n3002 = ~n2906 & ~n3001;
  assign n3003_1 = ppeaka_1_1_ & ~n2950_1;
  assign n3004 = \[5150]  & n2961;
  assign n3005 = \[13310]  & n2952;
  assign n3006 = ~n3004 & ~n3005;
  assign n3007 = \[13295]  & n2959;
  assign n3008_1 = \[14510]  & n2964;
  assign n3009 = ~n3007 & ~n3008_1;
  assign n3010 = \[8480]  & n2955_1;
  assign n3011 = n3009 & ~n3010;
  assign n3012 = n3006 & n3011;
  assign n3013_1 = ~n3003_1 & n3012;
  assign n3014 = n2907_1 & ~n3013_1;
  assign n3015 = ppeakb_1_1_ & ~n2989;
  assign n3016 = ~n3014 & ~n3015;
  assign n283 = n3002 | ~n3016;
  assign n3018_1 = \[12560]  & n2936;
  assign n3019 = n2857_1 & ~n2860;
  assign n3020 = n2850 & n3019;
  assign n3021 = n2907_1 & n3020;
  assign n3022 = \[15200]  & n3021;
  assign n3023_1 = n2857_1 & n2954;
  assign n3024 = n2907_1 & n3023_1;
  assign n3025 = \[11690]  & n3024;
  assign n3026 = ~n3022 & ~n3025;
  assign n3027 = ~n3018_1 & n3026;
  assign n3028_1 = ppeaka_6_6_ & ppeakb_6_6_;
  assign n3029 = n2912_1 & ~n3028_1;
  assign n3030 = n2871 & n2938;
  assign n3031 = n2907_1 & n3030;
  assign n3032 = \[5870]  & n3031;
  assign n3033_1 = ~n3029 & ~n3032;
  assign n3034 = n2958 & n2976;
  assign n3035 = ~n2931 & ~n3034;
  assign n3036 = ppeakp_6_6_ & ~n3035;
  assign n3037 = n3033_1 & ~n3036;
  assign n3038_1 = n3027 & n3037;
  assign n3039 = ~n2906 & ~n3038_1;
  assign n3040 = ppeaka_7_7_ & n2975_1;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042_1 = ~n2917 & n2988_1;
  assign n3043 = ppeaka_6_6_ & ~n3042_1;
  assign n3044 = n2915 & n2954;
  assign n3045 = \[4955]  & n3044;
  assign n3046_1 = n2873 & n2954;
  assign n3047 = ~n2949 & ~n3046_1;
  assign n3048 = \[7685]  & ~n3047;
  assign n3049 = n2873 & ~n2954;
  assign n3050 = ~n2955_1 & ~n3049;
  assign n3051_1 = ppeakb_6_6_ & ~n3050;
  assign n3052 = ~n3048 & ~n3051_1;
  assign n3053 = \[10745]  & n2964;
  assign n3054 = \[15935]  & n2961;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056_1 = n3052 & n3055;
  assign n3057 = ~n3045 & n3056_1;
  assign n3058 = n2907_1 & ~n3057;
  assign n3059 = ~n3043 & ~n3058;
  assign n287 = ~n3041 | ~n3059;
  assign n3061_1 = ~n2914 & n2947;
  assign n3062 = ~n2916_1 & ~n3061_1;
  assign n3063 = ~n3019 & ~n3062;
  assign n3064 = n2907_1 & ~n3063;
  assign n3065 = n2988_1 & ~n3064;
  assign n3066_1 = \[4295]  & ~n3065;
  assign n3067 = \[8825]  & n2931;
  assign n3068 = n2907_1 & n3046_1;
  assign n3069 = \[7655]  & n3068;
  assign n3070 = \[8540]  & n2917;
  assign n3071_1 = ~n3069 & ~n3070;
  assign n3072 = ~n3067 & n3071_1;
  assign n291 = n3066_1 | ~n3072;
  assign n3074 = \[4310]  & ~n3065;
  assign n3075 = \[7640]  & n3068;
  assign n3076_1 = ~n3074 & ~n3075;
  assign n3077 = \[14225]  & n2931;
  assign n3078 = \[8525]  & n2917;
  assign n3079 = ~n3077 & ~n3078;
  assign n296 = ~n3076_1 | ~n3079;
  assign n3081_1 = n2907_1 & n2952;
  assign n3082 = \[13055]  & n3081_1;
  assign n3083 = ~preset & n2906;
  assign n3084 = ~n2923 & n2925_1;
  assign n3085 = n2901 & n3084;
  assign n3086_1 = ~n2927 & n2930_1;
  assign n3087 = ~n3085 & ~n3086_1;
  assign n3088 = ~n2906 & ~n3087;
  assign n3089 = n2982 & ~n3088;
  assign n3090 = ~n3083 & n3089;
  assign n3091_1 = ppeaks_5_5_ & ~n3090;
  assign n3092 = \[15395]  & n2931;
  assign n3093 = \[11465]  & n3024;
  assign n3094 = \[13700]  & n2912_1;
  assign n3095 = n2923 & n2925_1;
  assign n3096_1 = \[11885]  & n3095;
  assign n3097 = ~n3094 & ~n3096_1;
  assign n3098 = \[14555]  & n2936;
  assign n3099 = \[5420]  & n2955_1;
  assign n3100 = \[10895]  & n2964;
  assign n3101_1 = \[13505]  & n2949;
  assign n3102 = ~n3100 & ~n3101_1;
  assign n3103 = ~n3099 & n3102;
  assign n3104 = \[13430]  & n2939;
  assign n3105 = \[6995]  & n3046_1;
  assign n3106_1 = ~n3104 & ~n3105;
  assign n3107 = \[6185]  & n2916_1;
  assign n3108 = n3106_1 & ~n3107;
  assign n3109 = \[7445]  & n2959;
  assign n3110 = \[10280]  & n2961;
  assign n3111_1 = ~n3109 & ~n3110;
  assign n3112 = \[9545]  & n3020;
  assign n3113 = n3111_1 & ~n3112;
  assign n3114 = n3108 & n3113;
  assign n3115 = n3103 & n3114;
  assign n3116_1 = n2907_1 & ~n3115;
  assign n3117 = ~n3098 & ~n3116_1;
  assign n3118 = n3097 & n3117;
  assign n3119 = ~n3093 & n3118;
  assign n3120 = ~n3092 & n3119;
  assign n3121_1 = ~n2906 & ~n3120;
  assign n3122 = ~n3091_1 & ~n3121_1;
  assign n301 = n3082 | ~n3122;
  assign n3124 = ~n2853_1 & n2860;
  assign n3125 = n2857_1 & ~n2914;
  assign n3126_1 = ~n3124 & ~n3125;
  assign n3127 = ~ppeakb_3_3_ & ~ppeakb_8_8_;
  assign n3128 = ~ppeakb_13_13_ & ~ppeakb_5_5_;
  assign n3129 = ~ppeakb_4_4_ & ~ppeakb_7_7_;
  assign n3130 = n3128 & n3129;
  assign n3131_1 = n3127 & n3130;
  assign n3132 = ~ppeakb_1_1_ & ~ppeakb_9_9_;
  assign n3133 = ~ppeakb_12_12_ & n3132;
  assign n3134 = ~ppeakb_6_6_ & n3133;
  assign n3135 = n3131_1 & n3134;
  assign n3136_1 = ~ppeakb_2_2_ & ~ppeakb_14_14_;
  assign n3137 = ~ppeakb_0_0_ & ~ppeakb_15_15_;
  assign n3138 = ~ppeakb_11_11_ & n3137;
  assign n3139 = ~ppeakb_10_10_ & n3138;
  assign n3140 = n3136_1 & n3139;
  assign n3141_1 = n3135 & n3140;
  assign n3142 = n2952 & n3141_1;
  assign n3143 = ~n3126_1 & ~n3142;
  assign n3144 = n2907_1 & ~n3143;
  assign n3145 = ~n3085 & ~n3144;
  assign n3146_1 = ~n3024 & n3145;
  assign n3147 = ~n3083 & n3146_1;
  assign n3148 = ppeakp_10_10_ & ~n3147;
  assign n3149 = \[4850]  & ~n2927;
  assign n3150_1 = \[12140]  & n3095;
  assign n3151 = ppeakb_10_10_ & n2917;
  assign n3152 = ~n3150_1 & ~n3151;
  assign n3153 = ~n3149 & n3152;
  assign n3154 = n2907_1 & n2958;
  assign n3155_1 = n3081_1 & ~n3141_1;
  assign n3156 = ~n3154 & ~n3155_1;
  assign n3157 = ppeaka_10_10_ & ~n3156;
  assign n3158 = \[6965]  & n3021;
  assign n3159_1 = ~n3157 & ~n3158;
  assign n3160 = n3153 & n3159_1;
  assign n305 = n3148 | ~n3160;
  assign n3162 = \[17453]  & ~\[18246] ;
  assign n3163 = ~\[4355]  & ~n3162;
  assign n3164_1 = ~pdata_0_0_ & n3162;
  assign n3165 = ~preset & ~n3164_1;
  assign n309 = ~n3163 & n3165;
  assign n3167 = ~\[4370]  & ~n3162;
  assign n3168 = ~pdata_11_11_ & n3162;
  assign n3169_1 = ~preset & ~n3168;
  assign n314 = ~n3167 & n3169_1;
  assign n3171 = ~\[18168]  & ~n2935_1;
  assign n3172 = ~\[18610]  & ~n2869;
  assign n3173 = n2862_1 & n2879;
  assign n3174_1 = n3172 & n3173;
  assign n3175 = n3171 & n3174_1;
  assign n3176 = ~\[4385]  & ~n3175;
  assign n3177 = ~preset & pdata_6_6_;
  assign n3178 = ~preset & ~n3175;
  assign n3179_1 = ~n3177 & ~n3178;
  assign n319 = ~n3176 & ~n3179_1;
  assign n3181 = \[17102]  & ~\[17154] ;
  assign n3182 = ~\[4400]  & ~n3181;
  assign n3183 = ~pdata_1_1_ & n3181;
  assign n3184_1 = ~preset & ~n3183;
  assign n324 = ~n3182 & n3184_1;
  assign n3186 = ~\[4415]  & ~n3181;
  assign n3187 = ~pdata_12_12_ & n3181;
  assign n3188 = ~preset & ~n3187;
  assign n329 = ~n3186 & n3188;
  assign n3190 = n2880 & n2961;
  assign n3191 = ~\[18285]  & n3190;
  assign n3192 = ~preset & n3191;
  assign n3193 = pdata_7_7_ & n3192;
  assign n3194_1 = ~preset & ~n3191;
  assign n3195 = \[4430]  & n3194_1;
  assign n334 = n3193 | n3195;
  assign n3197 = pdata_2_2_ & n3192;
  assign n3198 = \[4445]  & n3194_1;
  assign n339 = n3197 | n3198;
  assign n3200 = pdata_13_13_ & n3192;
  assign n3201 = \[4460]  & n3194_1;
  assign n344 = n3200 | n3201;
  assign n3203 = \[17167]  & ~\[17362] ;
  assign n3204_1 = ~\[4475]  & ~n3203;
  assign n3205 = ~pdata_8_8_ & n3203;
  assign n3206 = ~preset & ~n3205;
  assign n349 = ~n3204_1 & n3206;
  assign n3208 = \[17284]  & ~\[18376] ;
  assign n3209_1 = ~pdata_3_3_ & n3208;
  assign n3210 = ~\[4490]  & ~n3208;
  assign n3211 = ~preset & ~n3210;
  assign n354 = ~n3209_1 & n3211;
  assign n3213 = ~pdata_14_14_ & n3208;
  assign n3214_1 = ~\[4505]  & ~n3208;
  assign n3215 = ~preset & ~n3214_1;
  assign n359 = ~n3213 & n3215;
  assign n3217 = ~\[18493]  & n2959;
  assign n3218 = n2880 & n3217;
  assign n3219_1 = ~\[4520]  & ~n3218;
  assign n3220 = ~pdata_9_9_ & n3218;
  assign n3221 = ~preset & ~n3220;
  assign n364 = ~n3219_1 & n3221;
  assign n3223 = ~\[16920]  & n2880;
  assign n3224_1 = n2952 & n3223;
  assign n3225 = ~preset & ~n3224_1;
  assign n3226 = \[4535]  & n3225;
  assign n3963 = ~preset & n3224_1;
  assign n3228 = pdata_15_15_ & n3963;
  assign n369 = n3226 | n3228;
  assign n3230 = ~\[17297]  & n2939;
  assign n3231 = n2880 & n3230;
  assign n3232 = ~\[4550]  & ~n3231;
  assign n3233 = ~pdata_10_10_ & n3231;
  assign n3234_1 = ~preset & ~n3233;
  assign n374 = ~n3232 & n3234_1;
  assign n3236 = n2880 & n2916_1;
  assign n3237 = ~\[18506]  & n3236;
  assign n3238 = ~preset & n3237;
  assign n3239_1 = pdata_5_5_ & n3238;
  assign n3240 = ~preset & ~n3237;
  assign n3241 = \[4565]  & n3240;
  assign n379 = n3239_1 | n3241;
  assign n3243 = pdata_0_0_ & n3238;
  assign n3244_1 = \[4580]  & n3240;
  assign n384 = n3243 | n3244_1;
  assign n3246 = pdata_11_11_ & n3238;
  assign n3247 = \[4595]  & n3240;
  assign n389 = n3246 | n3247;
  assign n3249_1 = ~\[17310]  & \[17388] ;
  assign n3250 = ~\[4610]  & ~n3249_1;
  assign n3251 = ~pdata_6_6_ & n3249_1;
  assign n3252 = ~preset & ~n3251;
  assign n394 = ~n3250 & n3252;
  assign n3254_1 = ~\[17453]  & ~n2911;
  assign n3255 = ~preset & n2880;
  assign n3256 = n2862_1 & n3255;
  assign n3257 = n3172 & n3256;
  assign n4161 = n3254_1 & n3257;
  assign n3259_1 = ~n3191 & ~n3237;
  assign n3260 = n3174_1 & n3254_1;
  assign n3261 = ~n3231 & ~n3260;
  assign n3262 = ~n3218 & ~n3224_1;
  assign n3263 = n3261 & n3262;
  assign n3264_1 = n3259_1 & n3263;
  assign n3265 = ~\[18103]  & \[18168] ;
  assign n3266 = \[18285]  & ~\[18363] ;
  assign n3267 = ~\[18311]  & \[18506] ;
  assign n3268_1 = ~n3266 & ~n3267;
  assign n3269 = ~n3265 & n3268_1;
  assign n3270 = n3264_1 & n3269;
  assign n3271 = ppeaka_0_0_ & n3175;
  assign n3272_1 = ~\[17284]  & n2880;
  assign n3273 = n2955_1 & n3272_1;
  assign n3274 = n2880 & n2964;
  assign n3275 = ~\[16933]  & n3274;
  assign n3276_1 = ~n3273 & ~n3275;
  assign n3277 = ~n3271 & n3276_1;
  assign n3278 = n3270 & n3277;
  assign n3279 = ppeakb_0_0_ & n3175;
  assign n3280 = \[4310]  & n3237;
  assign n3281_1 = ~n3279 & ~n3280;
  assign n3282 = ppeaka_0_0_ & n3191;
  assign n3283 = \[8630]  & n3266;
  assign n3284 = \[10025]  & n3267;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286_1 = ~n3282 & n3285;
  assign n3287 = n3281_1 & n3286_1;
  assign n3288 = n3263 & ~n3265;
  assign n3289 = n3276_1 & n3288;
  assign n3290 = ppeaks_0_0_ & ~n3289;
  assign n3291_1 = n3287 & ~n3290;
  assign n3292 = ~n3278 & n3291_1;
  assign n3293 = ppeaks_1_1_ & ~n3289;
  assign n3294 = \[5030]  & n3237;
  assign n3295 = ppeaka_1_1_ & n3191;
  assign n3296_1 = ~n3294 & ~n3295;
  assign n3297 = \[10310]  & n3267;
  assign n3298 = \[9290]  & n3266;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ppeakb_1_1_ & n3175;
  assign n3301_1 = n3299 & ~n3300;
  assign n3302 = n3296_1 & n3301_1;
  assign n3303 = ~n3293 & n3302;
  assign n3304 = ppeaka_1_1_ & n3175;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306_1 = n3303 & n3304;
  assign n3307 = ~n3305 & ~n3306_1;
  assign n3308 = ~n3292 & ~n3307;
  assign n3309 = n3292 & n3307;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311_1 = n4161 & ~n3310;
  assign n3312 = ~preset & ~n3260;
  assign n3313 = \[4625]  & n3312;
  assign n399 = n3311_1 | n3313;
  assign n3315 = ppeaks_12_12_ & ~n3289;
  assign n3316_1 = \[15845]  & n3237;
  assign n3317 = \[10010]  & n3266;
  assign n3318 = \[6860]  & n3267;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = ~n3316_1 & n3319;
  assign n3321_1 = ppeaka_12_12_ & n3191;
  assign n3322 = ppeakb_12_12_ & n3175;
  assign n3323 = ~n3321_1 & ~n3322;
  assign n3324 = n3320 & n3323;
  assign n3325 = ~n3315 & n3324;
  assign n3326_1 = ~n3175 & n3278;
  assign n3327 = n3278 & ~n3304;
  assign n3328 = ~ppeaka_2_2_ & n3327;
  assign n3329 = ~ppeaka_3_3_ & n3328;
  assign n3330 = ~n3326_1 & ~n3329;
  assign n3331_1 = ppeaka_4_4_ & n3175;
  assign n3332 = ~n3330 & ~n3331_1;
  assign n3333 = ~ppeaka_5_5_ & n3332;
  assign n3334 = ~ppeaka_6_6_ & n3333;
  assign n3335 = ~n3326_1 & ~n3334;
  assign n3336_1 = ~n3175 & n3335;
  assign n3337 = ppeaka_7_7_ & n3175;
  assign n3338 = ~n3335 & ~n3337;
  assign n3339 = ~ppeaka_8_8_ & n3338;
  assign n3340 = ~ppeaka_9_9_ & n3339;
  assign n3341_1 = ppeaka_10_10_ & n3175;
  assign n3342 = n3340 & ~n3341_1;
  assign n3343 = ~n3175 & ~n3335;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~ppeaka_11_11_ & ~n3344;
  assign n3346_1 = ppeaka_12_12_ & ~n3345;
  assign n3347 = ~ppeaka_12_12_ & n3345;
  assign n3348 = ~n3343 & ~n3347;
  assign n3349 = ~n3346_1 & n3348;
  assign n3350 = ~n3336_1 & ~n3349;
  assign n3351_1 = ~n3325 & ~n3350;
  assign n3352 = n3325 & n3350;
  assign n3353 = ~n3351_1 & ~n3352;
  assign n3354 = ppeaks_11_11_ & ~n3289;
  assign n3355 = \[4295]  & n3237;
  assign n3356_1 = \[10595]  & n3267;
  assign n3357 = \[8645]  & n3266;
  assign n3358 = ~n3356_1 & ~n3357;
  assign n3359 = ~n3355 & n3358;
  assign n3360 = ppeaka_11_11_ & n3191;
  assign n3361_1 = ppeakb_11_11_ & n3175;
  assign n3362 = ~n3360 & ~n3361_1;
  assign n3363 = n3359 & n3362;
  assign n3364 = ~n3354 & n3363;
  assign n3365 = ppeaka_11_11_ & n3175;
  assign n3366_1 = ~n3342 & n3365;
  assign n3367 = ~n3344 & ~n3365;
  assign n3368 = ~n3366_1 & ~n3367;
  assign n3369 = ~n3364 & n3368;
  assign n3370 = n3364 & ~n3368;
  assign n3371_1 = ~n3340 & n3341_1;
  assign n3372 = n3344 & ~n3371_1;
  assign n3373 = ppeaks_9_9_ & ~n3289;
  assign n3374 = \[5720]  & n3237;
  assign n3375 = ppeaka_9_9_ & n3191;
  assign n3376_1 = ~n3374 & ~n3375;
  assign n3377 = \[7370]  & n3266;
  assign n3378 = \[10040]  & n3267;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = ppeakb_9_9_ & n3175;
  assign n3381_1 = n3379 & ~n3380;
  assign n3382 = n3376_1 & n3381_1;
  assign n3383 = ~n3373 & n3382;
  assign n3384 = ppeaka_9_9_ & ~n3339;
  assign n3385 = ~n3340 & ~n3384;
  assign n3386_1 = n3175 & n3385;
  assign n3387 = ~n3336_1 & ~n3386_1;
  assign n3388 = ~n3383 & ~n3387;
  assign n3389 = n3383 & n3387;
  assign n3390_1 = ppeaks_8_8_ & ~n3289;
  assign n3391 = \[6410]  & n3237;
  assign n3392 = \[8000]  & n3266;
  assign n3393 = ppeaka_8_8_ & n3191;
  assign n3394_1 = ~n3392 & ~n3393;
  assign n3395 = ~n3391 & n3394_1;
  assign n3396 = \[8750]  & n3267;
  assign n3397 = ppeakb_8_8_ & n3175;
  assign n3398_1 = ~n3396 & ~n3397;
  assign n3399 = n3395 & n3398_1;
  assign n3400 = ~n3390_1 & n3399;
  assign n3401 = ppeaka_8_8_ & n3175;
  assign n3402_1 = n3338 & ~n3401;
  assign n3403 = ~n3338 & n3401;
  assign n3404 = ~n3402_1 & ~n3403;
  assign n3405 = ~n3400 & n3404;
  assign n3406 = n3400 & ~n3404;
  assign n3407_1 = ppeaks_7_7_ & ~n3289;
  assign n3408 = \[7055]  & n3237;
  assign n3409 = \[6065]  & n3266;
  assign n3410 = \[9410]  & n3267;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412_1 = ~n3408 & n3411;
  assign n3413 = ppeaka_7_7_ & n3191;
  assign n3414 = ppeakb_7_7_ & n3175;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = n3412_1 & n3415;
  assign n3417_1 = ~n3407_1 & n3416;
  assign n3418 = ppeaks_6_6_ & ~n3289;
  assign n3419 = \[7685]  & n3237;
  assign n3420 = ppeaka_6_6_ & n3191;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422_1 = \[6740]  & n3266;
  assign n3423 = \[7475]  & n3267;
  assign n3424 = ~n3422_1 & ~n3423;
  assign n3425 = ppeakb_6_6_ & n3175;
  assign n3426 = n3424 & ~n3425;
  assign n3427_1 = n3421 & n3426;
  assign n3428 = ~n3418 & n3427_1;
  assign n3429 = ppeaka_6_6_ & n3175;
  assign n3430 = ~n3333 & n3429;
  assign n3431 = n3335 & ~n3430;
  assign n3432_1 = ~n3428 & n3431;
  assign n3433 = n3428 & ~n3431;
  assign n3434 = ppeaks_5_5_ & ~n3289;
  assign n3435 = ppeaka_5_5_ & n3191;
  assign n3436 = \[4670]  & n3266;
  assign n3437_1 = \[8330]  & n3237;
  assign n3438 = ~n3436 & ~n3437_1;
  assign n3439 = ~n3435 & n3438;
  assign n3440 = \[8105]  & n3267;
  assign n3441 = ppeakb_5_5_ & n3175;
  assign n3442_1 = ~n3440 & ~n3441;
  assign n3443 = n3439 & n3442_1;
  assign n3444 = ~n3434 & n3443;
  assign n3445 = ppeaka_5_5_ & n3175;
  assign n3446 = ~n3332 & ~n3445;
  assign n3447_1 = n3332 & n3445;
  assign n3448 = ~n3446 & ~n3447_1;
  assign n3449 = ~n3444 & ~n3448;
  assign n3450 = n3444 & n3448;
  assign n3451 = ~n3329 & n3331_1;
  assign n3452_1 = ~n3332 & ~n3451;
  assign n3453 = ppeaks_3_3_ & ~n3289;
  assign n3454 = \[15860]  & n3237;
  assign n3455 = \[9995]  & n3266;
  assign n3456 = \[6845]  & n3267;
  assign n3457_1 = ~n3455 & ~n3456;
  assign n3458 = ~n3454 & n3457_1;
  assign n3459 = ppeaka_3_3_ & n3191;
  assign n3460 = ppeakb_3_3_ & n3175;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462_1 = n3458 & n3461;
  assign n3463 = ~n3453 & n3462_1;
  assign n3464 = n3292 & ~n3305;
  assign n3465 = ~n3306_1 & ~n3464;
  assign n3466 = ~n3327 & n3465;
  assign n3467_1 = ppeaka_2_2_ & n3175;
  assign n3468 = n3466 & ~n3467_1;
  assign n3469 = ~n3327 & n3467_1;
  assign n3470 = n3327 & ~n3467_1;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472_1 = ~n3466 & ~n3471;
  assign n3473 = ppeaks_2_2_ & ~n3289;
  assign n3474 = ppeaka_2_2_ & n3191;
  assign n3475 = ppeakb_2_2_ & n3175;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477_1 = \[15515]  & n3237;
  assign n3478 = \[9725]  & n3266;
  assign n3479 = \[4760]  & n3267;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = ~n3477_1 & n3480;
  assign n3482_1 = n3476 & n3481;
  assign n3483 = ~n3473 & n3482_1;
  assign n3484 = ~n3472_1 & ~n3483;
  assign n3485 = ~n3468 & ~n3484;
  assign n3486 = ~n3463 & ~n3485;
  assign n3487_1 = n3463 & n3485;
  assign n3488 = ppeaka_3_3_ & n3175;
  assign n3489 = ~n3328 & n3488;
  assign n3490 = n3330 & ~n3489;
  assign n3491 = ~n3487_1 & n3490;
  assign n3492_1 = ~n3486 & ~n3491;
  assign n3493 = n3452_1 & ~n3492_1;
  assign n3494 = ~n3452_1 & n3492_1;
  assign n3495 = ppeaks_4_4_ & ~n3289;
  assign n3496 = \[14765]  & n3237;
  assign n3497_1 = ppeakb_4_4_ & n3175;
  assign n3498 = \[5375]  & n3266;
  assign n3499 = ~n3497_1 & ~n3498;
  assign n3500 = ~n3496 & n3499;
  assign n3501 = ppeaka_4_4_ & n3191;
  assign n3502_1 = \[6170]  & n3267;
  assign n3503 = ~n3501 & ~n3502_1;
  assign n3504 = n3500 & n3503;
  assign n3505 = ~n3495 & n3504;
  assign n3506 = ~n3494 & ~n3505;
  assign n3507_1 = ~n3493 & ~n3506;
  assign n3508 = ~n3450 & ~n3507_1;
  assign n3509 = ~n3449 & ~n3508;
  assign n3510 = ~n3433 & ~n3509;
  assign n3511 = ~n3432_1 & ~n3510;
  assign n3512_1 = ~n3417_1 & ~n3511;
  assign n3513 = n3417_1 & n3511;
  assign n3514 = ~n3334 & n3337;
  assign n3515 = ~n3338 & ~n3514;
  assign n3516 = ~n3513 & n3515;
  assign n3517_1 = ~n3512_1 & ~n3516;
  assign n3518 = ~n3406 & ~n3517_1;
  assign n3519 = ~n3405 & ~n3518;
  assign n3520 = ~n3389 & ~n3519;
  assign n3521_1 = ~n3388 & ~n3520;
  assign n3522 = n3372 & ~n3521_1;
  assign n3523 = ~n3372 & n3521_1;
  assign n3524 = ppeaks_10_10_ & ~n3289;
  assign n3525_1 = \[5015]  & n3237;
  assign n3526 = ppeaka_10_10_ & n3191;
  assign n3527 = ~n3525_1 & ~n3526;
  assign n3528 = \[9305]  & n3266;
  assign n3529_1 = \[9770]  & n3267;
  assign n3530 = ~n3528 & ~n3529_1;
  assign n3531 = ppeakb_10_10_ & n3175;
  assign n3532 = n3530 & ~n3531;
  assign n3533 = n3527 & n3532;
  assign n3534_1 = ~n3524 & n3533;
  assign n3535 = ~n3523 & ~n3534_1;
  assign n3536 = ~n3522 & ~n3535;
  assign n3537 = ~n3370 & ~n3536;
  assign n3538_1 = ~n3369 & ~n3537;
  assign n3539 = n3353 & ~n3538_1;
  assign n3540 = ~n3353 & n3538_1;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542_1 = n4161 & n3541;
  assign n3543 = \[4640]  & n3312;
  assign n404 = n3542_1 | n3543;
  assign n3545 = ~\[4655]  & ~n3265;
  assign n3546 = ~n3369 & ~n3370;
  assign n3547_1 = ~n3536 & ~n3546;
  assign n3548 = n3536 & n3546;
  assign n3549 = ~n3547_1 & ~n3548;
  assign n3550 = n3265 & n3549;
  assign n3551 = ~preset & ~n3550;
  assign n409 = ~n3545 & n3551;
  assign n3553 = ~n3449 & ~n3450;
  assign n3554 = n3507_1 & ~n3553;
  assign n3555 = ~n3507_1 & n3553;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557_1 = n3192 & n3556;
  assign n3558 = \[4670]  & n3194_1;
  assign n414 = n3557_1 | n3558;
  assign n3560 = ~\[4700]  & ~n3266;
  assign n3561 = ~n3522 & ~n3523;
  assign n3562_1 = n3534_1 & ~n3561;
  assign n3563 = ~n3534_1 & n3561;
  assign n3564 = ~n3562_1 & ~n3563;
  assign n3565 = n3266 & ~n3564;
  assign n3566 = ~preset & ~n3565;
  assign n419 = ~n3560 & n3566;
  assign n3568 = ~preset & n3273;
  assign n3569 = ~n3493 & ~n3494;
  assign n3570 = n3505 & ~n3569;
  assign n3571 = ~n3505 & n3569;
  assign n3572_1 = ~n3570 & ~n3571;
  assign n3573 = n3568 & n3572_1;
  assign n3574 = ~preset & ~n3273;
  assign n3575 = \[4715]  & n3574;
  assign n424 = n3573 | n3575;
  assign n3577_1 = \[4730]  & n3574;
  assign n3578 = ppeaks_15_15_ & ~n3289;
  assign n3579 = \[13550]  & n3237;
  assign n3580 = \[6755]  & n3266;
  assign n3581 = ppeaka_15_15_ & n3191;
  assign n3582_1 = ~n3580 & ~n3581;
  assign n3583 = ~n3579 & n3582_1;
  assign n3584 = \[8765]  & n3267;
  assign n3585 = ppeakb_15_15_ & n3175;
  assign n3586 = ~n3584 & ~n3585;
  assign n3587_1 = n3583 & n3586;
  assign n3588 = ~n3578 & n3587_1;
  assign n3589 = n3336_1 & ~n3347;
  assign n3590 = ~n3340 & n3589;
  assign n3591 = ppeaka_13_13_ & n3175;
  assign n3592_1 = ~n3348 & ~n3591;
  assign n3593 = ~ppeaka_14_14_ & ~n3592_1;
  assign n3594 = ~n3590 & ~n3593;
  assign n3595 = ppeaka_15_15_ & ~ppeaka_14_14_;
  assign n3596 = n3594 & n3595;
  assign n3597_1 = ~ppeaka_15_15_ & ppeaka_14_14_;
  assign n3598 = ~n3596 & ~n3597_1;
  assign n3599 = n3175 & ~n3598;
  assign n3600 = ~ppeaka_15_15_ & ~n3592_1;
  assign n3601 = ~n3590 & ~n3600;
  assign n3602_1 = ~n3599 & n3601;
  assign n3603 = n3588 & ~n3602_1;
  assign n3604 = ~n3588 & n3602_1;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~ppeaka_13_13_ & n3175;
  assign n3607_1 = n3347 & n3606;
  assign n3608 = ppeaka_14_14_ & n3607_1;
  assign n3609 = n3594 & ~n3608;
  assign n3610 = ppeaks_14_14_ & ~n3289;
  assign n3611 = \[15140]  & n3237;
  assign n3612_1 = ppeaka_14_14_ & n3191;
  assign n3613 = ~n3611 & ~n3612_1;
  assign n3614 = \[6080]  & n3266;
  assign n3615 = \[5480]  & n3267;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617_1 = ppeakb_14_14_ & n3175;
  assign n3618 = n3616 & ~n3617_1;
  assign n3619 = n3613 & n3618;
  assign n3620 = ~n3610 & n3619;
  assign n3621 = n3609 & n3620;
  assign n3622_1 = ~n3609 & ~n3620;
  assign n3623 = ~n3347 & n3591;
  assign n3624 = ~n3592_1 & ~n3623;
  assign n3625 = ~n3352 & ~n3538_1;
  assign n3626 = ~n3351_1 & ~n3625;
  assign n3627_1 = ~n3624 & n3626;
  assign n3628 = n3624 & ~n3626;
  assign n3629 = ppeaks_13_13_ & ~n3289;
  assign n3630 = \[15500]  & n3237;
  assign n3631 = ppeaka_13_13_ & n3191;
  assign n3632_1 = ~n3630 & ~n3631;
  assign n3633 = \[4775]  & n3267;
  assign n3634 = \[9740]  & n3266;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636_1 = ppeakb_13_13_ & n3175;
  assign n3637 = n3635 & ~n3636_1;
  assign n3638 = n3632_1 & n3637;
  assign n3639 = ~n3629 & n3638;
  assign n3640_1 = ~n3628 & n3639;
  assign n3641 = ~n3627_1 & ~n3640_1;
  assign n3642 = ~n3622_1 & ~n3641;
  assign n3643 = ~n3621 & ~n3642;
  assign n3644_1 = n3605 & n3643;
  assign n3645 = ~n3605 & ~n3643;
  assign n3646 = ~n3644_1 & ~n3645;
  assign n3647 = n3568 & ~n3646;
  assign n429 = n3577_1 | n3647;
  assign n3649_1 = ~\[4745]  & ~n3218;
  assign n3650 = ~n3388 & ~n3389;
  assign n3651 = n3519 & ~n3650;
  assign n3652 = ~n3519 & n3650;
  assign n3653_1 = ~n3651 & ~n3652;
  assign n3654 = n3218 & ~n3653_1;
  assign n3655 = ~preset & ~n3654;
  assign n434 = ~n3649_1 & n3655;
  assign n3657_1 = ~n3468 & ~n3472_1;
  assign n3658 = n3483 & ~n3657_1;
  assign n3659 = ~n3468 & n3484;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = n3238 & n3660;
  assign n3662_1 = \[4760]  & n3240;
  assign n439 = n3661 | n3662_1;
  assign n3664 = ~n3627_1 & ~n3628;
  assign n3665 = n3639 & n3664;
  assign n3666 = ~n3639 & ~n3664;
  assign n3667_1 = ~n3665 & ~n3666;
  assign n3668 = n3238 & ~n3667_1;
  assign n3669 = \[4775]  & n3240;
  assign n444 = n3668 | n3669;
  assign n3671 = ~preset & n3267;
  assign n3672_1 = ~n3512_1 & ~n3513;
  assign n3673 = ~n3515 & ~n3672_1;
  assign n3674 = n3515 & n3672_1;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = n3671 & n3675;
  assign n3677_1 = ~preset & ~n3267;
  assign n3678 = \[4790]  & n3677_1;
  assign n449 = n3676 | n3678;
  assign n3680 = ~preset & n3275;
  assign n3681 = ~n3310 & n3680;
  assign n3682_1 = ~preset & ~n3275;
  assign n3683 = \[4805]  & n3682_1;
  assign n454 = n3681 | n3683;
  assign n3685 = n3541 & n3680;
  assign n3686 = \[4820]  & n3682_1;
  assign n459 = n3685 | n3686;
  assign n3688 = ~pdn & ~n2923;
  assign n3689 = ~\[18467]  & ~n2930_1;
  assign n3690 = n3688 & n3689;
  assign n3691 = ~\[17817]  & n3690;
  assign n3692_1 = ~\[4835]  & ~n3691;
  assign n3693 = n2880 & n3023_1;
  assign n3694 = ~\[17206]  & n3693;
  assign n3695 = n2880 & n3046_1;
  assign n3696 = ~\[17180]  & n3695;
  assign n3697_1 = n2880 & n2949;
  assign n3698 = ~\[17115]  & n3697_1;
  assign n3699 = ~n3696 & ~n3698;
  assign n3700 = ~n3694 & n3699;
  assign n3701 = n2880 & n3020;
  assign n3702_1 = ~\[18025]  & n3701;
  assign n3703 = ~n3691 & ~n3702_1;
  assign n3704 = n3700 & n3703;
  assign n3705 = ppeaks_6_6_ & ~n3704;
  assign n3706 = ~\[17037]  & \[18025] ;
  assign n3707_1 = \[17635]  & ~\[17986] ;
  assign n3708 = n2930_1 & n3707_1;
  assign n3709 = ~n3706 & ~n3708;
  assign n3710 = ppeakp_6_6_ & ~n3709;
  assign n3711 = n2880 & n3044;
  assign n3712_1 = ~\[17245]  & n3711;
  assign n3713 = ppeaka_6_6_ & n3712_1;
  assign n3714 = ~n3710 & ~n3713;
  assign n3715 = \[9950]  & ~n2930_1;
  assign n3716 = n3707_1 & n3715;
  assign n3717_1 = \[17427]  & ~\[17648] ;
  assign n3718 = \[4835]  & n3717_1;
  assign n3719 = ~n3716 & ~n3718;
  assign n3720 = ~\[17999]  & \[18077] ;
  assign n3721 = \[14210]  & n3720;
  assign n3722_1 = n3719 & ~n3721;
  assign n3723 = n3714 & n3722_1;
  assign n3724 = \[17180]  & ~\[17232] ;
  assign n3725 = \[7625]  & n3724;
  assign n3726 = ppeakb_6_6_ & n3275;
  assign n3727_1 = ~n3725 & ~n3726;
  assign n3728 = n3723 & n3727_1;
  assign n3729 = ~n3705 & n3728;
  assign n3730 = ppeaka_6_6_ & n3275;
  assign n3731 = ppeaks_5_5_ & ~n3704;
  assign n3732_1 = ppeakp_5_5_ & ~n3709;
  assign n3733 = ppeaka_5_5_ & n3712_1;
  assign n3734 = ~n3732_1 & ~n3733;
  assign n3735 = \[10220]  & ~n2930_1;
  assign n3736 = n3707_1 & n3735;
  assign n3737_1 = \[15395]  & n3720;
  assign n3738 = ~n3736 & ~n3737_1;
  assign n3739 = \[6905]  & n3717_1;
  assign n3740 = n3738 & ~n3739;
  assign n3741 = n3734 & n3740;
  assign n3742_1 = \[6995]  & n3724;
  assign n3743 = ppeakb_5_5_ & n3275;
  assign n3744 = ~n3742_1 & ~n3743;
  assign n3745 = n3741 & n3744;
  assign n3746 = ~n3731 & n3745;
  assign n3747_1 = ppeaks_4_4_ & ~n3704;
  assign n3748 = ppeakb_4_4_ & n3275;
  assign n3749 = \[6230]  & n3717_1;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751_1 = ppeaka_4_4_ & n3712_1;
  assign n3752 = \[12245]  & n3724;
  assign n3753 = ~n3751_1 & ~n3752;
  assign n3754 = n3750 & n3753;
  assign n3755_1 = ppeakp_4_4_ & ~n3709;
  assign n3756 = \[10505]  & ~n2930_1;
  assign n3757 = n3707_1 & n3756;
  assign n3758 = ~n3755_1 & ~n3757;
  assign n3759_1 = \[15035]  & n3720;
  assign n3760 = n3758 & ~n3759_1;
  assign n3761 = n3754 & n3760;
  assign n3762 = ~n3747_1 & n3761;
  assign n3763 = ppeaks_3_3_ & ~n3704;
  assign n3764_1 = ppeakb_3_3_ & n3275;
  assign n3765 = \[10790]  & ~n2930_1;
  assign n3766 = n3707_1 & n3765;
  assign n3767 = \[12455]  & n3724;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769_1 = ~n3764_1 & n3768;
  assign n3770 = ppeaka_3_3_ & n3712_1;
  assign n3771 = ppeakp_3_3_ & ~n3709;
  assign n3772 = \[12845]  & n3720;
  assign n3773_1 = \[8165]  & n3717_1;
  assign n3774 = ~n3772 & ~n3773_1;
  assign n3775 = ~n3771 & n3774;
  assign n3776 = ~n3770 & n3775;
  assign n3777 = n3769_1 & n3776;
  assign n3778_1 = ~n3763 & n3777;
  assign n3779 = ppeaks_2_2_ & ~n3704;
  assign n3780 = ppeaka_2_2_ & n3712_1;
  assign n3781 = ppeakp_2_2_ & ~n3709;
  assign n3782 = ppeakb_2_2_ & n3275;
  assign n3783_1 = ~n3781 & ~n3782;
  assign n3784 = ~n3780 & n3783_1;
  assign n3785 = \[11060]  & ~n2930_1;
  assign n3786 = n3707_1 & n3785;
  assign n3787 = \[7535]  & n3717_1;
  assign n3788_1 = \[13100]  & n3720;
  assign n3789 = ~n3787 & ~n3788_1;
  assign n3790 = ~n3786 & n3789;
  assign n3791 = \[12680]  & n3724;
  assign n3792 = n3790 & ~n3791;
  assign n3793_1 = n3784 & n3792;
  assign n3794 = ~n3779 & n3793_1;
  assign n3795 = ppeaks_1_1_ & ~n3704;
  assign n3796 = ppeakp_1_1_ & ~n3709;
  assign n3797 = ppeakb_1_1_ & n3275;
  assign n3798_1 = ~n3796 & ~n3797;
  assign n3799 = \[11315]  & ~n2930_1;
  assign n3800 = n3707_1 & n3799;
  assign n3801 = \[12920]  & n3724;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803_1 = \[9485]  & n3717_1;
  assign n3804 = n3802 & ~n3803_1;
  assign n3805 = n3798_1 & n3804;
  assign n3806 = \[12380]  & n3720;
  assign n3807 = ppeaka_1_1_ & n3712_1;
  assign n3808_1 = ~n3806 & ~n3807;
  assign n3809 = n3805 & n3808_1;
  assign n3810 = ~n3795 & n3809;
  assign n3811 = ppeakb_0_0_ & n3275;
  assign n3812 = \[13175]  & n3724;
  assign n3813_1 = \[12605]  & n3720;
  assign n3814 = ~n3812 & ~n3813_1;
  assign n3815 = ~n3811 & n3814;
  assign n3816 = ppeaka_0_0_ & n3712_1;
  assign n3817 = \[11555]  & ~n2930_1;
  assign n3818_1 = n3707_1 & n3817;
  assign n3819 = ppeakp_0_0_ & ~n3709;
  assign n3820 = \[11630]  & n3717_1;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = ~n3818_1 & n3821;
  assign n3823_1 = ~n3816 & n3822;
  assign n3824 = n3815 & n3823_1;
  assign n3825 = ~n3706 & ~n3717_1;
  assign n3826 = ~n3707_1 & n3825;
  assign n3827 = ~n3720 & n3826;
  assign n3828_1 = ppeaka_0_0_ & n3275;
  assign n3829 = ~n3712_1 & ~n3828_1;
  assign n3830 = n3827 & n3829;
  assign n3831 = n3704 & n3830;
  assign n3832 = ~n3824 & ~n3831;
  assign n3833_1 = ppeaks_0_0_ & ~n3704;
  assign n3834 = ~n3832 & ~n3833_1;
  assign n3835 = ~n3810 & ~n3834;
  assign n3836 = n3810 & n3834;
  assign n3837 = ppeaka_1_1_ & n3275;
  assign n3838_1 = ~n3724 & ~n3837;
  assign n3839 = ~n3836 & ~n3838_1;
  assign n3840 = ~n3835 & ~n3839;
  assign n3841 = n3794 & n3840;
  assign n3842 = ~n3794 & ~n3840;
  assign n3843_1 = ppeaka_2_2_ & n3275;
  assign n3844 = ~n3842 & ~n3843_1;
  assign n3845 = ~n3841 & ~n3844;
  assign n3846 = ~n3778_1 & n3845;
  assign n3847 = n3778_1 & ~n3845;
  assign n3848_1 = ppeaka_3_3_ & n3275;
  assign n3849 = ~n3847 & n3848_1;
  assign n3850 = ~n3846 & ~n3849;
  assign n3851 = ~n3762 & ~n3850;
  assign n3852 = n3762 & n3850;
  assign n3853_1 = ppeaka_4_4_ & n3275;
  assign n3854 = ~n3852 & n3853_1;
  assign n3855 = ~n3851 & ~n3854;
  assign n3856 = ~n3746 & ~n3855;
  assign n3857_1 = n3746 & n3855;
  assign n3858 = ppeaka_5_5_ & n3275;
  assign n3859 = ~n3857_1 & n3858;
  assign n3860 = ~n3856 & ~n3859;
  assign n3861_1 = n3730 & ~n3860;
  assign n3862 = ~n3730 & n3860;
  assign n3863 = ~n3861_1 & ~n3862;
  assign n3864 = n3729 & n3863;
  assign n3865_1 = ~n3729 & ~n3863;
  assign n3866 = ~n3864 & ~n3865_1;
  assign n3867 = n3691 & n3866;
  assign n3868 = ~preset & ~n3867;
  assign n464 = ~n3692_1 & n3868;
  assign n3870_1 = ~\[4850]  & ~n3707_1;
  assign n3871 = ppeaks_10_10_ & ~n3704;
  assign n3872 = ppeakb_10_10_ & n3275;
  assign n3873 = \[11795]  & ~n2930_1;
  assign n3874 = n3707_1 & n3873;
  assign n3875_1 = \[9860]  & n3724;
  assign n3876 = ~n3874 & ~n3875_1;
  assign n3877 = ~n3872 & n3876;
  assign n3878 = \[10925]  & n3717_1;
  assign n3879_1 = ppeaka_10_10_ & n3712_1;
  assign n3880 = ppeakp_10_10_ & ~n3709;
  assign n3881 = \[12860]  & n3720;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = ~n3879_1 & n3882;
  assign n3884_1 = ~n3878 & n3883;
  assign n3885 = n3877 & n3884_1;
  assign n3886 = ~n3871 & n3885;
  assign n3887 = ppeaka_10_10_ & n3275;
  assign n3888 = ppeaks_9_9_ & ~n3704;
  assign n3889_1 = ppeakb_9_9_ & n3275;
  assign n3890 = ppeaka_9_9_ & n3712_1;
  assign n3891 = ~n3889_1 & ~n3890;
  assign n3892 = ppeakp_9_9_ & ~n3709;
  assign n3893 = \[13820]  & n3720;
  assign n3894_1 = \[9590]  & n3724;
  assign n3895 = ~n3893 & ~n3894_1;
  assign n3896 = \[11570]  & ~n2930_1;
  assign n3897 = n3707_1 & n3896;
  assign n3898 = \[11645]  & n3717_1;
  assign n3899_1 = ~n3897 & ~n3898;
  assign n3900 = n3895 & n3899_1;
  assign n3901 = ~n3892 & n3900;
  assign n3902 = n3891 & n3901;
  assign n3903 = ~n3888 & n3902;
  assign n3904_1 = ppeaks_8_8_ & ~n3704;
  assign n3905 = ppeakp_8_8_ & ~n3709;
  assign n3906 = ppeaka_8_8_ & n3712_1;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = \[11330]  & ~n2930_1;
  assign n3909_1 = n3707_1 & n3908;
  assign n3910 = \[13460]  & n3720;
  assign n3911 = ~n3909_1 & ~n3910;
  assign n3912 = \[8915]  & n3724;
  assign n3913 = n3911 & ~n3912;
  assign n3914_1 = n3907 & n3913;
  assign n3915 = \[11420]  & n3717_1;
  assign n3916 = ppeakb_8_8_ & n3275;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = n3914_1 & n3917;
  assign n3919_1 = ~n3904_1 & n3918;
  assign n3920 = ppeaks_7_7_ & ~n3704;
  assign n3921 = ppeakb_7_7_ & n3275;
  assign n3922 = \[11075]  & ~n2930_1;
  assign n3923 = n3707_1 & n3922;
  assign n3924_1 = \[5540]  & n3717_1;
  assign n3925 = ~n3923 & ~n3924_1;
  assign n3926 = ~n3921 & n3925;
  assign n3927 = ppeaka_7_7_ & n3712_1;
  assign n3928 = ppeakp_7_7_ & ~n3709;
  assign n3929_1 = \[14630]  & n3720;
  assign n3930 = \[8255]  & n3724;
  assign n3931 = ~n3929_1 & ~n3930;
  assign n3932 = ~n3928 & n3931;
  assign n3933 = ~n3927 & n3932;
  assign n3934_1 = n3926 & n3933;
  assign n3935 = ~n3920 & n3934_1;
  assign n3936 = ~n3729 & ~n3862;
  assign n3937 = ~n3861_1 & ~n3936;
  assign n3938 = ~n3935 & ~n3937;
  assign n3939_1 = n3935 & n3937;
  assign n3940 = ppeaka_7_7_ & n3275;
  assign n3941 = ~n3939_1 & n3940;
  assign n3942 = ~n3938 & ~n3941;
  assign n3943 = ~n3919_1 & ~n3942;
  assign n3944_1 = n3919_1 & n3942;
  assign n3945 = ppeaka_8_8_ & n3275;
  assign n3946 = ~n3944_1 & n3945;
  assign n3947 = ~n3943 & ~n3946;
  assign n3948 = ~n3903 & ~n3947;
  assign n3949_1 = n3903 & n3947;
  assign n3950 = ppeaka_9_9_ & n3275;
  assign n3951 = ~n3949_1 & n3950;
  assign n3952 = ~n3948 & ~n3951;
  assign n3953 = ~n3887 & n3952;
  assign n3954_1 = n3887 & ~n3952;
  assign n3955 = ~n3953 & ~n3954_1;
  assign n3956 = n3886 & n3955;
  assign n3957 = ~n3886 & ~n3955;
  assign n3958_1 = ~n3956 & ~n3957;
  assign n3959 = n3707_1 & n3958_1;
  assign n3960 = ~preset & ~n3959;
  assign n469 = ~n3870_1 & n3960;
  assign n3962 = ~preset & n3702_1;
  assign n3963_1 = ~n3851 & ~n3852;
  assign n3964 = ~n3853_1 & ~n3963_1;
  assign n3965 = n3853_1 & n3963_1;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = n3962 & n3966;
  assign n3968_1 = ~preset & ~n3702_1;
  assign n3969 = \[4865]  & n3968_1;
  assign n474 = n3967 | n3969;
  assign n3971 = \[4880]  & n3968_1;
  assign n3972 = ppeaka_15_15_ & n3275;
  assign n3973_1 = ppeaks_15_15_ & ~n3704;
  assign n3974 = ppeakb_15_15_ & n3275;
  assign n3975 = \[12470]  & ~n2930_1;
  assign n3976 = n3707_1 & n3975;
  assign n3977_1 = \[6320]  & n3724;
  assign n3978 = ~n3976 & ~n3977_1;
  assign n3979 = ~n3974 & n3978;
  assign n3980 = \[14615]  & n3717_1;
  assign n3981 = ppeaka_15_15_ & n3712_1;
  assign n3982_1 = ppeakp_15_15_ & ~n3709;
  assign n3983 = \[15050]  & n3720;
  assign n3984 = ~n3982_1 & ~n3983;
  assign n3985 = ~n3981 & n3984;
  assign n3986 = ~n3980 & n3985;
  assign n3987_1 = n3979 & n3986;
  assign n3988 = ~n3973_1 & n3987_1;
  assign n3989 = n3972 & ~n3988;
  assign n3990 = ~n3972 & n3988;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992_1 = ppeaks_14_14_ & ~n3704;
  assign n3993 = ppeaka_14_14_ & n3712_1;
  assign n3994 = \[10985]  & n3724;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ppeakb_14_14_ & n3275;
  assign n3997_1 = \[15410]  & n3720;
  assign n3998 = ~n3996 & ~n3997_1;
  assign n3999 = n3995 & n3998;
  assign n4000 = ppeakp_14_14_ & ~n3709;
  assign n4001 = \[12260]  & ~n2930_1;
  assign n4002_1 = n3707_1 & n4001;
  assign n4003 = ~n4000 & ~n4002_1;
  assign n4004 = \[13445]  & n3717_1;
  assign n4005 = n4003 & ~n4004;
  assign n4006 = n3999 & n4005;
  assign n4007_1 = ~n3992_1 & n4006;
  assign n4008 = ppeaks_13_13_ & ~n3704;
  assign n4009 = ppeakb_13_13_ & n3275;
  assign n4010 = \[12170]  & ~n2930_1;
  assign n4011 = n3707_1 & n4010;
  assign n4012_1 = \[10700]  & n3724;
  assign n4013 = ~n4011 & ~n4012_1;
  assign n4014 = ~n4009 & n4013;
  assign n4015 = \[13805]  & n3717_1;
  assign n4016 = ppeaka_13_13_ & n3712_1;
  assign n4017_1 = ppeakp_13_13_ & ~n3709;
  assign n4018 = \[12620]  & n3720;
  assign n4019 = ~n4017_1 & ~n4018;
  assign n4020 = ~n4016 & n4019;
  assign n4021 = ~n4015 & n4020;
  assign n4022_1 = n4014 & n4021;
  assign n4023 = ~n4008 & n4022_1;
  assign n4024 = ppeaks_12_12_ & ~n3704;
  assign n4025 = \[10415]  & n3724;
  assign n4026 = \[12395]  & n3720;
  assign n4027_1 = ~n4025 & ~n4026;
  assign n4028 = \[15755]  & n3717_1;
  assign n4029 = n4027_1 & ~n4028;
  assign n4030 = ~n4024 & n4029;
  assign n4031 = ppeaka_12_12_ & n3712_1;
  assign n4032_1 = ppeakb_12_12_ & n3275;
  assign n4033 = ~n4031 & ~n4032_1;
  assign n4034 = ppeakp_12_12_ & ~n3709;
  assign n4035 = \[12050]  & ~n2930_1;
  assign n4036 = n3707_1 & n4035;
  assign n4037_1 = ~n4034 & ~n4036;
  assign n4038 = n4033 & n4037_1;
  assign n4039 = n4030 & n4038;
  assign n4040 = ppeaks_11_11_ & ~n3704;
  assign n4041 = ppeakp_11_11_ & ~n3709;
  assign n4042_1 = ppeakb_11_11_ & n3275;
  assign n4043 = ~n4041 & ~n4042_1;
  assign n4044 = \[11915]  & ~n2930_1;
  assign n4045 = n3707_1 & n4044;
  assign n4046 = \[16100]  & n3717_1;
  assign n4047_1 = ~n4045 & ~n4046;
  assign n4048 = \[10130]  & n3724;
  assign n4049 = n4047_1 & ~n4048;
  assign n4050 = n4043 & n4049;
  assign n4051 = \[13115]  & n3720;
  assign n4052_1 = ppeaka_11_11_ & n3712_1;
  assign n4053 = ~n4051 & ~n4052_1;
  assign n4054 = n4050 & n4053;
  assign n4055 = ~n4040 & n4054;
  assign n4056 = ~n3886 & ~n3953;
  assign n4057_1 = ~n3954_1 & ~n4056;
  assign n4058 = n4055 & n4057_1;
  assign n4059 = ~n4055 & ~n4057_1;
  assign n4060 = ppeaka_11_11_ & n3275;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062_1 = ~n4058 & ~n4061;
  assign n4063 = ~n4039 & n4062_1;
  assign n4064 = n4039 & ~n4062_1;
  assign n4065 = ppeaka_12_12_ & n3275;
  assign n4066 = ~n4064 & n4065;
  assign n4067_1 = ~n4063 & ~n4066;
  assign n4068 = n4023 & n4067_1;
  assign n4069 = ~n4023 & ~n4067_1;
  assign n4070 = ppeaka_13_13_ & n3275;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072_1 = ~n4068 & ~n4071;
  assign n4073 = n4007_1 & ~n4072_1;
  assign n4074 = ~n4007_1 & n4072_1;
  assign n4075 = ppeaka_14_14_ & n3275;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077_1 = ~n4073 & ~n4076;
  assign n4078 = ~n3991 & n4077_1;
  assign n4079 = n3991 & ~n4077_1;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = n3962 & ~n4080;
  assign n479 = n3971 | n4081;
  assign n4083 = ~\[4895]  & ~n3706;
  assign n4084 = ~n3948 & ~n3949_1;
  assign n4085 = ~n3950 & ~n4084;
  assign n4086 = n3950 & n4084;
  assign n4087_1 = ~n4085 & ~n4086;
  assign n4088 = n3706 & ~n4087_1;
  assign n4089 = ~preset & ~n4088;
  assign n484 = ~n4083 & n4089;
  assign n4091 = ~preset & n3694;
  assign n4092_1 = ~n3846 & ~n3847;
  assign n4093 = n3848_1 & n4092_1;
  assign n4094 = ~n3848_1 & ~n4092_1;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = n4091 & n4095;
  assign n4097_1 = ~preset & ~n3694;
  assign n4098 = \[4910]  & n4097_1;
  assign n489 = n4096 | n4098;
  assign n4100 = \[4925]  & n3682_1;
  assign n4101 = ~n3835 & ~n3836;
  assign n4102_1 = n3838_1 & ~n4101;
  assign n4103 = ~n3838_1 & n4101;
  assign n4104 = ~n4102_1 & ~n4103;
  assign n4105 = n3680 & n4104;
  assign n494 = n4100 | n4105;
  assign n4107_1 = \[4940]  & n3682_1;
  assign n4108 = ~n4063 & ~n4064;
  assign n4109 = ~n4065 & ~n4108;
  assign n4110 = n4065 & n4108;
  assign n4111 = ~n4109 & ~n4110;
  assign n4112_1 = n3680 & n4111;
  assign n499 = n4107_1 | n4112_1;
  assign n4114 = ~preset & n3712_1;
  assign n4115 = ~n3866 & n4114;
  assign n4116 = ~preset & ~n3712_1;
  assign n4117_1 = \[4955]  & n4116;
  assign n504 = n4115 | n4117_1;
  assign n4119 = ~\[4970]  & ~n2843;
  assign n4120 = ~pdata_1_1_ & n2843;
  assign n4121 = ~preset & ~n4120;
  assign n509 = ~n4119 & n4121;
  assign n4123 = ppeakb_0_0_ & ~n2989;
  assign n4124 = n2907_1 & ~n2950_1;
  assign n4125 = ppeaka_0_0_ & n4124;
  assign n4126 = ~n4123 & ~n4125;
  assign n4127_1 = \[4355]  & n2912_1;
  assign n4128 = \[4310]  & n2931;
  assign n4129 = \[8405]  & n2936;
  assign n4130 = \[15995]  & n2939;
  assign n4131 = \[4580]  & n2916_1;
  assign n4132_1 = ~n4130 & ~n4131;
  assign n4133 = \[15605]  & n2961;
  assign n4134 = \[10550]  & n2964;
  assign n4135 = ~n4133 & ~n4134;
  assign n4136 = \[5900]  & n2959;
  assign n4137_1 = \[7835]  & n2955_1;
  assign n4138 = ~n4136 & ~n4137_1;
  assign n4139 = n4135 & n4138;
  assign n4140 = n4132_1 & n4139;
  assign n4141 = n2907_1 & ~n4140;
  assign n4142_1 = ~n4129 & ~n4141;
  assign n4143 = ~n4128 & n4142_1;
  assign n4144 = ~n4127_1 & n4143;
  assign n4145 = ~n2906 & ~n4144;
  assign n4146 = \[13655]  & n3081_1;
  assign n4147_1 = ~n4145 & ~n4146;
  assign n514 = ~n4126 | ~n4147_1;
  assign n4149 = \[10970]  & n3024;
  assign n4150 = ppeakp_7_7_ & ~n3035;
  assign n4151_1 = ppeaka_7_7_ & ppeakb_7_7_;
  assign n4152 = n2912_1 & ~n4151_1;
  assign n4153 = \[12335]  & n2936;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = ~n4150 & n4154;
  assign n4156_1 = ~n4149 & n4155;
  assign n4157 = ~n2906 & ~n4156_1;
  assign n4158 = ppeaka_8_8_ & n2975_1;
  assign n4159 = ~n4157 & ~n4158;
  assign n4160 = ppeaka_7_7_ & ~n3042_1;
  assign n4161_1 = \[7025]  & n3044;
  assign n4162 = \[7055]  & ~n3047;
  assign n4163 = \[13985]  & n3020;
  assign n4164 = \[5180]  & n3030;
  assign n4165 = ~n4163 & ~n4164;
  assign n4166_1 = ~n4162 & n4165;
  assign n4167 = ppeakb_7_7_ & ~n3050;
  assign n4168 = \[4430]  & n2961;
  assign n4169 = \[10460]  & n2964;
  assign n4170_1 = ~n4168 & ~n4169;
  assign n4171 = ~n4167 & n4170_1;
  assign n4172 = n4166_1 & n4171;
  assign n4173 = ~n4161_1 & n4172;
  assign n4174 = n2907_1 & ~n4173;
  assign n4175_1 = ~n4160 & ~n4174;
  assign n518 = ~n4159 | ~n4175_1;
  assign n4177 = \[5015]  & ~n3065;
  assign n4178 = \[9620]  & n3068;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180_1 = \[8180]  & n2931;
  assign n4181 = \[9200]  & n2917;
  assign n4182 = ~n4180_1 & ~n4181;
  assign n522 = ~n4179 | ~n4182;
  assign n4184 = \[5030]  & ~n3065;
  assign n4185_1 = \[9185]  & n2917;
  assign n4186 = ~n4184 & ~n4185_1;
  assign n4187 = \[13835]  & n2931;
  assign n4188 = \[9605]  & n3068;
  assign n4189 = ~n4187 & ~n4188;
  assign n527 = ~n4186 | ~n4189;
  assign n4191 = \[12350]  & n3081_1;
  assign n4192 = ppeaks_4_4_ & ~n3090;
  assign n4193 = \[14975]  & n2936;
  assign n4194 = \[11120]  & n2912_1;
  assign n4195_1 = ~n4193 & ~n4194;
  assign n4196 = \[15035]  & n2931;
  assign n4197 = \[5615]  & n3024;
  assign n4198 = \[11765]  & n3095;
  assign n4199 = \[12245]  & n3046_1;
  assign n4200_1 = \[13790]  & n2939;
  assign n4201 = ~n4199 & ~n4200_1;
  assign n4202 = \[9785]  & n2916_1;
  assign n4203 = n4201 & ~n4202;
  assign n4204_1 = \[14675]  & n2949;
  assign n4205 = \[8015]  & n2961;
  assign n4206 = ~n4204_1 & ~n4205;
  assign n4207 = \[4865]  & n3020;
  assign n4208 = n4206 & ~n4207;
  assign n4209_1 = \[4715]  & n2955_1;
  assign n4210 = \[9380]  & n2959;
  assign n4211 = \[6875]  & n2964;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = ~n4209_1 & n4212;
  assign n4214_1 = n4208 & n4213;
  assign n4215 = n4203 & n4214_1;
  assign n4216 = n2907_1 & ~n4215;
  assign n4217 = ~n4198 & ~n4216;
  assign n4218 = ~n4197 & n4217;
  assign n4219_1 = ~n4196 & n4218;
  assign n4220 = n4195_1 & n4219_1;
  assign n4221 = ~n2906 & ~n4220;
  assign n4222 = ~n4192 & ~n4221;
  assign n532 = n4191 | ~n4222;
  assign n4224_1 = ppeakp_11_11_ & ~n3147;
  assign n4225 = \[5555]  & ~n2927;
  assign n4226 = \[12020]  & n3095;
  assign n4227 = ppeakb_11_11_ & n2917;
  assign n4228_1 = ~n4226 & ~n4227;
  assign n4229 = ~n4225 & n4228_1;
  assign n4230 = ppeaka_11_11_ & ~n3156;
  assign n4231 = \[6290]  & n3021;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233_1 = n4229 & n4232;
  assign n536 = n4224_1 | ~n4233_1;
  assign n4235 = ~\[5075]  & ~n3162;
  assign n4236 = ~pdata_1_1_ & n3162;
  assign n4237 = ~preset & ~n4236;
  assign n540 = ~n4235 & n4237;
  assign n4239 = ~\[5090]  & ~n3162;
  assign n4240 = ~pdata_10_10_ & n3162;
  assign n4241 = ~preset & ~n4240;
  assign n545 = ~n4239 & n4241;
  assign n4243_1 = ~\[5105]  & ~n3181;
  assign n4244 = ~pdata_2_2_ & n3181;
  assign n4245 = ~preset & ~n4244;
  assign n550 = ~n4243_1 & n4245;
  assign n4247 = ~\[5120]  & ~n3181;
  assign n4248_1 = ~pdata_11_11_ & n3181;
  assign n4249 = ~preset & ~n4248_1;
  assign n555 = ~n4247 & n4249;
  assign n4251 = pdata_8_8_ & n3192;
  assign n4252_1 = \[5135]  & n3194_1;
  assign n560 = n4251 | n4252_1;
  assign n4254 = pdata_1_1_ & n3192;
  assign n4255 = \[5150]  & n3194_1;
  assign n565 = n4254 | n4255;
  assign n4257_1 = pdata_14_14_ & n3192;
  assign n4258 = \[5165]  & n3194_1;
  assign n570 = n4257_1 | n4258;
  assign n4260 = ~\[5180]  & ~n3203;
  assign n4261 = ~pdata_7_7_ & n3203;
  assign n4262_1 = ~preset & ~n4261;
  assign n575 = ~n4260 & n4262_1;
  assign n4264 = ~pdata_4_4_ & n3208;
  assign n4265 = ~\[5195]  & ~n3208;
  assign n4266_1 = ~preset & ~n4265;
  assign n580 = ~n4264 & n4266_1;
  assign n4268 = ~pdata_13_13_ & n3208;
  assign n4269 = ~\[5210]  & ~n3208;
  assign n4270 = ~preset & ~n4269;
  assign n585 = ~n4268 & n4270;
  assign n4272 = ~\[5225]  & ~n3218;
  assign n4273 = ~pdata_10_10_ & n3218;
  assign n4274 = ~preset & ~n4273;
  assign n590 = ~n4272 & n4274;
  assign n4276_1 = \[5240]  & n3225;
  assign n4277 = pdata_5_5_ & n3963;
  assign n595 = n4276_1 | n4277;
  assign n4279 = ~\[5255]  & ~n3231;
  assign n4280 = ~pdata_11_11_ & n3231;
  assign n4281_1 = ~preset & ~n4280;
  assign n600 = ~n4279 & n4281_1;
  assign n4283 = pdata_4_4_ & n3238;
  assign n4284 = \[5270]  & n3240;
  assign n605 = n4283 | n4284;
  assign n4286_1 = pdata_1_1_ & n3238;
  assign n4287 = \[5285]  & n3240;
  assign n610 = n4286_1 | n4287;
  assign n4289 = pdata_10_10_ & n3238;
  assign n4290 = \[5300]  & n3240;
  assign n615 = n4289 | n4290;
  assign n4292 = ~\[5315]  & ~n3249_1;
  assign n4293 = ~pdata_7_7_ & n3249_1;
  assign n4294 = ~preset & ~n4293;
  assign n620 = ~n4292 & n4294;
  assign n4296_1 = \[5330]  & n3312;
  assign n4297 = n3278 & ~n3287;
  assign n4298 = ~n3292 & ~n4297;
  assign n4299 = n4161 & ~n4298;
  assign n625 = n4296_1 | n4299;
  assign n4301_1 = n4161 & ~n3667_1;
  assign n4302 = \[5345]  & n3312;
  assign n630 = n4301_1 | n4302;
  assign n4304 = ~\[5360]  & ~n3265;
  assign n4305_1 = n3265 & ~n3541;
  assign n4306 = ~preset & ~n4305_1;
  assign n635 = ~n4304 & n4306;
  assign n4308 = n3192 & n3572_1;
  assign n4309 = \[5375]  & n3194_1;
  assign n640 = n4308 | n4309;
  assign n4311 = ~\[5390]  & ~n3266;
  assign n4312 = n3266 & n4298;
  assign n4313 = ~preset & ~n4312;
  assign n645 = ~n4311 & n4313;
  assign n4315_1 = ~\[5405]  & ~n3266;
  assign n4316 = n3266 & ~n3653_1;
  assign n4317 = ~preset & ~n4316;
  assign n650 = ~n4315_1 & n4317;
  assign n4319 = n3556 & n3568;
  assign n4320_1 = \[5420]  & n3574;
  assign n655 = n4319 | n4320_1;
  assign n4322 = \[5435]  & n3574;
  assign n4323 = ~n3621 & ~n3622_1;
  assign n4324 = n3641 & ~n4323;
  assign n4325_1 = ~n3641 & n4323;
  assign n4326 = ~n4324 & ~n4325_1;
  assign n4327 = n3568 & ~n4326;
  assign n660 = n4322 | n4327;
  assign n4329_1 = ~\[5450]  & ~n3218;
  assign n4330 = n3218 & ~n3564;
  assign n4331 = ~preset & ~n4330;
  assign n665 = ~n4329_1 & n4331;
  assign n4333 = ~\[5465]  & ~n3231;
  assign n4334_1 = n3231 & ~n3653_1;
  assign n4335 = ~preset & ~n4334_1;
  assign n670 = ~n4333 & n4335;
  assign n4337 = n3238 & ~n4326;
  assign n4338 = \[5480]  & n3240;
  assign n675 = n4337 | n4338;
  assign n4340 = \[5495]  & n3677_1;
  assign n4341 = ~n3432_1 & ~n3433;
  assign n4342 = ~n3509 & ~n4341;
  assign n4343 = n3509 & n4341;
  assign n4344_1 = ~n4342 & ~n4343;
  assign n4345 = n3671 & ~n4344_1;
  assign n680 = n4340 | n4345;
  assign n4347 = n3660 & n3680;
  assign n4348 = \[5510]  & n3682_1;
  assign n685 = n4347 | n4348;
  assign n4350 = ~n3549 & n3680;
  assign n4351 = \[5525]  & n3682_1;
  assign n690 = n4350 | n4351;
  assign n4353 = ~\[5540]  & ~n3691;
  assign n4354_1 = ~n3938 & ~n3939_1;
  assign n4355 = ~n3940 & ~n4354_1;
  assign n4356 = n3940 & n4354_1;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = n3691 & ~n4357;
  assign n4359_1 = ~preset & ~n4358;
  assign n695 = ~n4353 & n4359_1;
  assign n4361 = ~\[5555]  & ~n3707_1;
  assign n4362 = ~n4058 & ~n4059;
  assign n4363 = ~n4060 & n4362;
  assign n4364_1 = n4060 & ~n4362;
  assign n4365 = ~n4363 & ~n4364_1;
  assign n4366 = n3707_1 & n4365;
  assign n4367 = ~preset & ~n4366;
  assign n700 = ~n4361 & n4367;
  assign n4369_1 = \[5570]  & n3968_1;
  assign n4370 = n3962 & n4095;
  assign n705 = n4369_1 | n4370;
  assign n4372 = ~\[5600]  & ~n3706;
  assign n4373 = ~n3943 & ~n3944_1;
  assign n4374_1 = ~n3945 & ~n4373;
  assign n4375 = n3945 & n4373;
  assign n4376 = ~n4374_1 & ~n4375;
  assign n4377 = n3706 & ~n4376;
  assign n4378 = ~preset & ~n4377;
  assign n710 = ~n4372 & n4378;
  assign n4380 = n3966 & n4091;
  assign n4381 = \[5615]  & n4097_1;
  assign n715 = n4380 | n4381;
  assign n4082 = ~preset & n3724;
  assign n4384_1 = n4376 & n4082;
  assign n4385 = ~preset & ~n3724;
  assign n4386 = \[5630]  & n4385;
  assign n720 = n4384_1 | n4386;
  assign n4388_1 = \[5645]  & n3682_1;
  assign n4389 = ~n4068 & ~n4069;
  assign n4390 = ~n4070 & n4389;
  assign n4391 = n4070 & ~n4389;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393_1 = n3680 & ~n4392;
  assign n725 = n4388_1 | n4393_1;
  assign n4395 = \[5660]  & n4116;
  assign n4396 = ~n3856 & ~n3857_1;
  assign n4397 = ~n3858 & ~n4396;
  assign n4398_1 = n3858 & n4396;
  assign n4399 = ~n4397 & ~n4398_1;
  assign n4400 = n4114 & n4399;
  assign n730 = n4395 | n4400;
  assign n4402 = ~\[5675]  & ~n2843;
  assign n4403_1 = ~pdata_0_0_ & n2843;
  assign n4404 = ~preset & ~n4403_1;
  assign n735 = ~n4402 & n4404;
  assign n4406 = ppeakb_10_10_ & ~n2989;
  assign n4407 = ppeaka_10_10_ & n4124;
  assign n4408_1 = ~n4406 & ~n4407;
  assign n4409 = \[14810]  & n2936;
  assign n4410 = \[5015]  & n2931;
  assign n4411 = \[5090]  & n2912_1;
  assign n4412 = \[10850]  & n2964;
  assign n4413_1 = \[4550]  & n2939;
  assign n4414 = ~n4412 & ~n4413_1;
  assign n4415 = \[5225]  & n2959;
  assign n4416 = \[15230]  & n2961;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418_1 = \[7220]  & n2955_1;
  assign n4419 = \[5300]  & n2916_1;
  assign n4420 = ~n4418_1 & ~n4419;
  assign n4421 = n4417 & n4420;
  assign n4422 = n4414 & n4421;
  assign n4423_1 = n2907_1 & ~n4422;
  assign n4424 = ~n4411 & ~n4423_1;
  assign n4425 = ~n4410 & n4424;
  assign n4426 = ~n4409 & n4425;
  assign n4427 = ~n2906 & ~n4426;
  assign n4428_1 = \[14060]  & n3081_1;
  assign n4429 = ~n4427 & ~n4428_1;
  assign n740 = ~n4408_1 | ~n4429;
  assign n4431 = \[4475]  & n3030;
  assign n4432 = \[10175]  & n2964;
  assign n4433_1 = \[6350]  & n3044;
  assign n4434 = ~n4432 & ~n4433_1;
  assign n4435 = \[14405]  & n3020;
  assign n4436 = \[5135]  & n2961;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438_1 = n4434 & n4437;
  assign n4439 = ~n4431 & n4438_1;
  assign n4440 = n2907_1 & ~n4439;
  assign n4441 = ppeakp_8_8_ & ~n3035;
  assign n4442 = \[15695]  & n2936;
  assign n4443_1 = ppeaka_8_8_ & ppeakb_8_8_;
  assign n4444 = n2912_1 & ~n4443_1;
  assign n4445 = \[11225]  & n3024;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = ~n4442 & n4446;
  assign n4448_1 = ~n4441 & n4447;
  assign n4449 = ~n4440 & n4448_1;
  assign n4450 = ~n2906 & ~n4449;
  assign n4451 = n2907_1 & ~n3050;
  assign n4452 = ppeakb_8_8_ & n4451;
  assign n4453_1 = n2907_1 & ~n3047;
  assign n4454 = \[6410]  & n4453_1;
  assign n4455 = ~n4452 & ~n4454;
  assign n4456 = ~n4450 & n4455;
  assign n4457 = ppeaka_8_8_ & ~n3042_1;
  assign n4458_1 = ppeaka_9_9_ & n2975_1;
  assign n4459 = ~n4457 & ~n4458_1;
  assign n744 = ~n4456 | ~n4459;
  assign n4461 = \[5720]  & ~n3065;
  assign n4462 = \[7265]  & n2917;
  assign n4463_1 = ~n4461 & ~n4462;
  assign n4464 = \[7550]  & n2931;
  assign n4465 = \[8945]  & n3068;
  assign n4466 = ~n4464 & ~n4465;
  assign n748 = ~n4463_1 | ~n4466;
  assign n4468 = ppeaks_14_14_ & ~n3090;
  assign n4469 = \[13070]  & n3081_1;
  assign n4470 = \[16070]  & n2959;
  assign n4471_1 = \[14270]  & n2949;
  assign n4472 = \[6215]  & n2964;
  assign n4473 = ~n4471_1 & ~n4472;
  assign n4474 = ~n4470 & n4473;
  assign n4475 = \[8735]  & n2939;
  assign n4476_1 = \[5435]  & n2955_1;
  assign n4477 = ~n4475 & ~n4476_1;
  assign n4478 = \[7400]  & n2961;
  assign n4479 = n4477 & ~n4478;
  assign n4480 = \[10985]  & n3046_1;
  assign n4481_1 = \[9560]  & n3020;
  assign n4482 = \[10055]  & n2916_1;
  assign n4483 = ~n4481_1 & ~n4482;
  assign n4484 = ~n4480 & n4483;
  assign n4485 = n4479 & n4484;
  assign n4486_1 = n4474 & n4485;
  assign n4487 = n2907_1 & ~n4486_1;
  assign n4488 = \[15410]  & n2931;
  assign n4489 = \[6725]  & n2936;
  assign n4490_1 = \[11900]  & n3095;
  assign n4491 = ~n4489 & ~n4490_1;
  assign n4492 = \[11375]  & n2912_1;
  assign n4493 = \[12650]  & n3024;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495_1 = n4491 & n4494;
  assign n4496 = ~n4488 & n4495_1;
  assign n4497 = ~n4487 & n4496;
  assign n4498 = ~n2906 & ~n4497;
  assign n4499 = ~n4469 & ~n4498;
  assign n753 = n4468 | ~n4499;
  assign n4501 = ppeaks_7_7_ & ~n3090;
  assign n4502 = \[15005]  & n3081_1;
  assign n4503 = \[13745]  & n2936;
  assign n4504 = \[6785]  & n2955_1;
  assign n4505_1 = \[8255]  & n3046_1;
  assign n4506 = \[12905]  & n2949;
  assign n4507 = ~n4505_1 & ~n4506;
  assign n4508 = ~n4504 & n4507;
  assign n4509 = \[6770]  & n2961;
  assign n4510_1 = \[11405]  & n2964;
  assign n4511 = ~n4509 & ~n4510_1;
  assign n4512 = \[12830]  & n2939;
  assign n4513 = n4511 & ~n4512;
  assign n4514 = \[6140]  & n2959;
  assign n4515_1 = \[8225]  & n3020;
  assign n4516 = \[4790]  & n2916_1;
  assign n4517 = ~n4515_1 & ~n4516;
  assign n4518 = ~n4514 & n4517;
  assign n4519_1 = n4513 & n4518;
  assign n4520 = n4508 & n4519_1;
  assign n4521 = n2907_1 & ~n4520;
  assign n4522 = ~n4503 & ~n4521;
  assign n4523 = \[9275]  & n2912_1;
  assign n4524_1 = \[11540]  & n3095;
  assign n4525 = ~n4149 & ~n4524_1;
  assign n4526 = ~n4523 & n4525;
  assign n4527 = \[14630]  & n2931;
  assign n4528 = n4526 & ~n4527;
  assign n4529_1 = n4522 & n4528;
  assign n4530 = ~n2906 & ~n4529_1;
  assign n4531 = ~n4502 & ~n4530;
  assign n757 = n4501 | ~n4531;
  assign n4533 = ppeakp_12_12_ & ~n3147;
  assign n4534_1 = ppeaka_12_12_ & ~n3156;
  assign n4535 = ppeakb_12_12_ & n2917;
  assign n4536 = ~n4534_1 & ~n4535;
  assign n4537 = ~n4533 & n4536;
  assign n4538_1 = \[11030]  & n3095;
  assign n4539 = \[11210]  & n3021;
  assign n4540 = \[8855]  & ~n2927;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~n4538_1 & n4541;
  assign n761 = ~n4537 | ~n4542;
  assign n4544 = ~\[5780]  & ~n3162;
  assign n4545 = ~pdata_2_2_ & n3162;
  assign n4546 = ~preset & ~n4545;
  assign n765 = ~n4544 & n4546;
  assign n4548_1 = ~pdata_4_4_ & n3175;
  assign n4549 = ~\[5795]  & ~n3175;
  assign n4550 = ~preset & ~n4549;
  assign n770 = ~n4548_1 & n4550;
  assign n4552 = ~pdata_8_8_ & n3175;
  assign n4553_1 = ~\[5810]  & ~n3175;
  assign n4554 = ~preset & ~n4553_1;
  assign n775 = ~n4552 & n4554;
  assign n4556 = pdata_9_9_ & n3192;
  assign n4557 = \[5825]  & n3194_1;
  assign n780 = n4556 | n4557;
  assign n4559 = pdata_4_4_ & n3192;
  assign n4560 = \[5840]  & n3194_1;
  assign n785 = n4559 | n4560;
  assign n4562_1 = pdata_11_11_ & n3192;
  assign n4563 = \[5855]  & n3194_1;
  assign n790 = n4562_1 | n4563;
  assign n4565 = ~\[5870]  & ~n3203;
  assign n4566_1 = ~pdata_6_6_ & n3203;
  assign n4567 = ~preset & ~n4566_1;
  assign n795 = ~n4565 & n4567;
  assign n4569 = ~pdata_5_5_ & n3208;
  assign n4570 = ~\[5885]  & ~n3208;
  assign n4571_1 = ~preset & ~n4570;
  assign n800 = ~n4569 & n4571_1;
  assign n4573 = ~\[5900]  & ~n3218;
  assign n4574 = ~pdata_0_0_ & n3218;
  assign n4575_1 = ~preset & ~n4574;
  assign n805 = ~n4573 & n4575_1;
  assign n4577 = ~\[5915]  & ~n3218;
  assign n4578 = ~pdata_7_7_ & n3218;
  assign n4579 = ~preset & ~n4578;
  assign n810 = ~n4577 & n4579;
  assign n4581 = ~\[5930]  & ~n3218;
  assign n4582 = ~pdata_11_11_ & n3218;
  assign n4583 = ~preset & ~n4582;
  assign n815 = ~n4581 & n4583;
  assign n4585_1 = ~\[5945]  & ~n3231;
  assign n4586 = ~pdata_12_12_ & n3231;
  assign n4587 = ~preset & ~n4586;
  assign n820 = ~n4585_1 & n4587;
  assign n4589 = pdata_7_7_ & n3238;
  assign n4590_1 = \[5960]  & n3240;
  assign n825 = n4589 | n4590_1;
  assign n4592 = pdata_14_14_ & n3238;
  assign n4593 = \[5975]  & n3240;
  assign n830 = n4592 | n4593;
  assign n4595_1 = pdata_9_9_ & n3238;
  assign n4596 = \[5990]  & n3240;
  assign n835 = n4595_1 | n4596;
  assign n4598 = ~\[6005]  & ~n3249_1;
  assign n4599_1 = ~pdata_8_8_ & n3249_1;
  assign n4600 = ~preset & ~n4599_1;
  assign n840 = ~n4598 & n4600;
  assign n4602 = ~n3486 & ~n3487_1;
  assign n4603 = ~n3490 & ~n4602;
  assign n4604 = n3490 & n4602;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = n4161 & n4605;
  assign n4607 = \[6020]  & n3312;
  assign n845 = n4606 | n4607;
  assign n4609 = n4161 & n3564;
  assign n4610 = \[6035]  & n3312;
  assign n850 = n4609 | n4610;
  assign n4612 = ~\[6050]  & ~n3265;
  assign n4613 = n3265 & n3667_1;
  assign n4614 = ~preset & ~n4613;
  assign n855 = ~n4612 & n4614;
  assign n4616 = n3192 & n3675;
  assign n4617 = \[6065]  & n3194_1;
  assign n860 = n4616 | n4617;
  assign n4619 = n3192 & ~n4326;
  assign n4620 = \[6080]  & n3194_1;
  assign n865 = n4619 | n4620;
  assign n4622 = ~\[6095]  & ~n3266;
  assign n4623 = n3405 & ~n3517_1;
  assign n4624 = n3406 & n3517_1;
  assign n4625 = n3519 & ~n4624;
  assign n4626 = ~n4623 & ~n4625;
  assign n4627 = n3266 & n4626;
  assign n4628 = ~preset & ~n4627;
  assign n870 = ~n4622 & n4628;
  assign n4630 = \[6110]  & n3574;
  assign n4631 = n3568 & ~n4344_1;
  assign n875 = n4630 | n4631;
  assign n4633 = ~\[6125]  & ~n3218;
  assign n4634 = n3218 & n4298;
  assign n4635 = ~preset & ~n4634;
  assign n880 = ~n4633 & n4635;
  assign n4637 = ~\[6140]  & ~n3218;
  assign n4638 = n3218 & ~n3675;
  assign n4639 = ~preset & ~n4638;
  assign n885 = ~n4637 & n4639;
  assign n4641 = ~\[6155]  & ~n3231;
  assign n4642 = n3231 & ~n3564;
  assign n4643 = ~preset & ~n4642;
  assign n890 = ~n4641 & n4643;
  assign n4645 = n3238 & n3572_1;
  assign n4646 = \[6170]  & n3240;
  assign n895 = n4645 | n4646;
  assign n4648 = n3556 & n3671;
  assign n4649 = \[6185]  & n3677_1;
  assign n900 = n4648 | n4649;
  assign n4651 = \[6200]  & n3682_1;
  assign n4652 = n3680 & n4605;
  assign n905 = n4651 | n4652;
  assign n4654 = \[6215]  & n3682_1;
  assign n4655 = n3680 & ~n4326;
  assign n910 = n4654 | n4655;
  assign n4657 = ~\[6230]  & ~n3691;
  assign n4658 = n3691 & ~n3966;
  assign n4659 = ~preset & ~n4658;
  assign n915 = ~n4657 & n4659;
  assign n4661 = ~\[6245]  & ~n3720;
  assign n4662 = n3720 & ~n4357;
  assign n4663 = ~preset & ~n4662;
  assign n920 = ~n4661 & n4663;
  assign n4665 = ~\[6260]  & ~n3707_1;
  assign n4666 = n3707_1 & ~n4104;
  assign n4667 = ~preset & ~n4666;
  assign n925 = ~n4665 & n4667;
  assign n4669 = ~\[6275]  & ~n3706;
  assign n4670 = ~n3831 & ~n3833_1;
  assign n4671 = n3824 & ~n4670;
  assign n4672 = ~n3832 & ~n4671;
  assign n4673 = n3706 & ~n4672;
  assign n4674 = ~preset & ~n4673;
  assign n930 = ~n4669 & n4674;
  assign n4676 = ~\[6290]  & ~n3706;
  assign n4677 = n3706 & n4365;
  assign n4678 = ~preset & ~n4677;
  assign n935 = ~n4676 & n4678;
  assign n4680 = \[6305]  & n4097_1;
  assign n4681 = n4091 & n4104;
  assign n940 = n4680 | n4681;
  assign n4683 = ~preset & ~n3696;
  assign n4684 = \[6320]  & n4683;
  assign n4685 = ~preset & n3696;
  assign n4686 = ~n4080 & n4685;
  assign n945 = n4684 | n4686;
  assign n4688 = \[6335]  & n3682_1;
  assign n4689 = ~n4073 & ~n4074;
  assign n4690 = ~n4075 & n4689;
  assign n4691 = n4075 & ~n4689;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = n3680 & ~n4692;
  assign n950 = n4688 | n4693;
  assign n4695 = \[6350]  & n4116;
  assign n4696 = n4114 & n4376;
  assign n955 = n4695 | n4696;
  assign n4698 = \[6365]  & n4116;
  assign n4699 = ~n4080 & n4114;
  assign n960 = n4698 | n4699;
  assign n4701 = ppeakb_11_11_ & ~n2989;
  assign n4702 = \[14480]  & n3081_1;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = \[15890]  & n2936;
  assign n4705 = \[4295]  & n2931;
  assign n4706 = \[4370]  & n2912_1;
  assign n4707 = \[4595]  & n2916_1;
  assign n4708 = \[5855]  & n2961;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = \[5930]  & n2959;
  assign n4711 = \[5255]  & n2939;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = \[14090]  & n2964;
  assign n4714 = \[9155]  & n2955_1;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4712 & n4715;
  assign n4717 = n4709 & n4716;
  assign n4718 = n2907_1 & ~n4717;
  assign n4719 = ~n4706 & ~n4718;
  assign n4720 = ~n4705 & n4719;
  assign n4721 = ~n4704 & n4720;
  assign n4722 = ~n2906 & ~n4721;
  assign n4723 = ppeaka_11_11_ & n4124;
  assign n4724 = ~n4722 & ~n4723;
  assign n965 = ~n4703 | ~n4724;
  assign n4726 = ppeakb_2_2_ & ~n2989;
  assign n4727 = \[14465]  & n3081_1;
  assign n4728 = ~n4726 & ~n4727;
  assign n4729 = \[5780]  & n2912_1;
  assign n4730 = \[15515]  & n2931;
  assign n4731 = \[7130]  & n2936;
  assign n4732 = \[4445]  & n2961;
  assign n4733 = \[8555]  & n2916_1;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = \[7310]  & n2964;
  assign n4736 = \[9140]  & n2955_1;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = \[15290]  & n2939;
  assign n4739 = \[13640]  & n2959;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = n4737 & n4740;
  assign n4742 = n4734 & n4741;
  assign n4743 = n2907_1 & ~n4742;
  assign n4744 = ~n4731 & ~n4743;
  assign n4745 = ~n4730 & n4744;
  assign n4746 = ~n4729 & n4745;
  assign n4747 = ~n2906 & ~n4746;
  assign n4748 = ppeaka_2_2_ & n4124;
  assign n4749 = ~n4747 & ~n4748;
  assign n969 = ~n4728 | ~n4749;
  assign n4751 = \[6410]  & ~n3065;
  assign n4752 = \[5630]  & n3068;
  assign n4753 = ~n4751 & ~n4752;
  assign n4754 = \[6920]  & n2931;
  assign n4755 = \[7895]  & n2917;
  assign n4756 = ~n4754 & ~n4755;
  assign n973 = ~n4753 | ~n4756;
  assign n4758 = \[7355]  & n2936;
  assign n4759 = \[15050]  & n2931;
  assign n4760 = \[12425]  & n3024;
  assign n4761 = \[10580]  & n2961;
  assign n4762 = \[6320]  & n3046_1;
  assign n4763 = \[4730]  & n2955_1;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = ~n4761 & n4764;
  assign n4766 = \[13880]  & n2949;
  assign n4767 = \[11180]  & n2964;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = \[9395]  & n2939;
  assign n4770 = n4768 & ~n4769;
  assign n4771 = \[4880]  & n3020;
  assign n4772 = \[8150]  & n2916_1;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = \[15725]  & n2959;
  assign n4775 = n4773 & ~n4774;
  assign n4776 = n4770 & n4775;
  assign n4777 = n4765 & n4776;
  assign n4778 = n2907_1 & ~n4777;
  assign n4779 = ~n4760 & ~n4778;
  assign n4780 = \[15320]  & n2912_1;
  assign n4781 = \[11780]  & n3095;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = n4779 & n4782;
  assign n4784 = ~n4759 & n4783;
  assign n4785 = ~n4758 & n4784;
  assign n4786 = ~n2906 & ~n4785;
  assign n4787 = ppeaks_15_15_ & ~n3090;
  assign n4788 = \[12365]  & n3081_1;
  assign n4789 = ~n4787 & ~n4788;
  assign n978 = n4786 | ~n4789;
  assign n4791 = \[14210]  & n2931;
  assign n4792 = \[14135]  & n2936;
  assign n4793 = \[8870]  & n3021;
  assign n4794 = ~n3025 & ~n4793;
  assign n4795 = \[8615]  & n2912_1;
  assign n4796 = n4794 & ~n4795;
  assign n4797 = ~n4792 & n4796;
  assign n4798 = \[5495]  & n2917;
  assign n4799 = \[13085]  & n2940_1;
  assign n4800 = ~n4798 & ~n4799;
  assign n4801 = \[11300]  & n3095;
  assign n4802 = \[11165]  & n2964;
  assign n4803 = \[8075]  & n2959;
  assign n4804 = \[10565]  & n2961;
  assign n4805 = \[13865]  & n2949;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~n4803 & n4806;
  assign n4808 = \[7625]  & n3046_1;
  assign n4809 = \[6110]  & n2955_1;
  assign n4810 = ~n4808 & ~n4809;
  assign n4811 = n4807 & n4810;
  assign n4812 = ~n4802 & n4811;
  assign n4813 = n2907_1 & ~n4812;
  assign n4814 = ~n4801 & ~n4813;
  assign n4815 = n4800 & n4814;
  assign n4816 = n4797 & n4815;
  assign n4817 = ~n4791 & n4816;
  assign n4818 = ~n2906 & ~n4817;
  assign n4819 = ppeaks_6_6_ & ~n3090;
  assign n4820 = \[16085]  & n3081_1;
  assign n4821 = ~n4819 & ~n4820;
  assign n982 = n4818 | ~n4821;
  assign n4823 = ppeakp_13_13_ & ~n3147;
  assign n4824 = ppeaka_13_13_ & ~n3156;
  assign n4825 = ppeakb_13_13_ & n2917;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = ~n4823 & n4826;
  assign n4828 = \[10760]  & n3095;
  assign n4829 = \[10955]  & n3021;
  assign n4830 = \[9530]  & ~n2927;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = ~n4828 & n4831;
  assign n986 = ~n4827 | ~n4832;
  assign n4834 = ~\[6470]  & ~n3162;
  assign n4835 = ~pdata_12_12_ & n3162;
  assign n4836 = ~preset & ~n4835;
  assign n990 = ~n4834 & n4836;
  assign n4838 = ~pdata_5_5_ & n3175;
  assign n4839 = ~\[6485]  & ~n3175;
  assign n4840 = ~preset & ~n4839;
  assign n995 = ~n4838 & n4840;
  assign n4842 = ~pdata_7_7_ & n3175;
  assign n4843 = ~\[6500]  & ~n3175;
  assign n4844 = ~preset & ~n4843;
  assign n1000 = ~n4842 & n4844;
  assign n4846 = pdata_10_10_ & n3192;
  assign n4847 = \[6515]  & n3194_1;
  assign n1005 = n4846 | n4847;
  assign n4849 = pdata_3_3_ & n3192;
  assign n4850 = \[6530]  & n3194_1;
  assign n1010 = n4849 | n4850;
  assign n4852 = pdata_12_12_ & n3192;
  assign n4853 = \[6545]  & n3194_1;
  assign n1015 = n4852 | n4853;
  assign n4855 = ~\[6560]  & ~n3203;
  assign n4856 = ~pdata_5_5_ & n3203;
  assign n4857 = ~preset & ~n4856;
  assign n1020 = ~n4855 & n4857;
  assign n4859 = ~pdata_6_6_ & n3208;
  assign n4860 = ~\[6575]  & ~n3208;
  assign n4861 = ~preset & ~n4860;
  assign n1025 = ~n4859 & n4861;
  assign n4863 = ~pdata_15_15_ & n3208;
  assign n4864 = ~\[6590]  & ~n3208;
  assign n4865 = ~preset & ~n4864;
  assign n1030 = ~n4863 & n4865;
  assign n4867 = ~\[6605]  & ~n3218;
  assign n4868 = ~pdata_8_8_ & n3218;
  assign n4869 = ~preset & ~n4868;
  assign n1035 = ~n4867 & n4869;
  assign n4871 = ~\[6620]  & ~n3231;
  assign n4872 = ~pdata_13_13_ & n3231;
  assign n4873 = ~preset & ~n4872;
  assign n1040 = ~n4871 & n4873;
  assign n4875 = n3177 & n3237;
  assign n4876 = \[6635]  & n3240;
  assign n1045 = n4875 | n4876;
  assign n4878 = pdata_15_15_ & n3238;
  assign n4879 = \[6650]  & n3240;
  assign n1050 = n4878 | n4879;
  assign n4881 = pdata_8_8_ & n3238;
  assign n4882 = \[6665]  & n3240;
  assign n1055 = n4881 | n4882;
  assign n4884 = ~\[6680]  & ~n3249_1;
  assign n4885 = ~pdata_9_9_ & n3249_1;
  assign n4886 = ~preset & ~n4885;
  assign n1060 = ~n4884 & n4886;
  assign n4888 = n4161 & n3660;
  assign n4889 = \[6695]  & n3312;
  assign n1065 = n4888 | n4889;
  assign n4891 = n4161 & ~n3549;
  assign n4892 = \[6710]  & n3312;
  assign n1070 = n4891 | n4892;
  assign n4894 = ~\[6725]  & ~n3265;
  assign n4895 = n3265 & n4326;
  assign n4896 = ~preset & ~n4895;
  assign n1075 = ~n4894 & n4896;
  assign n4898 = n3192 & ~n4344_1;
  assign n4899 = \[6740]  & n3194_1;
  assign n1080 = n4898 | n4899;
  assign n4901 = n3192 & ~n3646;
  assign n4902 = \[6755]  & n3194_1;
  assign n1085 = n4901 | n4902;
  assign n4904 = ~\[6770]  & ~n3266;
  assign n4905 = n3266 & ~n3675;
  assign n4906 = ~preset & ~n4905;
  assign n1090 = ~n4904 & n4906;
  assign n4908 = n3568 & n3675;
  assign n4909 = \[6785]  & n3574;
  assign n1095 = n4908 | n4909;
  assign n4911 = ~\[6815]  & ~n3218;
  assign n4912 = n3218 & n4626;
  assign n4913 = ~preset & ~n4912;
  assign n1100 = ~n4911 & n4913;
  assign n4915 = ~\[6830]  & ~n3231;
  assign n4916 = n3231 & n3549;
  assign n4917 = ~preset & ~n4916;
  assign n1105 = ~n4915 & n4917;
  assign n4919 = n3238 & n4605;
  assign n4920 = \[6845]  & n3240;
  assign n1110 = n4919 | n4920;
  assign n4922 = n3238 & n3541;
  assign n4923 = \[6860]  & n3240;
  assign n1115 = n4922 | n4923;
  assign n4925 = n3572_1 & n3680;
  assign n4926 = \[6875]  & n3682_1;
  assign n1120 = n4925 | n4926;
  assign n4928 = ~n3667_1 & n3680;
  assign n4929 = \[6890]  & n3682_1;
  assign n1125 = n4928 | n4929;
  assign n4931 = ~\[6905]  & ~n3691;
  assign n4932 = n3691 & ~n4399;
  assign n4933 = ~preset & ~n4932;
  assign n1130 = ~n4931 & n4933;
  assign n4935 = ~\[6920]  & ~n3720;
  assign n4936 = n3720 & ~n4376;
  assign n4937 = ~preset & ~n4936;
  assign n1135 = ~n4935 & n4937;
  assign n4939 = ~\[6935]  & ~n3707_1;
  assign n4940 = n3707_1 & ~n4672;
  assign n4941 = ~preset & ~n4940;
  assign n1140 = ~n4939 & n4941;
  assign n4943 = ~\[6950]  & ~n3706;
  assign n4944 = n3706 & ~n4104;
  assign n4945 = ~preset & ~n4944;
  assign n1145 = ~n4943 & n4945;
  assign n4947 = ~\[6965]  & ~n3706;
  assign n4948 = n3706 & n3958_1;
  assign n4949 = ~preset & ~n4948;
  assign n1150 = ~n4947 & n4949;
  assign n4951 = \[6980]  & n4097_1;
  assign n4952 = ~n3841 & ~n3842;
  assign n4953 = n3843_1 & ~n4952;
  assign n4954 = ~n3843_1 & n4952;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = n4091 & ~n4955;
  assign n1155 = n4951 | n4956;
  assign n4958 = n4399 & n4685;
  assign n4959 = \[6995]  & n4683;
  assign n1160 = n4958 | n4959;
  assign n4961 = \[7010]  & n3682_1;
  assign n4962 = n3680 & ~n4080;
  assign n1165 = n4961 | n4962;
  assign n4964 = \[7025]  & n4116;
  assign n4965 = n4114 & n4357;
  assign n1170 = n4964 | n4965;
  assign n4967 = \[7055]  & ~n3065;
  assign n4968 = \[11240]  & n3068;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = \[6245]  & n2931;
  assign n4971 = \[5960]  & n2917;
  assign n4972 = ~n4970 & ~n4971;
  assign n1175 = ~n4969 | ~n4972;
  assign n4974 = \[13775]  & n3081_1;
  assign n4975 = ppeaks_12_12_ & ~n3090;
  assign n4976 = \[12395]  & n2931;
  assign n4977 = \[14660]  & n3024;
  assign n4978 = \[10625]  & n2916_1;
  assign n4979 = \[8675]  & n2961;
  assign n4980 = \[10415]  & n3046_1;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = ~n4978 & n4981;
  assign n4983 = \[11615]  & n2959;
  assign n4984 = \[7460]  & n2939;
  assign n4985 = \[9365]  & n2955_1;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = ~n4983 & n4986;
  assign n4988 = \[9845]  & n3020;
  assign n4989 = \[4820]  & n2964;
  assign n4990 = \[15065]  & n2949;
  assign n4991 = ~n4989 & ~n4990;
  assign n4992 = ~n4988 & n4991;
  assign n4993 = n4987 & n4992;
  assign n4994 = n4982 & n4993;
  assign n4995 = n2907_1 & ~n4994;
  assign n4996 = \[4640]  & n2912_1;
  assign n4997 = \[5360]  & n2936;
  assign n4998 = \[9680]  & n3095;
  assign n4999 = ~n4997 & ~n4998;
  assign n5000 = ~n4996 & n4999;
  assign n5001 = ~n4995 & n5000;
  assign n5002 = ~n4977 & n5001;
  assign n5003 = ~n4976 & n5002;
  assign n5004 = ~n2906 & ~n5003;
  assign n5005 = ~n4975 & ~n5004;
  assign n1180 = n4974 | ~n5005;
  assign n5007 = \[14570]  & n3081_1;
  assign n5008 = ppeaks_1_1_ & ~n3090;
  assign n5009 = \[6305]  & n3024;
  assign n5010 = \[12380]  & n2931;
  assign n5011 = \[4625]  & n2912_1;
  assign n5012 = \[9665]  & n3095;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = \[16055]  & n2936;
  assign n5015 = \[4805]  & n2964;
  assign n5016 = \[8120]  & n2916_1;
  assign n5017 = \[8660]  & n2961;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = ~n5015 & n5018;
  assign n5020 = \[8045]  & n2955_1;
  assign n5021 = \[12005]  & n2949;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = \[15020]  & n2939;
  assign n5024 = n5022 & ~n5023;
  assign n5025 = \[11150]  & n2959;
  assign n5026 = \[12920]  & n3046_1;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = \[9830]  & n3020;
  assign n5029 = n5027 & ~n5028;
  assign n5030 = n5024 & n5029;
  assign n5031 = n5019 & n5030;
  assign n5032 = n2907_1 & ~n5031;
  assign n5033 = ~n5014 & ~n5032;
  assign n5034 = n5013 & n5033;
  assign n5035 = ~n5010 & n5034;
  assign n5036 = ~n5009 & n5035;
  assign n5037 = ~n2906 & ~n5036;
  assign n5038 = ~n5008 & ~n5037;
  assign n1184 = n5007 | ~n5038;
  assign n5040 = ppeakp_3_3_ & ~n3147;
  assign n5041 = ppeaka_3_3_ & ~n3156;
  assign n5042 = ppeakb_3_3_ & n2917;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = ~n5040 & n5043;
  assign n5045 = \[15785]  & n3095;
  assign n5046 = \[11195]  & n3021;
  assign n5047 = \[7565]  & ~n2927;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = ~n5045 & n5048;
  assign n1188 = ~n5044 | ~n5049;
  assign n5051 = ~\[7115]  & ~n3162;
  assign n5052 = ~pdata_7_7_ & n3162;
  assign n5053 = ~preset & ~n5052;
  assign n1192 = ~n5051 & n5053;
  assign n5055 = ~pdata_2_2_ & n3175;
  assign n5056 = ~\[7130]  & ~n3175;
  assign n5057 = ~preset & ~n5056;
  assign n1197 = ~n5055 & n5057;
  assign n5059 = \[7145]  & n3194_1;
  assign n1202 = n4562_1 | n5059;
  assign n5061 = n3177 & n3191;
  assign n5062 = \[7160]  & n3194_1;
  assign n1207 = n5061 | n5062;
  assign n5064 = ~\[7175]  & ~n3203;
  assign n5065 = ~pdata_1_1_ & n3203;
  assign n5066 = ~preset & ~n5065;
  assign n1212 = ~n5064 & n5066;
  assign n5068 = ~\[7190]  & ~n3203;
  assign n5069 = ~pdata_12_12_ & n3203;
  assign n5070 = ~preset & ~n5069;
  assign n1217 = ~n5068 & n5070;
  assign n5072 = ~\[7205]  & ~n3203;
  assign n5073 = ~pdata_15_15_ & n3203;
  assign n5074 = ~preset & ~n5073;
  assign n1222 = ~n5072 & n5074;
  assign n5076 = ~pdata_10_10_ & n3208;
  assign n5077 = ~\[7220]  & ~n3208;
  assign n5078 = ~preset & ~n5077;
  assign n1227 = ~n5076 & n5078;
  assign n5080 = ~\[7235]  & ~n3218;
  assign n5081 = ~pdata_5_5_ & n3218;
  assign n5082 = ~preset & ~n5081;
  assign n1232 = ~n5080 & n5082;
  assign n5084 = ~\[7250]  & ~n3231;
  assign n5085 = ~pdata_14_14_ & n3231;
  assign n5086 = ~preset & ~n5085;
  assign n1237 = ~n5084 & n5086;
  assign n5088 = \[7265]  & n3240;
  assign n1242 = n4595_1 | n5088;
  assign n5090 = \[7280]  & n3240;
  assign n1247 = n4283 | n5090;
  assign n5092 = \[7295]  & n3240;
  assign n1252 = n4878 | n5092;
  assign n5094 = ~\[7310]  & ~n3249_1;
  assign n5095 = ~pdata_2_2_ & n3249_1;
  assign n5096 = ~preset & ~n5095;
  assign n1257 = ~n5094 & n5096;
  assign n5098 = ~\[7325]  & ~n3249_1;
  assign n5099 = ~pdata_13_13_ & n3249_1;
  assign n5100 = ~preset & ~n5099;
  assign n1262 = ~n5098 & n5100;
  assign n5102 = n4161 & ~n4626;
  assign n5103 = \[7340]  & n3312;
  assign n1267 = n5102 | n5103;
  assign n5105 = ~\[7355]  & ~n3265;
  assign n5106 = n3265 & n3646;
  assign n5107 = ~preset & ~n5106;
  assign n1272 = ~n5105 & n5107;
  assign n5109 = n3192 & n3653_1;
  assign n5110 = \[7370]  & n3194_1;
  assign n1277 = n5109 | n5110;
  assign n5112 = ~\[7385]  & ~n3266;
  assign n5113 = n3266 & ~n4605;
  assign n5114 = ~preset & ~n5113;
  assign n1282 = ~n5112 & n5114;
  assign n5116 = ~\[7400]  & ~n3266;
  assign n5117 = n3266 & n4326;
  assign n5118 = ~preset & ~n5117;
  assign n1287 = ~n5116 & n5118;
  assign n5120 = \[7415]  & n3574;
  assign n5121 = n3568 & ~n4298;
  assign n1292 = n5120 | n5121;
  assign n5123 = ~n3549 & n3568;
  assign n5124 = \[7430]  & n3574;
  assign n1297 = n5123 | n5124;
  assign n5126 = ~\[7445]  & ~n3218;
  assign n5127 = n3218 & ~n3556;
  assign n5128 = ~preset & ~n5127;
  assign n1302 = ~n5126 & n5128;
  assign n5130 = ~\[7460]  & ~n3231;
  assign n5131 = n3231 & ~n3541;
  assign n5132 = ~preset & ~n5131;
  assign n1307 = ~n5130 & n5132;
  assign n5134 = n3238 & ~n4344_1;
  assign n5135 = \[7475]  & n3240;
  assign n1312 = n5134 | n5135;
  assign n5137 = \[7490]  & n3677_1;
  assign n5138 = n3671 & ~n4298;
  assign n1317 = n5137 | n5138;
  assign n5140 = ~n3549 & n3671;
  assign n5141 = \[7505]  & n3677_1;
  assign n1322 = n5140 | n5141;
  assign n5143 = n3680 & ~n4626;
  assign n5144 = \[7520]  & n3682_1;
  assign n1327 = n5143 | n5144;
  assign n5146 = ~\[7535]  & ~n3691;
  assign n5147 = n3691 & n4955;
  assign n5148 = ~preset & ~n5147;
  assign n1332 = ~n5146 & n5148;
  assign n5150 = ~\[7550]  & ~n3720;
  assign n5151 = n3720 & ~n4087_1;
  assign n5152 = ~preset & ~n5151;
  assign n1337 = ~n5150 & n5152;
  assign n5154 = ~\[7565]  & ~n3707_1;
  assign n5155 = n3707_1 & ~n4095;
  assign n5156 = ~preset & ~n5155;
  assign n1342 = ~n5154 & n5156;
  assign n5158 = ~\[7580]  & ~n3707_1;
  assign n5159 = n3707_1 & n4692;
  assign n5160 = ~preset & ~n5159;
  assign n1347 = ~n5158 & n5160;
  assign n5162 = \[7595]  & n3968_1;
  assign n5163 = n3962 & n4376;
  assign n1352 = n5162 | n5163;
  assign n5165 = ~n3866 & n4685;
  assign n5166 = \[7625]  & n4683;
  assign n1357 = n5165 | n5166;
  assign n5168 = n4082 & n4672;
  assign n5169 = \[7640]  & n4385;
  assign n1362 = n5168 | n5169;
  assign n5171 = ~n4365 & n4082;
  assign n5172 = \[7655]  & n4385;
  assign n1367 = n5171 | n5172;
  assign n5174 = \[7670]  & n3682_1;
  assign n5175 = n3680 & n4399;
  assign n1372 = n5174 | n5175;
  assign n5177 = \[7685]  & ~n3065;
  assign n5178 = \[10430]  & n3068;
  assign n5179 = ~n5177 & ~n5178;
  assign n5180 = \[12410]  & n2931;
  assign n5181 = \[6635]  & n2917;
  assign n5182 = ~n5180 & ~n5181;
  assign n1377 = ~n5179 | ~n5182;
  assign n5184 = ppeaks_13_13_ & ~n3090;
  assign n5185 = \[12815]  & n3081_1;
  assign n5186 = \[12620]  & n2931;
  assign n5187 = \[5345]  & n2912_1;
  assign n5188 = \[12035]  & n3095;
  assign n5189 = \[14690]  & n2949;
  assign n5190 = \[8030]  & n2961;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = \[8885]  & n3020;
  assign n5193 = \[14990]  & n2959;
  assign n5194 = ~n5192 & ~n5193;
  assign n5195 = \[8705]  & n2955_1;
  assign n5196 = \[10700]  & n3046_1;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = \[6890]  & n2964;
  assign n5199 = n5197 & ~n5198;
  assign n5200 = n5194 & n5199;
  assign n5201 = n5191 & n5200;
  assign n5202 = \[8090]  & n2939;
  assign n5203 = n5201 & ~n5202;
  assign n5204 = n2907_1 & ~n5203;
  assign n5205 = ~n5188 & ~n5204;
  assign n5206 = ~n5187 & n5205;
  assign n5207 = \[6050]  & n2936;
  assign n5208 = \[14240]  & n3024;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = \[10340]  & n2917;
  assign n5211 = n5209 & ~n5210;
  assign n5212 = n5206 & n5211;
  assign n5213 = ~n5186 & n5212;
  assign n5214 = ~n2906 & ~n5213;
  assign n5215 = ~n5185 & ~n5214;
  assign n1382 = n5184 | ~n5215;
  assign n5217 = ppeakp_7_7_ & ~n3147;
  assign n5218 = \[14285]  & n3095;
  assign n5219 = ppeaka_7_7_ & ~n3156;
  assign n5220 = ppeakb_7_7_ & n2917;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = \[8900]  & n3021;
  assign n5223 = \[9815]  & ~n2927;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = n5221 & n5224;
  assign n5226 = ~n5218 & n5225;
  assign n1386 = n5217 | ~n5226;
  assign n5228 = ppeakp_2_2_ & ~n3147;
  assign n5229 = ppeaka_2_2_ & ~n3156;
  assign n5230 = \[10940]  & n3021;
  assign n5231 = ~n5229 & ~n5230;
  assign n5232 = ~n5228 & n5231;
  assign n5233 = ndout & n3095;
  assign n5234 = ppeakb_2_2_ & n2917;
  assign n5235 = \[8195]  & ~n2927;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = ~n5233 & n5236;
  assign n1390 = ~n5232 | ~n5237;
  assign n5239 = ~\[7745]  & ~n3162;
  assign n5240 = ~pdata_6_6_ & n3162;
  assign n5241 = ~preset & ~n5240;
  assign n1394 = ~n5239 & n5241;
  assign n5243 = ~pdata_3_3_ & n3175;
  assign n5244 = ~\[7760]  & ~n3175;
  assign n5245 = ~preset & ~n5244;
  assign n1399 = ~n5243 & n5245;
  assign n5247 = \[7775]  & n3194_1;
  assign n1404 = n4852 | n5247;
  assign n5249 = pdata_5_5_ & n3192;
  assign n5250 = \[7790]  & n3194_1;
  assign n1409 = n5249 | n5250;
  assign n5252 = ~\[7805]  & ~n3203;
  assign n5253 = ~pdata_2_2_ & n3203;
  assign n5254 = ~preset & ~n5253;
  assign n1414 = ~n5252 & n5254;
  assign n5256 = ~\[7820]  & ~n3203;
  assign n5257 = ~pdata_11_11_ & n3203;
  assign n5258 = ~preset & ~n5257;
  assign n1419 = ~n5256 & n5258;
  assign n5260 = ~pdata_0_0_ & n3208;
  assign n5261 = ~\[7835]  & ~n3208;
  assign n5262 = ~preset & ~n5261;
  assign n1424 = ~n5260 & n5262;
  assign n5264 = ~pdata_9_9_ & n3208;
  assign n5265 = ~\[7850]  & ~n3208;
  assign n5266 = ~preset & ~n5265;
  assign n1429 = ~n5264 & n5266;
  assign n5268 = ~\[7865]  & ~n3218;
  assign n5269 = ~pdata_6_6_ & n3218;
  assign n5270 = ~preset & ~n5269;
  assign n1434 = ~n5268 & n5270;
  assign n5272 = ~\[7880]  & ~n3231;
  assign n5273 = ~pdata_15_15_ & n3231;
  assign n5274 = ~preset & ~n5273;
  assign n1439 = ~n5272 & n5274;
  assign n5276 = \[7895]  & n3240;
  assign n1444 = n4881 | n5276;
  assign n5278 = \[7910]  & n3240;
  assign n1449 = n3239_1 | n5278;
  assign n5280 = \[7925]  & n3240;
  assign n1454 = n4592 | n5280;
  assign n5282 = ~\[7940]  & ~n3249_1;
  assign n5283 = ~pdata_3_3_ & n3249_1;
  assign n5284 = ~preset & ~n5283;
  assign n1459 = ~n5282 & n5284;
  assign n5286 = ~\[7955]  & ~n3249_1;
  assign n5287 = ~pdata_12_12_ & n3249_1;
  assign n5288 = ~preset & ~n5287;
  assign n1464 = ~n5286 & n5288;
  assign n5290 = n4161 & n3653_1;
  assign n5291 = \[7970]  & n3312;
  assign n1469 = n5290 | n5291;
  assign n5293 = n3192 & ~n4626;
  assign n5294 = \[8000]  & n3194_1;
  assign n1474 = n5293 | n5294;
  assign n5296 = ~\[8015]  & ~n3266;
  assign n5297 = n3266 & ~n3572_1;
  assign n5298 = ~preset & ~n5297;
  assign n1479 = ~n5296 & n5298;
  assign n5300 = ~\[8030]  & ~n3266;
  assign n5301 = n3266 & n3667_1;
  assign n5302 = ~preset & ~n5301;
  assign n1484 = ~n5300 & n5302;
  assign n5304 = ~n3310 & n3568;
  assign n5305 = \[8045]  & n3574;
  assign n1489 = n5304 | n5305;
  assign n5307 = n3564 & n3568;
  assign n5308 = \[8060]  & n3574;
  assign n1494 = n5307 | n5308;
  assign n5310 = ~\[8075]  & ~n3218;
  assign n5311 = n3218 & n4344_1;
  assign n5312 = ~preset & ~n5311;
  assign n1499 = ~n5310 & n5312;
  assign n5314 = ~\[8090]  & ~n3231;
  assign n5315 = n3231 & n3667_1;
  assign n5316 = ~preset & ~n5315;
  assign n1504 = ~n5314 & n5316;
  assign n5318 = n3238 & n3556;
  assign n5319 = \[8105]  & n3240;
  assign n1509 = n5318 | n5319;
  assign n5321 = \[8120]  & n3677_1;
  assign n5322 = ~n3310 & n3671;
  assign n1514 = n5321 | n5322;
  assign n5324 = n3564 & n3671;
  assign n5325 = \[8135]  & n3677_1;
  assign n1519 = n5324 | n5325;
  assign n5327 = \[8150]  & n3677_1;
  assign n5328 = ~n3646 & n3671;
  assign n1524 = n5327 | n5328;
  assign n5330 = ~\[8165]  & ~n3691;
  assign n5331 = n3691 & ~n4095;
  assign n5332 = ~preset & ~n5331;
  assign n1529 = ~n5330 & n5332;
  assign n5334 = ~\[8180]  & ~n3720;
  assign n5335 = n3720 & n3958_1;
  assign n5336 = ~preset & ~n5335;
  assign n1534 = ~n5334 & n5336;
  assign n5338 = ~\[8195]  & ~n3707_1;
  assign n5339 = n3707_1 & n4955;
  assign n5340 = ~preset & ~n5339;
  assign n1539 = ~n5338 & n5340;
  assign n5342 = ~\[8210]  & ~n3707_1;
  assign n5343 = n3707_1 & n4080;
  assign n5344 = ~preset & ~n5343;
  assign n1544 = ~n5342 & n5344;
  assign n5346 = \[8225]  & n3968_1;
  assign n5347 = n3962 & n4357;
  assign n1549 = n5346 | n5347;
  assign n5349 = \[8240]  & n4097_1;
  assign n5350 = n4091 & n4672;
  assign n1554 = n5349 | n5350;
  assign n5352 = n4357 & n4685;
  assign n5353 = \[8255]  & n4683;
  assign n1559 = n5352 | n5353;
  assign n5355 = n4111 & n4082;
  assign n5356 = \[8285]  & n4385;
  assign n1564 = n5355 | n5356;
  assign n5358 = \[8300]  & n3682_1;
  assign n5359 = n3680 & n3966;
  assign n1569 = n5358 | n5359;
  assign n5361 = \[8315]  & n4116;
  assign n5362 = n4114 & ~n4692;
  assign n1574 = n5361 | n5362;
  assign n5364 = \[8330]  & ~n3065;
  assign n5365 = \[4565]  & n2917;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = \[12635]  & n2931;
  assign n5368 = \[10715]  & n3068;
  assign n5369 = ~n5367 & ~n5368;
  assign n1579 = ~n5366 | ~n5369;
  assign n5371 = \[12575]  & n3081_1;
  assign n5372 = ppeaks_3_3_ & ~n3090;
  assign n5373 = \[15350]  & n2936;
  assign n5374 = \[4910]  & n3024;
  assign n5375 = \[12155]  & n3095;
  assign n5376 = ~n5374 & ~n5375;
  assign n5377 = ~n5373 & n5376;
  assign n5378 = \[12845]  & n2931;
  assign n5379 = \[6020]  & n2912_1;
  assign n5380 = \[8720]  & n2959;
  assign n5381 = \[6200]  & n2964;
  assign n5382 = \[10610]  & n2916_1;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = ~n5380 & n5383;
  assign n5385 = \[12455]  & n3046_1;
  assign n5386 = \[14255]  & n2949;
  assign n5387 = \[14180]  & n2939;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = ~n5385 & n5388;
  assign n5390 = \[5570]  & n3020;
  assign n5391 = \[9350]  & n2955_1;
  assign n5392 = \[7385]  & n2961;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394 = ~n5390 & n5393;
  assign n5395 = n5389 & n5394;
  assign n5396 = n5384 & n5395;
  assign n5397 = n2907_1 & ~n5396;
  assign n5398 = ~n5379 & ~n5397;
  assign n5399 = ~n5378 & n5398;
  assign n5400 = n5377 & n5399;
  assign n5401 = ~n2906 & ~n5400;
  assign n5402 = ~n5372 & ~n5401;
  assign n1584 = n5371 | ~n5402;
  assign n5404 = ppeakp_8_8_ & ~n3147;
  assign n5405 = ppeaka_8_8_ & ~n3156;
  assign n5406 = \[5600]  & n3021;
  assign n5407 = ~n5405 & ~n5406;
  assign n5408 = ~n5404 & n5407;
  assign n5409 = \[13895]  & n3095;
  assign n5410 = ppeakb_8_8_ & n2917;
  assign n5411 = \[10655]  & ~n2927;
  assign n5412 = ~n5410 & ~n5411;
  assign n5413 = ~n5409 & n5412;
  assign n1588 = ~n5408 | ~n5413;
  assign n5415 = ppeakp_1_1_ & ~n3147;
  assign n5416 = ppeaka_1_1_ & ~n3156;
  assign n5417 = \[6950]  & n3021;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = ~n5415 & n5418;
  assign n5420 = \[4970]  & n3095;
  assign n5421 = ppeakb_1_1_ & n2917;
  assign n5422 = \[6260]  & ~n2927;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = ~n5420 & n5423;
  assign n1592 = ~n5419 | ~n5424;
  assign n5426 = ~\[8390]  & ~n3162;
  assign n5427 = ~pdata_9_9_ & n3162;
  assign n5428 = ~preset & ~n5427;
  assign n1596 = ~n5426 & n5428;
  assign n5430 = ~pdata_0_0_ & n3175;
  assign n5431 = ~\[8405]  & ~n3175;
  assign n5432 = ~preset & ~n5431;
  assign n1601 = ~n5430 & n5432;
  assign n5434 = \[8420]  & n3194_1;
  assign n1606 = n3200 | n5434;
  assign n5436 = \[8435]  & n3194_1;
  assign n1611 = n4251 | n5436;
  assign n5438 = pdata_15_15_ & n3192;
  assign n5439 = \[8450]  & n3194_1;
  assign n1616 = n5438 | n5439;
  assign n5441 = ~\[8465]  & ~n3203;
  assign n5442 = ~pdata_10_10_ & n3203;
  assign n5443 = ~preset & ~n5442;
  assign n1621 = ~n5441 & n5443;
  assign n5445 = ~pdata_1_1_ & n3208;
  assign n5446 = ~\[8480]  & ~n3208;
  assign n5447 = ~preset & ~n5446;
  assign n1626 = ~n5445 & n5447;
  assign n5449 = ~pdata_12_12_ & n3208;
  assign n5450 = ~\[8495]  & ~n3208;
  assign n5451 = ~preset & ~n5450;
  assign n1631 = ~n5449 & n5451;
  assign n5453 = ~\[8510]  & ~n3218;
  assign n5454 = ~pdata_3_3_ & n3218;
  assign n5455 = ~preset & ~n5454;
  assign n1636 = ~n5453 & n5455;
  assign n5457 = \[8525]  & n3240;
  assign n1641 = n3243 | n5457;
  assign n5459 = \[8540]  & n3240;
  assign n1646 = n3246 | n5459;
  assign n5461 = pdata_2_2_ & n3238;
  assign n5462 = \[8555]  & n3240;
  assign n1651 = n5461 | n5462;
  assign n5464 = pdata_13_13_ & n3238;
  assign n5465 = \[8570]  & n3240;
  assign n1656 = n5464 | n5465;
  assign n5467 = ~\[8585]  & ~n3249_1;
  assign n5468 = ~pdata_4_4_ & n3249_1;
  assign n5469 = ~preset & ~n5468;
  assign n1661 = ~n5467 & n5469;
  assign n5471 = ~\[8600]  & ~n3249_1;
  assign n5472 = ~pdata_15_15_ & n3249_1;
  assign n5473 = ~preset & ~n5472;
  assign n1666 = ~n5471 & n5473;
  assign n5475 = n4161 & ~n4344_1;
  assign n5476 = \[8615]  & n3312;
  assign n1671 = n5475 | n5476;
  assign n5478 = \[8630]  & n3194_1;
  assign n5479 = n3192 & ~n4298;
  assign n1676 = n5478 | n5479;
  assign n5481 = n3192 & ~n3549;
  assign n5482 = \[8645]  & n3194_1;
  assign n1681 = n5481 | n5482;
  assign n5484 = ~\[8660]  & ~n3266;
  assign n5485 = n3266 & n3310;
  assign n5486 = ~preset & ~n5485;
  assign n1686 = ~n5484 & n5486;
  assign n5488 = ~\[8675]  & ~n3266;
  assign n5489 = n3266 & ~n3541;
  assign n5490 = ~preset & ~n5489;
  assign n1691 = ~n5488 & n5490;
  assign n5492 = n3568 & n3660;
  assign n5493 = \[8690]  & n3574;
  assign n1696 = n5492 | n5493;
  assign n5495 = n3568 & ~n3667_1;
  assign n5496 = \[8705]  & n3574;
  assign n1701 = n5495 | n5496;
  assign n5498 = ~\[8720]  & ~n3218;
  assign n5499 = n3218 & ~n4605;
  assign n5500 = ~preset & ~n5499;
  assign n1706 = ~n5498 & n5500;
  assign n5502 = ~\[8735]  & ~n3231;
  assign n5503 = n3231 & n4326;
  assign n5504 = ~preset & ~n5503;
  assign n1711 = ~n5502 & n5504;
  assign n5506 = n3238 & ~n4626;
  assign n5507 = \[8750]  & n3240;
  assign n1716 = n5506 | n5507;
  assign n5509 = n3238 & ~n3646;
  assign n5510 = \[8765]  & n3240;
  assign n1721 = n5509 | n5510;
  assign n5512 = \[8780]  & n3677_1;
  assign n5513 = n3653_1 & n3671;
  assign n1726 = n5512 | n5513;
  assign n5515 = n3564 & n3680;
  assign n5516 = \[8810]  & n3682_1;
  assign n1731 = n5515 | n5516;
  assign n5518 = ~\[8825]  & ~n3720;
  assign n5519 = n3720 & n4365;
  assign n5520 = ~preset & ~n5519;
  assign n1736 = ~n5518 & n5520;
  assign n5522 = ~\[8840]  & ~n3707_1;
  assign n5523 = n3707_1 & ~n4399;
  assign n5524 = ~preset & ~n5523;
  assign n1741 = ~n5522 & n5524;
  assign n5526 = ~\[8855]  & ~n3707_1;
  assign n5527 = n3707_1 & ~n4111;
  assign n5528 = ~preset & ~n5527;
  assign n1746 = ~n5526 & n5528;
  assign n5530 = ~n3866 & n3962;
  assign n5531 = \[8870]  & n3968_1;
  assign n1751 = n5530 | n5531;
  assign n5533 = \[8885]  & n3968_1;
  assign n5534 = n3962 & ~n4392;
  assign n1756 = n5533 | n5534;
  assign n5536 = ~\[8900]  & ~n3706;
  assign n5537 = n3706 & ~n4357;
  assign n5538 = ~preset & ~n5537;
  assign n1761 = ~n5536 & n5538;
  assign n5540 = n4376 & n4685;
  assign n5541 = \[8915]  & n4683;
  assign n1766 = n5540 | n5541;
  assign n5543 = n4082 & ~n4955;
  assign n5544 = \[8930]  & n4385;
  assign n1771 = n5543 | n5544;
  assign n5546 = n4087_1 & n4082;
  assign n5547 = \[8945]  & n4385;
  assign n1776 = n5546 | n5547;
  assign n5549 = \[8960]  & n3682_1;
  assign n5550 = n3680 & n4095;
  assign n1781 = n5549 | n5550;
  assign n5552 = n3966 & n4114;
  assign n5553 = \[8975]  & n4116;
  assign n1786 = n5552 | n5553;
  assign n5555 = \[6710]  & n2912_1;
  assign n5556 = \[13115]  & n2931;
  assign n5557 = \[4655]  & n2936;
  assign n5558 = \[13490]  & n3024;
  assign n5559 = \[10490]  & n3095;
  assign n5560 = \[12125]  & n2949;
  assign n5561 = \[7430]  & n2955_1;
  assign n5562 = \[10130]  & n3046_1;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = ~n5560 & n5563;
  assign n5565 = \[11390]  & n2959;
  assign n5566 = \[5525]  & n2964;
  assign n5567 = \[7505]  & n2916_1;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5565 & n5568;
  assign n5570 = \[10115]  & n3020;
  assign n5571 = \[9335]  & n2961;
  assign n5572 = ~n5570 & ~n5571;
  assign n5573 = \[6830]  & n2939;
  assign n5574 = n5572 & ~n5573;
  assign n5575 = n5569 & n5574;
  assign n5576 = n5564 & n5575;
  assign n5577 = n2907_1 & ~n5576;
  assign n5578 = ~n5559 & ~n5577;
  assign n5579 = ~n5558 & n5578;
  assign n5580 = ~n5557 & n5579;
  assign n5581 = ~n5556 & n5580;
  assign n5582 = ~n5555 & n5581;
  assign n5583 = ~n2906 & ~n5582;
  assign n5584 = ppeaks_11_11_ & ~n3090;
  assign n5585 = \[13415]  & n3081_1;
  assign n5586 = ~n5584 & ~n5585;
  assign n1791 = n5583 | ~n5586;
  assign n5588 = \[6980]  & n3024;
  assign n5589 = \[13100]  & n2931;
  assign n5590 = \[15710]  & n2936;
  assign n5591 = \[10325]  & n2916_1;
  assign n5592 = \[15425]  & n2949;
  assign n5593 = \[12680]  & n3046_1;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = ~n5591 & n5594;
  assign n5596 = \[9320]  & n2961;
  assign n5597 = \[8690]  & n2955_1;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = \[14600]  & n2939;
  assign n5600 = n5598 & ~n5599;
  assign n5601 = \[10100]  & n3020;
  assign n5602 = \[5510]  & n2964;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = \[10880]  & n2959;
  assign n5605 = n5603 & ~n5604;
  assign n5606 = n5600 & n5605;
  assign n5607 = n5595 & n5606;
  assign n5608 = n2907_1 & ~n5607;
  assign n5609 = ~n5590 & ~n5608;
  assign n5610 = \[6695]  & n2912_1;
  assign n5611 = \[10475]  & n3095;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = n5609 & n5612;
  assign n5614 = ~n5589 & n5613;
  assign n5615 = ~n5588 & n5614;
  assign n5616 = ~n2906 & ~n5615;
  assign n5617 = ppeaks_2_2_ & ~n3090;
  assign n5618 = \[14150]  & n3081_1;
  assign n5619 = ~n5617 & ~n5618;
  assign n1795 = n5616 | ~n5619;
  assign n5621 = ppeakp_9_9_ & ~n3147;
  assign n5622 = \[10370]  & ~n2927;
  assign n5623 = \[11750]  & n3095;
  assign n5624 = ppeakb_9_9_ & n2917;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~n5622 & n5625;
  assign n5627 = ppeaka_9_9_ & ~n3156;
  assign n5628 = \[4895]  & n3021;
  assign n5629 = ~n5627 & ~n5628;
  assign n5630 = n5626 & n5629;
  assign n1799 = n5621 | ~n5630;
  assign n5632 = ppeakp_0_0_ & ~n3147;
  assign n5633 = \[6935]  & ~n2927;
  assign n5634 = \[5675]  & n3095;
  assign n5635 = \[6275]  & n3021;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n5633 & n5636;
  assign n5638 = ppeaka_0_0_ & ~n3156;
  assign n5639 = ppeakb_0_0_ & n2917;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = n5637 & n5640;
  assign n1803 = n5632 | ~n5641;
  assign n5643 = ~\[9050]  & ~n3162;
  assign n5644 = ~pdata_8_8_ & n3162;
  assign n5645 = ~preset & ~n5644;
  assign n1807 = ~n5643 & n5645;
  assign n5647 = ~pdata_1_1_ & n3175;
  assign n5648 = ~\[9065]  & ~n3175;
  assign n5649 = ~preset & ~n5648;
  assign n1812 = ~n5647 & n5649;
  assign n5651 = \[9080]  & n3194_1;
  assign n1817 = n4257_1 | n5651;
  assign n5653 = \[9095]  & n3194_1;
  assign n1822 = n3193 | n5653;
  assign n5655 = ~\[9110]  & ~n3203;
  assign n5656 = ~pdata_0_0_ & n3203;
  assign n5657 = ~preset & ~n5656;
  assign n1827 = ~n5655 & n5657;
  assign n5659 = ~\[9125]  & ~n3203;
  assign n5660 = ~pdata_9_9_ & n3203;
  assign n5661 = ~preset & ~n5660;
  assign n1832 = ~n5659 & n5661;
  assign n5663 = ~pdata_2_2_ & n3208;
  assign n5664 = ~\[9140]  & ~n3208;
  assign n5665 = ~preset & ~n5664;
  assign n1837 = ~n5663 & n5665;
  assign n5667 = ~pdata_11_11_ & n3208;
  assign n5668 = ~\[9155]  & ~n3208;
  assign n5669 = ~preset & ~n5668;
  assign n1842 = ~n5667 & n5669;
  assign n5671 = ~\[9170]  & ~n3218;
  assign n5672 = ~pdata_4_4_ & n3218;
  assign n5673 = ~preset & ~n5672;
  assign n1847 = ~n5671 & n5673;
  assign n5675 = \[9185]  & n3240;
  assign n1852 = n4286_1 | n5675;
  assign n5677 = \[9200]  & n3240;
  assign n1857 = n4289 | n5677;
  assign n5679 = pdata_3_3_ & n3238;
  assign n5680 = \[9215]  & n3240;
  assign n1862 = n5679 | n5680;
  assign n5682 = pdata_12_12_ & n3238;
  assign n5683 = \[9230]  & n3240;
  assign n1867 = n5682 | n5683;
  assign n5685 = ~\[9245]  & ~n3249_1;
  assign n5686 = ~pdata_5_5_ & n3249_1;
  assign n5687 = ~preset & ~n5686;
  assign n1872 = ~n5685 & n5687;
  assign n5689 = ~\[9260]  & ~n3249_1;
  assign n5690 = ~pdata_14_14_ & n3249_1;
  assign n5691 = ~preset & ~n5690;
  assign n1877 = ~n5689 & n5691;
  assign n5693 = n4161 & n3675;
  assign n5694 = \[9275]  & n3312;
  assign n1882 = n5693 | n5694;
  assign n5696 = n3192 & ~n3310;
  assign n5697 = \[9290]  & n3194_1;
  assign n1887 = n5696 | n5697;
  assign n5699 = n3192 & n3564;
  assign n5700 = \[9305]  & n3194_1;
  assign n1892 = n5699 | n5700;
  assign n5702 = ~\[9320]  & ~n3266;
  assign n5703 = n3266 & ~n3660;
  assign n5704 = ~preset & ~n5703;
  assign n1897 = ~n5702 & n5704;
  assign n5706 = ~\[9335]  & ~n3266;
  assign n5707 = n3266 & n3549;
  assign n5708 = ~preset & ~n5707;
  assign n1902 = ~n5706 & n5708;
  assign n5710 = \[9350]  & n3574;
  assign n5711 = n3568 & n4605;
  assign n1907 = n5710 | n5711;
  assign n5713 = n3541 & n3568;
  assign n5714 = \[9365]  & n3574;
  assign n1912 = n5713 | n5714;
  assign n5716 = ~\[9380]  & ~n3218;
  assign n5717 = n3218 & ~n3572_1;
  assign n5718 = ~preset & ~n5717;
  assign n1917 = ~n5716 & n5718;
  assign n5720 = ~\[9395]  & ~n3231;
  assign n5721 = n3231 & n3646;
  assign n5722 = ~preset & ~n5721;
  assign n1922 = ~n5720 & n5722;
  assign n5724 = n3238 & n3675;
  assign n5725 = \[9410]  & n3240;
  assign n1927 = n5724 | n5725;
  assign n5727 = n3671 & ~n4626;
  assign n5728 = \[9440]  & n3677_1;
  assign n1932 = n5727 | n5728;
  assign n5730 = \[9455]  & n3682_1;
  assign n5731 = n3680 & ~n4298;
  assign n1937 = n5730 | n5731;
  assign n5733 = n3653_1 & n3680;
  assign n5734 = \[9470]  & n3682_1;
  assign n1942 = n5733 | n5734;
  assign n5736 = ~\[9485]  & ~n3691;
  assign n5737 = n3691 & ~n4104;
  assign n5738 = ~preset & ~n5737;
  assign n1947 = ~n5736 & n5738;
  assign n5740 = ~\[9500]  & ~n3720;
  assign n5741 = n3720 & ~n4111;
  assign n5742 = ~preset & ~n5741;
  assign n1952 = ~n5740 & n5742;
  assign n5744 = ~\[9515]  & ~n3707_1;
  assign n5745 = n3707_1 & ~n3966;
  assign n5746 = ~preset & ~n5745;
  assign n1957 = ~n5744 & n5746;
  assign n5748 = ~\[9530]  & ~n3707_1;
  assign n5749 = n3707_1 & n4392;
  assign n5750 = ~preset & ~n5749;
  assign n1962 = ~n5748 & n5750;
  assign n5752 = \[9545]  & n3968_1;
  assign n5753 = n3962 & n4399;
  assign n1967 = n5752 | n5753;
  assign n5755 = \[9560]  & n3968_1;
  assign n5756 = n3962 & ~n4692;
  assign n1972 = n5755 | n5756;
  assign n5758 = ~\[9575]  & ~n3706;
  assign n5759 = n3706 & n3866;
  assign n5760 = ~preset & ~n5759;
  assign n1977 = ~n5758 & n5760;
  assign n5762 = n4087_1 & n4685;
  assign n5763 = \[9590]  & n4683;
  assign n1982 = n5762 | n5763;
  assign n5765 = ~n4101 & n4082;
  assign n5766 = \[9605]  & n4385;
  assign n1987 = n5765 | n5766;
  assign n5768 = ~n3958_1 & n4082;
  assign n5769 = \[9620]  & n4385;
  assign n1992 = n5768 | n5769;
  assign n5771 = \[9635]  & n3682_1;
  assign n5772 = n3680 & ~n4955;
  assign n1997 = n5771 | n5772;
  assign n5774 = \[9650]  & n3682_1;
  assign n5775 = n3680 & ~n4365;
  assign n2002 = n5774 | n5775;
  assign n5777 = \[17414]  & ~\[17505] ;
  assign n5778 = ~\[9665]  & ~n5777;
  assign n5779 = ~pdata_1_1_ & n5777;
  assign n5780 = ~preset & ~n5779;
  assign n2007 = ~n5778 & n5780;
  assign n5782 = ~\[9680]  & ~n5777;
  assign n5783 = ~pdata_12_12_ & n5777;
  assign n5784 = ~preset & ~n5783;
  assign n2012 = ~n5782 & n5784;
  assign n5786 = \[12185]  & ~n2927;
  assign n5787 = ppeaki_10_10_ & ~n2861;
  assign n5788 = ppeaki_14_14_ & n2862_1;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = n2907_1 & ~n5789;
  assign n5791 = ~n5786 & ~n5790;
  assign n5792 = ~preset & ppeaki_6_6_;
  assign n5793 = ~n2984 & n5792;
  assign n2017 = ~n5791 | n5793;
  assign n5795 = \[9710]  & n3240;
  assign n2021 = n5461 | n5795;
  assign n5797 = n3192 & n3660;
  assign n5798 = \[9725]  & n3194_1;
  assign n2026 = n5797 | n5798;
  assign n5800 = n3192 & ~n3667_1;
  assign n5801 = \[9740]  & n3194_1;
  assign n2031 = n5800 | n5801;
  assign n5803 = n3238 & n3564;
  assign n5804 = \[9770]  & n3240;
  assign n2036 = n5803 | n5804;
  assign n5806 = n3572_1 & n3671;
  assign n5807 = \[9785]  & n3677_1;
  assign n2041 = n5806 | n5807;
  assign n5809 = ~\[9800]  & ~n3720;
  assign n5810 = n3720 & n4392;
  assign n5811 = ~preset & ~n5810;
  assign n2046 = ~n5809 & n5811;
  assign n5813 = ~\[9815]  & ~n3707_1;
  assign n5814 = n3707_1 & ~n4357;
  assign n5815 = ~preset & ~n5814;
  assign n2051 = ~n5813 & n5815;
  assign n5817 = \[9830]  & n3968_1;
  assign n5818 = n3962 & n4104;
  assign n2056 = n5817 | n5818;
  assign n5820 = \[9845]  & n3968_1;
  assign n5821 = n3962 & n4111;
  assign n2061 = n5820 | n5821;
  assign n5823 = ~n3958_1 & n4685;
  assign n5824 = \[9860]  & n4683;
  assign n2066 = n5823 | n5824;
  assign n5826 = n3966 & n4082;
  assign n5827 = \[9875]  & n4385;
  assign n2071 = n5826 | n5827;
  assign n5829 = ~n4080 & n4082;
  assign n5830 = \[9890]  & n4385;
  assign n2076 = n5829 | n5830;
  assign n5832 = \[9905]  & n3682_1;
  assign n5833 = n3680 & n4087_1;
  assign n2081 = n5832 | n5833;
  assign n5835 = n4095 & n4114;
  assign n5836 = \[9920]  & n4116;
  assign n2086 = n5835 | n5836;
  assign n5838 = ~\[9935]  & ~n5777;
  assign n5839 = ~pdata_0_0_ & n5777;
  assign n5840 = ~preset & ~n5839;
  assign n2091 = ~n5838 & n5840;
  assign n5842 = ~\[18142]  & \[18220] ;
  assign n5843 = ~\[9950]  & ~n5842;
  assign n5844 = ~pdata_6_6_ & n5842;
  assign n5845 = ~preset & ~n5844;
  assign n2096 = ~n5843 & n5845;
  assign n5847 = \[9980]  & n3240;
  assign n2101 = n5682 | n5847;
  assign n5849 = n3192 & n4605;
  assign n5850 = \[9995]  & n3194_1;
  assign n2106 = n5849 | n5850;
  assign n5852 = n3192 & n3541;
  assign n5853 = \[10010]  & n3194_1;
  assign n2111 = n5852 | n5853;
  assign n5855 = \[10025]  & n3240;
  assign n5856 = n3238 & ~n4298;
  assign n2116 = n5855 | n5856;
  assign n5858 = n3238 & n3653_1;
  assign n5859 = \[10040]  & n3240;
  assign n2121 = n5858 | n5859;
  assign n5861 = \[10055]  & n3677_1;
  assign n5862 = n3671 & ~n4326;
  assign n2126 = n5861 | n5862;
  assign n5864 = ~\[10070]  & ~n3720;
  assign n5865 = n3720 & n4692;
  assign n5866 = ~preset & ~n5865;
  assign n2131 = ~n5864 & n5866;
  assign n5868 = ~\[10085]  & ~n3707_1;
  assign n5869 = n3707_1 & n3866;
  assign n5870 = ~preset & ~n5869;
  assign n2136 = ~n5868 & n5870;
  assign n5872 = \[10100]  & n3968_1;
  assign n5873 = n3962 & ~n4955;
  assign n2141 = n5872 | n5873;
  assign n5875 = \[10115]  & n3968_1;
  assign n5876 = n3962 & ~n4365;
  assign n2146 = n5875 | n5876;
  assign n5878 = ~n4365 & n4685;
  assign n5879 = \[10130]  & n4683;
  assign n2151 = n5878 | n5879;
  assign n5881 = n4095 & n4082;
  assign n5882 = \[10145]  & n4385;
  assign n2156 = n5881 | n5882;
  assign n5884 = \[10175]  & n3682_1;
  assign n5885 = n3680 & n4376;
  assign n2161 = n5884 | n5885;
  assign n5887 = \[10190]  & n4116;
  assign n5888 = n4114 & ~n4392;
  assign n2166 = n5887 | n5888;
  assign n5890 = ~\[10205]  & ~n5777;
  assign n5891 = ~pdata_10_10_ & n5777;
  assign n5892 = ~preset & ~n5891;
  assign n2171 = ~n5890 & n5892;
  assign n5894 = ~\[10220]  & ~n5842;
  assign n5895 = ~pdata_5_5_ & n5842;
  assign n5896 = ~preset & ~n5895;
  assign n2176 = ~n5894 & n5896;
  assign n5898 = \[12200]  & ~n2927;
  assign n5899 = ppeaki_15_15_ & n2985;
  assign n2181 = n5898 | n5899;
  assign n5901 = ppeaki_4_4_ & n2985;
  assign n5902 = \[11930]  & ~n2927;
  assign n5903 = ppeaki_12_12_ & n2862_1;
  assign n5904 = ppeaki_8_8_ & ~n2861;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = n2907_1 & ~n5905;
  assign n5907 = ~n5902 & ~n5906;
  assign n2185 = n5901 | ~n5907;
  assign n5909 = \[10265]  & n3240;
  assign n2189 = n4875 | n5909;
  assign n5911 = ~\[10280]  & ~n3266;
  assign n5912 = n3266 & ~n3556;
  assign n5913 = ~preset & ~n5912;
  assign n2194 = ~n5911 & n5913;
  assign n5915 = n3238 & ~n3310;
  assign n5916 = \[10310]  & n3240;
  assign n2199 = n5915 | n5916;
  assign n5918 = n3660 & n3671;
  assign n5919 = \[10325]  & n3677_1;
  assign n2204 = n5918 | n5919;
  assign n5921 = ~n3667_1 & n3671;
  assign n5922 = \[10340]  & n3677_1;
  assign n2209 = n5921 | n5922;
  assign n5924 = ~\[10355]  & ~n3720;
  assign n5925 = n3720 & n4080;
  assign n5926 = ~preset & ~n5925;
  assign n2214 = ~n5924 & n5926;
  assign n5928 = ~\[10370]  & ~n3707_1;
  assign n5929 = n3707_1 & ~n4087_1;
  assign n5930 = ~preset & ~n5929;
  assign n2219 = ~n5928 & n5930;
  assign n5932 = ~n3958_1 & n3962;
  assign n5933 = \[10400]  & n3968_1;
  assign n2224 = n5932 | n5933;
  assign n5935 = n4111 & n4685;
  assign n5936 = \[10415]  & n4683;
  assign n2229 = n5935 | n5936;
  assign n5938 = ~n3866 & n4082;
  assign n5939 = \[10430]  & n4385;
  assign n2234 = n5938 | n5939;
  assign n5941 = n4082 & ~n4392;
  assign n5942 = \[10445]  & n4385;
  assign n2239 = n5941 | n5942;
  assign n5944 = \[10460]  & n3682_1;
  assign n5945 = n3680 & n4357;
  assign n2244 = n5944 | n5945;
  assign n5947 = ~\[10475]  & ~n5777;
  assign n5948 = ~pdata_2_2_ & n5777;
  assign n5949 = ~preset & ~n5948;
  assign n2249 = ~n5947 & n5949;
  assign n5951 = ~\[10490]  & ~n5777;
  assign n5952 = ~pdata_11_11_ & n5777;
  assign n5953 = ~preset & ~n5952;
  assign n2254 = ~n5951 & n5953;
  assign n5955 = ~\[10505]  & ~n5842;
  assign n5956 = ~pdata_4_4_ & n5842;
  assign n5957 = ~preset & ~n5956;
  assign n2259 = ~n5955 & n5957;
  assign n5959 = \[12080]  & ~n2927;
  assign n5960 = ppeaki_14_14_ & n2985;
  assign n2264 = n5959 | n5960;
  assign n5962 = \[11810]  & ~n2927;
  assign n5963 = ppeaki_13_13_ & n2862_1;
  assign n5964 = ppeaki_9_9_ & ~n2861;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = n2907_1 & ~n5965;
  assign n5967 = ~n5962 & ~n5966;
  assign n5968 = ~preset & ppeaki_5_5_;
  assign n5969 = ~n2984 & n5968;
  assign n2268 = ~n5967 | n5969;
  assign n5971 = ~\[10550]  & ~n3249_1;
  assign n5972 = ~pdata_0_0_ & n3249_1;
  assign n5973 = ~preset & ~n5972;
  assign n2272 = ~n5971 & n5973;
  assign n5975 = ~\[10565]  & ~n3266;
  assign n5976 = n3266 & n4344_1;
  assign n5977 = ~preset & ~n5976;
  assign n2277 = ~n5975 & n5977;
  assign n5979 = ~\[10580]  & ~n3266;
  assign n5980 = n3266 & n3646;
  assign n5981 = ~preset & ~n5980;
  assign n2282 = ~n5979 & n5981;
  assign n5983 = n3238 & ~n3549;
  assign n5984 = \[10595]  & n3240;
  assign n2287 = n5983 | n5984;
  assign n5986 = \[10610]  & n3677_1;
  assign n5987 = n3671 & n4605;
  assign n2292 = n5986 | n5987;
  assign n5989 = \[10625]  & n3677_1;
  assign n5990 = n3541 & n3671;
  assign n2297 = n5989 | n5990;
  assign n5992 = ~\[10655]  & ~n3707_1;
  assign n5993 = n3707_1 & ~n4376;
  assign n5994 = ~preset & ~n5993;
  assign n2302 = ~n5992 & n5994;
  assign n5996 = \[10670]  & n3968_1;
  assign n5997 = n3962 & n4672;
  assign n2307 = n5996 | n5997;
  assign n5999 = \[10685]  & n3968_1;
  assign n6000 = n3962 & n4087_1;
  assign n2312 = n5999 | n6000;
  assign n6002 = ~n4392 & n4685;
  assign n6003 = \[10700]  & n4683;
  assign n2317 = n6002 | n6003;
  assign n6005 = n4082 & n4399;
  assign n6006 = \[10715]  & n4385;
  assign n2322 = n6005 | n6006;
  assign n6008 = n4082 & ~n4692;
  assign n6009 = \[10730]  & n4385;
  assign n2327 = n6008 | n6009;
  assign n6011 = \[10745]  & n3682_1;
  assign n6012 = n3680 & ~n3866;
  assign n2332 = n6011 | n6012;
  assign n6014 = ~\[10760]  & ~n2843;
  assign n6015 = ~pdata_13_13_ & n2843;
  assign n6016 = ~preset & ~n6015;
  assign n2337 = ~n6014 & n6016;
  assign n6018 = ~\[10775]  & ~n5777;
  assign n6019 = ~pdata_8_8_ & n5777;
  assign n6020 = ~preset & ~n6019;
  assign n2342 = ~n6018 & n6020;
  assign n6022 = ~\[10790]  & ~n5842;
  assign n6023 = ~pdata_3_3_ & n5842;
  assign n6024 = ~preset & ~n6023;
  assign n2347 = ~n6022 & n6024;
  assign n6026 = \[17570]  & ~\[17635] ;
  assign n6027 = ~\[10805]  & ~n6026;
  assign n6028 = ~pdata_1_1_ & n6026;
  assign n6029 = ~preset & ~n6028;
  assign n2352 = ~n6027 & n6029;
  assign n6031 = ~\[10820]  & ~n6026;
  assign n6032 = ~pdata_12_12_ & n6026;
  assign n6033 = ~preset & ~n6032;
  assign n2357 = ~n6031 & n6033;
  assign n6035 = ~\[10850]  & ~n3249_1;
  assign n6036 = ~pdata_10_10_ & n3249_1;
  assign n6037 = ~preset & ~n6036;
  assign n2362 = ~n6035 & n6037;
  assign n6039 = n3568 & ~n4626;
  assign n6040 = \[10865]  & n3574;
  assign n2367 = n6039 | n6040;
  assign n6042 = ~\[10880]  & ~n3218;
  assign n6043 = n3218 & ~n3660;
  assign n6044 = ~preset & ~n6043;
  assign n2372 = ~n6042 & n6044;
  assign n6046 = n3556 & n3680;
  assign n6047 = \[10895]  & n3682_1;
  assign n2377 = n6046 | n6047;
  assign n6049 = ~\[10925]  & ~n3691;
  assign n6050 = n3691 & n3958_1;
  assign n6051 = ~preset & ~n6050;
  assign n2382 = ~n6049 & n6051;
  assign n6053 = ~\[10940]  & ~n3706;
  assign n6054 = n3706 & n4955;
  assign n6055 = ~preset & ~n6054;
  assign n2387 = ~n6053 & n6055;
  assign n6057 = ~\[10955]  & ~n3706;
  assign n6058 = n3706 & n4392;
  assign n6059 = ~preset & ~n6058;
  assign n2392 = ~n6057 & n6059;
  assign n6061 = \[10970]  & n4097_1;
  assign n6062 = n4091 & n4357;
  assign n2397 = n6061 | n6062;
  assign n6064 = n4685 & ~n4692;
  assign n6065 = \[10985]  & n4683;
  assign n2402 = n6064 | n6065;
  assign n6067 = ~n3958_1 & n4114;
  assign n6068 = \[11015]  & n4116;
  assign n2407 = n6067 | n6068;
  assign n6070 = ~\[11030]  & ~n2843;
  assign n6071 = ~pdata_12_12_ & n2843;
  assign n6072 = ~preset & ~n6071;
  assign n2412 = ~n6070 & n6072;
  assign n6074 = ~\[11045]  & ~n5777;
  assign n6075 = ~pdata_9_9_ & n5777;
  assign n6076 = ~preset & ~n6075;
  assign n2417 = ~n6074 & n6076;
  assign n6078 = ~\[11060]  & ~n5842;
  assign n6079 = ~pdata_2_2_ & n5842;
  assign n6080 = ~preset & ~n6079;
  assign n2422 = ~n6078 & n6080;
  assign n6082 = ~\[11075]  & ~n5842;
  assign n6083 = ~pdata_7_7_ & n5842;
  assign n6084 = ~preset & ~n6083;
  assign n2427 = ~n6082 & n6084;
  assign n6086 = ~\[11090]  & ~n6026;
  assign n6087 = ~pdata_13_13_ & n6026;
  assign n6088 = ~preset & ~n6087;
  assign n2432 = ~n6086 & n6088;
  assign n6090 = n4161 & n3572_1;
  assign n6091 = \[11120]  & n3312;
  assign n2437 = n6090 | n6091;
  assign n6093 = \[11135]  & n3574;
  assign n6094 = n3568 & n3653_1;
  assign n2442 = n6093 | n6094;
  assign n6096 = ~\[11150]  & ~n3218;
  assign n6097 = n3218 & n3310;
  assign n6098 = ~preset & ~n6097;
  assign n2447 = ~n6096 & n6098;
  assign n6100 = \[11165]  & n3682_1;
  assign n6101 = n3680 & ~n4344_1;
  assign n2452 = n6100 | n6101;
  assign n6103 = ~n3646 & n3680;
  assign n6104 = \[11180]  & n3682_1;
  assign n2457 = n6103 | n6104;
  assign n6106 = ~\[11195]  & ~n3706;
  assign n6107 = n3706 & ~n4095;
  assign n6108 = ~preset & ~n6107;
  assign n2462 = ~n6106 & n6108;
  assign n6110 = ~\[11210]  & ~n3706;
  assign n6111 = n3706 & ~n4111;
  assign n6112 = ~preset & ~n6111;
  assign n2467 = ~n6110 & n6112;
  assign n6114 = \[11225]  & n4097_1;
  assign n6115 = n4091 & n4376;
  assign n2472 = n6114 | n6115;
  assign n6117 = n4357 & n4082;
  assign n6118 = \[11240]  & n4385;
  assign n2477 = n6117 | n6118;
  assign n6120 = \[11255]  & n4116;
  assign n6121 = n4114 & n4672;
  assign n2482 = n6120 | n6121;
  assign n6123 = n4087_1 & n4114;
  assign n6124 = \[11270]  & n4116;
  assign n2487 = n6123 | n6124;
  assign n6126 = ~\[11285]  & ~n2843;
  assign n6127 = ~pdata_15_15_ & n2843;
  assign n6128 = ~preset & ~n6127;
  assign n2492 = ~n6126 & n6128;
  assign n6130 = ~\[11300]  & ~n5777;
  assign n6131 = ~pdata_6_6_ & n5777;
  assign n6132 = ~preset & ~n6131;
  assign n2497 = ~n6130 & n6132;
  assign n6134 = ~\[11315]  & ~n5842;
  assign n6135 = ~pdata_1_1_ & n5842;
  assign n6136 = ~preset & ~n6135;
  assign n2502 = ~n6134 & n6136;
  assign n6138 = ~\[11330]  & ~n5842;
  assign n6139 = ~pdata_8_8_ & n5842;
  assign n6140 = ~preset & ~n6139;
  assign n2507 = ~n6138 & n6140;
  assign n6142 = ~\[11345]  & ~n6026;
  assign n6143 = ~pdata_3_3_ & n6026;
  assign n6144 = ~preset & ~n6143;
  assign n2512 = ~n6142 & n6144;
  assign n6146 = n4161 & ~n4326;
  assign n6147 = \[11375]  & n3312;
  assign n2517 = n6146 | n6147;
  assign n6149 = ~\[11390]  & ~n3218;
  assign n6150 = n3218 & n3549;
  assign n6151 = ~preset & ~n6150;
  assign n2522 = ~n6149 & n6151;
  assign n6153 = n3675 & n3680;
  assign n6154 = \[11405]  & n3682_1;
  assign n2527 = n6153 | n6154;
  assign n6156 = ~\[11420]  & ~n3691;
  assign n6157 = n3691 & ~n4376;
  assign n6158 = ~preset & ~n6157;
  assign n2532 = ~n6156 & n6158;
  assign n6160 = ~\[11435]  & ~n3706;
  assign n6161 = n3706 & ~n3966;
  assign n6162 = ~preset & ~n6161;
  assign n2537 = ~n6160 & n6162;
  assign n6164 = ~\[11450]  & ~n3706;
  assign n6165 = n3706 & n4080;
  assign n6166 = ~preset & ~n6165;
  assign n2542 = ~n6164 & n6166;
  assign n6168 = \[11465]  & n4097_1;
  assign n6169 = n4091 & n4399;
  assign n2547 = n6168 | n6169;
  assign n6171 = \[11480]  & n3682_1;
  assign n6172 = n3680 & n4672;
  assign n2552 = n6171 | n6172;
  assign n6174 = n4104 & n4114;
  assign n6175 = \[11495]  & n4116;
  assign n2557 = n6174 | n6175;
  assign n6177 = n4111 & n4114;
  assign n6178 = \[11510]  & n4116;
  assign n2562 = n6177 | n6178;
  assign n6180 = ~\[11525]  & ~n2843;
  assign n6181 = ~pdata_14_14_ & n2843;
  assign n6182 = ~preset & ~n6181;
  assign n2567 = ~n6180 & n6182;
  assign n6184 = ~\[11540]  & ~n5777;
  assign n6185 = ~pdata_7_7_ & n5777;
  assign n6186 = ~preset & ~n6185;
  assign n2572 = ~n6184 & n6186;
  assign n6188 = ~\[11555]  & ~n5842;
  assign n6189 = ~pdata_0_0_ & n5842;
  assign n6190 = ~preset & ~n6189;
  assign n2577 = ~n6188 & n6190;
  assign n6192 = ~\[11570]  & ~n5842;
  assign n6193 = ~pdata_9_9_ & n5842;
  assign n6194 = ~preset & ~n6193;
  assign n2582 = ~n6192 & n6194;
  assign n6196 = ~\[11585]  & ~n6026;
  assign n6197 = ~pdata_2_2_ & n6026;
  assign n6198 = ~preset & ~n6197;
  assign n2587 = ~n6196 & n6198;
  assign n6200 = ~\[11600]  & ~n6026;
  assign n6201 = ~pdata_11_11_ & n6026;
  assign n6202 = ~preset & ~n6201;
  assign n2592 = ~n6200 & n6202;
  assign n6204 = ~\[11615]  & ~n3218;
  assign n6205 = n3218 & ~n3541;
  assign n6206 = ~preset & ~n6205;
  assign n2597 = ~n6204 & n6206;
  assign n6208 = ~\[11630]  & ~n3691;
  assign n6209 = n3691 & ~n4672;
  assign n6210 = ~preset & ~n6209;
  assign n2602 = ~n6208 & n6210;
  assign n6212 = ~\[11645]  & ~n3691;
  assign n6213 = n3691 & ~n4087_1;
  assign n6214 = ~preset & ~n6213;
  assign n2607 = ~n6212 & n6214;
  assign n6216 = ~\[11660]  & ~n3706;
  assign n6217 = n3706 & ~n4399;
  assign n6218 = ~preset & ~n6217;
  assign n2612 = ~n6216 & n6218;
  assign n6220 = ~\[11675]  & ~n3706;
  assign n6221 = n3706 & n4692;
  assign n6222 = ~preset & ~n6221;
  assign n2617 = ~n6220 & n6222;
  assign n6224 = ~n3866 & n4091;
  assign n6225 = \[11690]  & n4097_1;
  assign n2622 = n6224 | n6225;
  assign n6227 = \[11705]  & n3682_1;
  assign n6228 = n3680 & ~n3958_1;
  assign n2627 = n6227 | n6228;
  assign n6230 = \[11720]  & n4116;
  assign n6231 = n4114 & ~n4955;
  assign n2632 = n6230 | n6231;
  assign n6233 = \[11735]  & n4116;
  assign n6234 = n4114 & ~n4365;
  assign n2637 = n6233 | n6234;
  assign n6236 = ~\[11750]  & ~n2843;
  assign n6237 = ~pdata_9_9_ & n2843;
  assign n6238 = ~preset & ~n6237;
  assign n2642 = ~n6236 & n6238;
  assign n6240 = ~\[11765]  & ~n5777;
  assign n6241 = ~pdata_4_4_ & n5777;
  assign n6242 = ~preset & ~n6241;
  assign n2647 = ~n6240 & n6242;
  assign n6244 = ~\[11780]  & ~n5777;
  assign n6245 = ~pdata_15_15_ & n5777;
  assign n6246 = ~preset & ~n6245;
  assign n2652 = ~n6244 & n6246;
  assign n6248 = ~\[11795]  & ~n5842;
  assign n6249 = ~pdata_10_10_ & n5842;
  assign n6250 = ~preset & ~n6249;
  assign n2657 = ~n6248 & n6250;
  assign n6252 = ~\[11810]  & ~n6026;
  assign n6253 = ~pdata_5_5_ & n6026;
  assign n6254 = ~preset & ~n6253;
  assign n2662 = ~n6252 & n6254;
  assign n6256 = ppeaki_9_9_ & n2985;
  assign n6257 = \[12275]  & ~n2927;
  assign n6258 = ppeaki_13_13_ & ~n2861;
  assign n6259 = n2907_1 & n6258;
  assign n6260 = ~n6257 & ~n6259;
  assign n2667 = n6256 | ~n6260;
  assign n6262 = ppeakb_14_14_ & ~n2989;
  assign n6263 = ppeaka_14_14_ & n4124;
  assign n6264 = ~n6262 & ~n6263;
  assign n6265 = \[13235]  & n2912_1;
  assign n6266 = \[15140]  & n2931;
  assign n6267 = \[13250]  & n2936;
  assign n6268 = \[4505]  & n2955_1;
  assign n6269 = \[5165]  & n2961;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = \[15965]  & n2959;
  assign n6272 = \[7925]  & n2916_1;
  assign n6273 = ~n6271 & ~n6272;
  assign n6274 = \[9260]  & n2964;
  assign n6275 = \[7250]  & n2939;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = n6273 & n6276;
  assign n6278 = n6270 & n6277;
  assign n6279 = n2907_1 & ~n6278;
  assign n6280 = ~n6267 & ~n6279;
  assign n6281 = ~n6266 & n6280;
  assign n6282 = ~n6265 & n6281;
  assign n6283 = ~n2906 & ~n6282;
  assign n6284 = \[12770]  & n3081_1;
  assign n6285 = ~n6283 & ~n6284;
  assign n2671 = ~n6264 | ~n6285;
  assign n6287 = ~\[11885]  & ~n5777;
  assign n6288 = ~pdata_5_5_ & n5777;
  assign n6289 = ~preset & ~n6288;
  assign n2675 = ~n6287 & n6289;
  assign n6291 = ~\[11900]  & ~n5777;
  assign n6292 = ~pdata_14_14_ & n5777;
  assign n6293 = ~preset & ~n6292;
  assign n2680 = ~n6291 & n6293;
  assign n6295 = ~\[11915]  & ~n5842;
  assign n6296 = ~pdata_11_11_ & n5842;
  assign n6297 = ~preset & ~n6296;
  assign n2685 = ~n6295 & n6297;
  assign n6299 = ~\[11930]  & ~n6026;
  assign n6300 = ~pdata_4_4_ & n6026;
  assign n6301 = ~preset & ~n6300;
  assign n2690 = ~n6299 & n6301;
  assign n6303 = ppeaki_8_8_ & n2985;
  assign n6304 = ppeaki_12_12_ & ~n2861;
  assign n6305 = n2907_1 & n6304;
  assign n6306 = \[12485]  & ~n2927;
  assign n6307 = ~n6305 & ~n6306;
  assign n2695 = n6303 | ~n6307;
  assign n6309 = ppeakb_15_15_ & ~n2989;
  assign n6310 = \[13580]  & n2912_1;
  assign n6311 = \[14390]  & n2936;
  assign n6312 = ppeaka_15_15_ & ~n2950_1;
  assign n6313 = \[4535]  & n2952;
  assign n6314 = \[7880]  & n2939;
  assign n6315 = \[6590]  & n2955_1;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = \[8450]  & n2961;
  assign n6318 = n6316 & ~n6317;
  assign n6319 = ~n6313 & n6318;
  assign n6320 = \[15620]  & n2959;
  assign n6321 = \[7295]  & n2916_1;
  assign n6322 = \[8600]  & n2964;
  assign n6323 = ~n6321 & ~n6322;
  assign n6324 = ~n6320 & n6323;
  assign n6325 = n6319 & n6324;
  assign n6326 = ~n6312 & n6325;
  assign n6327 = n2907_1 & ~n6326;
  assign n6328 = \[13550]  & n2931;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = ~n6311 & n6329;
  assign n6331 = ~n6310 & n6330;
  assign n2699 = n6309 | ~n6331;
  assign n6333 = ~preset & n3698;
  assign n6334 = n4104 & n6333;
  assign n6335 = ~preset & ~n3698;
  assign n6336 = \[12005]  & n6335;
  assign n2703 = n6334 | n6336;
  assign n6338 = ~\[12020]  & ~n2843;
  assign n6339 = ~pdata_11_11_ & n2843;
  assign n6340 = ~preset & ~n6339;
  assign n2708 = ~n6338 & n6340;
  assign n6342 = ~\[12035]  & ~n5777;
  assign n6343 = ~pdata_13_13_ & n5777;
  assign n6344 = ~preset & ~n6343;
  assign n2713 = ~n6342 & n6344;
  assign n6346 = ~\[12050]  & ~n5842;
  assign n6347 = ~pdata_12_12_ & n5842;
  assign n6348 = ~preset & ~n6347;
  assign n2718 = ~n6346 & n6348;
  assign n6350 = ~\[12065]  & ~n6026;
  assign n6351 = ~pdata_7_7_ & n6026;
  assign n6352 = ~preset & ~n6351;
  assign n2723 = ~n6350 & n6352;
  assign n6354 = ~\[12080]  & ~n6026;
  assign n6355 = ~pdata_14_14_ & n6026;
  assign n6356 = ~preset & ~n6355;
  assign n2728 = ~n6354 & n6356;
  assign n6358 = \[12065]  & ~n2927;
  assign n6359 = ppeaki_11_11_ & ~n2861;
  assign n6360 = ppeaki_15_15_ & n2862_1;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = n2907_1 & ~n6361;
  assign n6363 = ~n6358 & ~n6362;
  assign n6364 = ~preset & ppeaki_7_7_;
  assign n6365 = ~n2984 & n6364;
  assign n2733 = ~n6363 | n6365;
  assign n6367 = ~n4365 & n6333;
  assign n6368 = \[12125]  & n6335;
  assign n2737 = n6367 | n6368;
  assign n6370 = ~\[12140]  & ~n2843;
  assign n6371 = ~pdata_10_10_ & n2843;
  assign n6372 = ~preset & ~n6371;
  assign n2742 = ~n6370 & n6372;
  assign n6374 = ~\[12155]  & ~n5777;
  assign n6375 = ~pdata_3_3_ & n5777;
  assign n6376 = ~preset & ~n6375;
  assign n2747 = ~n6374 & n6376;
  assign n6378 = ~\[12170]  & ~n5842;
  assign n6379 = ~pdata_13_13_ & n5842;
  assign n6380 = ~preset & ~n6379;
  assign n2752 = ~n6378 & n6380;
  assign n6382 = ~\[12185]  & ~n6026;
  assign n6383 = ~pdata_6_6_ & n6026;
  assign n6384 = ~preset & ~n6383;
  assign n2757 = ~n6382 & n6384;
  assign n6386 = ~\[12200]  & ~n6026;
  assign n6387 = ~pdata_15_15_ & n6026;
  assign n6388 = ~preset & ~n6387;
  assign n2762 = ~n6386 & n6388;
  assign n6390 = ppeakb_13_13_ & ~n2989;
  assign n6391 = \[13595]  & n2936;
  assign n6392 = ppeaka_13_13_ & ~n2950_1;
  assign n6393 = \[6620]  & n2939;
  assign n6394 = \[5210]  & n2955_1;
  assign n6395 = \[7325]  & n2964;
  assign n6396 = ~n6394 & ~n6395;
  assign n6397 = ~n6393 & n6396;
  assign n6398 = \[13670]  & n2952;
  assign n6399 = \[4460]  & n2961;
  assign n6400 = \[8570]  & n2916_1;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = ~n6398 & n6401;
  assign n6403 = \[14885]  & n2959;
  assign n6404 = n6402 & ~n6403;
  assign n6405 = n6397 & n6404;
  assign n6406 = ~n6392 & n6405;
  assign n6407 = n2907_1 & ~n6406;
  assign n6408 = ~n6391 & ~n6407;
  assign n6409 = \[14375]  & n2912_1;
  assign n6410 = \[15500]  & n2931;
  assign n6411 = ~n6409 & ~n6410;
  assign n6412 = n6408 & n6411;
  assign n2767 = n6390 | ~n6412;
  assign n6414 = n3966 & n4685;
  assign n6415 = \[12245]  & n4683;
  assign n2771 = n6414 | n6415;
  assign n6417 = ~\[12260]  & ~n5842;
  assign n6418 = ~pdata_14_14_ & n5842;
  assign n6419 = ~preset & ~n6418;
  assign n2776 = ~n6417 & n6419;
  assign n6421 = ~\[12275]  & ~n6026;
  assign n6422 = ~pdata_9_9_ & n6026;
  assign n6423 = ~preset & ~n6422;
  assign n2781 = ~n6421 & n6423;
  assign n6425 = \[11090]  & ~n2927;
  assign n6426 = ppeaki_13_13_ & n2985;
  assign n2786 = n6425 | n6426;
  assign n6428 = \[11585]  & ~n2927;
  assign n6429 = ppeaki_10_10_ & n2862_1;
  assign n6430 = ppeaki_6_6_ & ~n2861;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = n2907_1 & ~n6431;
  assign n6433 = ~n6428 & ~n6432;
  assign n6434 = ~preset & ppeaki_2_2_;
  assign n6435 = ~n2984 & n6434;
  assign n2790 = ~n6433 | n6435;
  assign n4428 = n3171 & n3257;
  assign n6438 = n3675 & n4428;
  assign n6439 = \[12335]  & n3178;
  assign n2794 = n6438 | n6439;
  assign n6441 = n3963 & n3572_1;
  assign n6442 = \[12350]  & n3225;
  assign n2799 = n6441 | n6442;
  assign n6444 = n3963 & ~n3646;
  assign n6445 = \[12365]  & n3225;
  assign n2804 = n6444 | n6445;
  assign n6447 = ~\[12380]  & ~n3717_1;
  assign n6448 = n3717_1 & ~n4104;
  assign n6449 = ~preset & ~n6448;
  assign n2809 = ~n6447 & n6449;
  assign n6451 = ~\[12395]  & ~n3717_1;
  assign n6452 = n3717_1 & ~n4111;
  assign n6453 = ~preset & ~n6452;
  assign n2814 = ~n6451 & n6453;
  assign n6455 = ~\[12410]  & ~n3720;
  assign n6456 = n3720 & n3866;
  assign n6457 = ~preset & ~n6456;
  assign n2819 = ~n6455 & n6457;
  assign n6459 = \[12425]  & n4097_1;
  assign n6460 = ~n4080 & n4091;
  assign n2824 = n6459 | n6460;
  assign n6462 = n4087_1 & n6333;
  assign n6463 = \[12440]  & n6335;
  assign n2829 = n6462 | n6463;
  assign n6465 = n4095 & n4685;
  assign n6466 = \[12455]  & n4683;
  assign n2834 = n6465 | n6466;
  assign n6468 = ~\[12470]  & ~n5842;
  assign n6469 = ~pdata_15_15_ & n5842;
  assign n6470 = ~preset & ~n6469;
  assign n2839 = ~n6468 & n6470;
  assign n6472 = ~\[12485]  & ~n6026;
  assign n6473 = ~pdata_8_8_ & n6026;
  assign n6474 = ~preset & ~n6473;
  assign n2844 = ~n6472 & n6474;
  assign n6476 = \[10820]  & ~n2927;
  assign n6477 = ppeaki_12_12_ & n2985;
  assign n2849 = n6476 | n6477;
  assign n6479 = ppeaki_3_3_ & n2985;
  assign n6480 = ppeaki_7_7_ & ~n2861;
  assign n6481 = ppeaki_11_11_ & n2862_1;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = n2907_1 & ~n6482;
  assign n6484 = \[11345]  & ~n2927;
  assign n6485 = ~n6483 & ~n6484;
  assign n2853 = n6479 | ~n6485;
  assign n6487 = \[12545]  & n3225;
  assign n6488 = pdata_4_4_ & n3963;
  assign n2857 = n6487 | n6488;
  assign n6490 = ~n4344_1 & n4428;
  assign n6491 = \[12560]  & n3178;
  assign n2862 = n6490 | n6491;
  assign n6493 = n3963 & n4605;
  assign n6494 = \[12575]  & n3225;
  assign n2867 = n6493 | n6494;
  assign n6496 = ~\[12590]  & ~n3231;
  assign n6497 = n3231 & n4626;
  assign n6498 = ~preset & ~n6497;
  assign n2872 = ~n6496 & n6498;
  assign n6500 = ~\[12605]  & ~n3717_1;
  assign n6501 = n3717_1 & ~n4672;
  assign n6502 = ~preset & ~n6501;
  assign n2877 = ~n6500 & n6502;
  assign n6504 = ~\[12620]  & ~n3717_1;
  assign n6505 = n3717_1 & n4392;
  assign n6506 = ~preset & ~n6505;
  assign n2882 = ~n6504 & n6506;
  assign n6508 = ~\[12635]  & ~n3720;
  assign n6509 = n3720 & ~n4399;
  assign n6510 = ~preset & ~n6509;
  assign n2887 = ~n6508 & n6510;
  assign n6512 = \[12650]  & n4097_1;
  assign n6513 = n4091 & ~n4692;
  assign n2892 = n6512 | n6513;
  assign n6515 = ~n3958_1 & n6333;
  assign n6516 = \[12665]  & n6335;
  assign n2897 = n6515 | n6516;
  assign n6518 = n4685 & ~n4955;
  assign n6519 = \[12680]  & n4683;
  assign n2902 = n6518 | n6519;
  assign n6521 = ~\[12695]  & ~n6026;
  assign n6522 = ~pdata_0_0_ & n6026;
  assign n6523 = ~preset & ~n6522;
  assign n2907 = ~n6521 & n6523;
  assign n6525 = ppeaki_11_11_ & n2985;
  assign n6526 = \[11600]  & ~n2927;
  assign n6527 = ppeaki_15_15_ & ~n2861;
  assign n6528 = n2907_1 & n6527;
  assign n6529 = ~n6526 & ~n6528;
  assign n2912 = n6525 | ~n6529;
  assign n6531 = ppeaki_0_0_ & n2985;
  assign n6532 = ppeaki_8_8_ & n2862_1;
  assign n6533 = ppeaki_4_4_ & ~n2861;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = n2907_1 & ~n6534;
  assign n6536 = \[12695]  & ~n2927;
  assign n6537 = ~n6535 & ~n6536;
  assign n2916 = n6531 | ~n6537;
  assign n6539 = \[12770]  & n3225;
  assign n6540 = pdata_14_14_ & n3963;
  assign n2920 = n6539 | n6540;
  assign n6542 = ~\[12800]  & ~n3265;
  assign n6543 = n3265 & ~n3564;
  assign n6544 = ~preset & ~n6543;
  assign n2925 = ~n6542 & n6544;
  assign n6546 = n3963 & ~n3667_1;
  assign n6547 = \[12815]  & n3225;
  assign n2930 = n6546 | n6547;
  assign n6549 = ~\[12830]  & ~n3231;
  assign n6550 = n3231 & ~n3675;
  assign n6551 = ~preset & ~n6550;
  assign n2935 = ~n6549 & n6551;
  assign n6553 = ~\[12845]  & ~n3717_1;
  assign n6554 = n3717_1 & ~n4095;
  assign n6555 = ~preset & ~n6554;
  assign n2940 = ~n6553 & n6555;
  assign n6557 = ~\[12860]  & ~n3717_1;
  assign n6558 = n3717_1 & n3958_1;
  assign n6559 = ~preset & ~n6558;
  assign n2945 = ~n6557 & n6559;
  assign n6561 = ~\[12875]  & ~n3720;
  assign n6562 = n3720 & ~n3966;
  assign n6563 = ~preset & ~n6562;
  assign n2950 = ~n6561 & n6563;
  assign n6565 = n4672 & n6333;
  assign n6566 = \[12890]  & n6335;
  assign n2955 = n6565 | n6566;
  assign n6568 = n4357 & n6333;
  assign n6569 = \[12905]  & n6335;
  assign n2960 = n6568 | n6569;
  assign n6571 = n4104 & n4685;
  assign n6572 = \[12920]  & n4683;
  assign n2965 = n6571 | n6572;
  assign n6574 = ~\[12935]  & ~n6026;
  assign n6575 = ~pdata_10_10_ & n6026;
  assign n6576 = ~preset & ~n6575;
  assign n2970 = ~n6574 & n6576;
  assign n6578 = ppeaki_10_10_ & n2985;
  assign n6579 = ppeaki_14_14_ & ~n2861;
  assign n6580 = n2907_1 & n6579;
  assign n6581 = \[12935]  & ~n2927;
  assign n6582 = ~n6580 & ~n6581;
  assign n2975 = n6578 | ~n6582;
  assign n6584 = ppeaki_1_1_ & n2985;
  assign n6585 = \[10805]  & ~n2927;
  assign n6586 = ppeaki_9_9_ & n2862_1;
  assign n6587 = ppeaki_5_5_ & ~n2861;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = n2907_1 & ~n6588;
  assign n6590 = ~n6585 & ~n6589;
  assign n2979 = n6584 | ~n6590;
  assign n6592 = ~\[13010]  & ~n3231;
  assign n6593 = ~pdata_8_8_ & n3231;
  assign n6594 = ~preset & ~n6593;
  assign n2983 = ~n6592 & n6594;
  assign n6596 = ~\[13025]  & ~n3265;
  assign n6597 = n3265 & n4298;
  assign n6598 = ~preset & ~n6597;
  assign n2988 = ~n6596 & n6598;
  assign n6600 = ~\[13040]  & ~n3265;
  assign n6601 = n3265 & ~n3653_1;
  assign n6602 = ~preset & ~n6601;
  assign n2993 = ~n6600 & n6602;
  assign n6604 = n3963 & n3556;
  assign n6605 = \[13055]  & n3225;
  assign n2998 = n6604 | n6605;
  assign n6607 = n3963 & ~n4326;
  assign n6608 = \[13070]  & n3225;
  assign n3003 = n6607 | n6608;
  assign n6610 = ~\[13085]  & ~n3231;
  assign n6611 = n3231 & n4344_1;
  assign n6612 = ~preset & ~n6611;
  assign n3008 = ~n6610 & n6612;
  assign n6614 = ~\[13100]  & ~n3717_1;
  assign n6615 = n3717_1 & n4955;
  assign n6616 = ~preset & ~n6615;
  assign n3013 = ~n6614 & n6616;
  assign n6618 = ~\[13115]  & ~n3717_1;
  assign n6619 = n3717_1 & n4365;
  assign n6620 = ~preset & ~n6619;
  assign n3018 = ~n6618 & n6620;
  assign n6622 = ~\[13130]  & ~n3720;
  assign n6623 = n3720 & ~n4095;
  assign n6624 = ~preset & ~n6623;
  assign n3023 = ~n6622 & n6624;
  assign n6626 = n4376 & n6333;
  assign n6627 = \[13160]  & n6335;
  assign n3028 = n6626 | n6627;
  assign n6629 = n4672 & n4685;
  assign n6630 = \[13175]  & n4683;
  assign n3033 = n6629 | n6630;
  assign n6632 = ppeakb_4_4_ & ~n2989;
  assign n6633 = \[12545]  & n3081_1;
  assign n6634 = ~n6632 & ~n6633;
  assign n6635 = \[14360]  & n2912_1;
  assign n6636 = \[14765]  & n2931;
  assign n6637 = \[5795]  & n2936;
  assign n6638 = \[14495]  & n2939;
  assign n6639 = \[7280]  & n2916_1;
  assign n6640 = ~n6638 & ~n6639;
  assign n6641 = \[9170]  & n2959;
  assign n6642 = \[8585]  & n2964;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = \[5840]  & n2961;
  assign n6645 = \[5195]  & n2955_1;
  assign n6646 = ~n6644 & ~n6645;
  assign n6647 = n6643 & n6646;
  assign n6648 = n6640 & n6647;
  assign n6649 = n2907_1 & ~n6648;
  assign n6650 = ~n6637 & ~n6649;
  assign n6651 = ~n6636 & n6650;
  assign n6652 = ~n6635 & n6651;
  assign n6653 = ~n2906 & ~n6652;
  assign n6654 = ppeaka_4_4_ & n4124;
  assign n6655 = ~n6653 & ~n6654;
  assign n3038 = ~n6634 | ~n6655;
  assign n6657 = ppeakp_9_9_ & ~n3035;
  assign n6658 = ppeaka_9_9_ & ppeakb_9_9_;
  assign n6659 = n2912_1 & ~n6658;
  assign n6660 = \[16040]  & n2936;
  assign n6661 = \[11270]  & n3044;
  assign n6662 = \[13265]  & n3020;
  assign n6663 = \[5825]  & n2961;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = \[9125]  & n3030;
  assign n6666 = \[9905]  & n2964;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = n6664 & n6667;
  assign n6669 = ~n6661 & n6668;
  assign n6670 = n2907_1 & ~n6669;
  assign n6671 = ~n6660 & ~n6670;
  assign n6672 = \[15770]  & n3024;
  assign n6673 = n6671 & ~n6672;
  assign n6674 = ~n6659 & n6673;
  assign n6675 = ~n6657 & n6674;
  assign n6676 = ~n2906 & ~n6675;
  assign n6677 = \[5720]  & n4453_1;
  assign n6678 = ppeakb_9_9_ & n4451;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = ~n6676 & n6679;
  assign n6681 = ppeaka_9_9_ & ~n3042_1;
  assign n6682 = ppeaka_10_10_ & n2975_1;
  assign n6683 = ~n6681 & ~n6682;
  assign n3042 = ~n6680 | ~n6683;
  assign n6685 = ~\[13220]  & ~n3162;
  assign n6686 = ~pdata_3_3_ & n3162;
  assign n6687 = ~preset & ~n6686;
  assign n3046 = ~n6685 & n6687;
  assign n6689 = ~\[13235]  & ~n3162;
  assign n6690 = ~pdata_14_14_ & n3162;
  assign n6691 = ~preset & ~n6690;
  assign n3051 = ~n6689 & n6691;
  assign n6693 = ~pdata_14_14_ & n3175;
  assign n6694 = ~\[13250]  & ~n3175;
  assign n6695 = ~preset & ~n6694;
  assign n3056 = ~n6693 & n6695;
  assign n6697 = ~\[13265]  & ~n3181;
  assign n6698 = ~pdata_9_9_ & n3181;
  assign n6699 = ~preset & ~n6698;
  assign n3061 = ~n6697 & n6699;
  assign n6701 = \[13280]  & n3194_1;
  assign n3066 = n4559 | n6701;
  assign n6703 = ~\[13295]  & ~n3218;
  assign n6704 = ~pdata_1_1_ & n3218;
  assign n6705 = ~preset & ~n6704;
  assign n3071 = ~n6703 & n6705;
  assign n6707 = \[13310]  & n3225;
  assign n6708 = pdata_1_1_ & n3963;
  assign n3076 = n6707 | n6708;
  assign n6710 = \[13325]  & n3225;
  assign n6711 = pdata_12_12_ & n3963;
  assign n3081 = n6710 | n6711;
  assign n6713 = ~\[13340]  & ~n3231;
  assign n6714 = ~pdata_7_7_ & n3231;
  assign n6715 = ~preset & ~n6714;
  assign n3086 = ~n6713 & n6715;
  assign n6717 = n4605 & n4428;
  assign n6718 = \[13355]  & n3178;
  assign n3091 = n6717 | n6718;
  assign n6720 = ~n4326 & n4428;
  assign n6721 = \[13370]  & n3178;
  assign n3096 = n6720 | n6721;
  assign n6723 = ~\[13385]  & ~n3265;
  assign n6724 = n3265 & n4626;
  assign n6725 = ~preset & ~n6724;
  assign n3101 = ~n6723 & n6725;
  assign n6727 = n3963 & ~n4298;
  assign n6728 = \[13400]  & n3225;
  assign n3106 = n6727 | n6728;
  assign n6730 = n3963 & ~n3549;
  assign n6731 = \[13415]  & n3225;
  assign n3111 = n6730 | n6731;
  assign n6733 = ~\[13430]  & ~n3231;
  assign n6734 = n3231 & ~n3556;
  assign n6735 = ~preset & ~n6734;
  assign n3116 = ~n6733 & n6735;
  assign n6737 = ~\[13445]  & ~n3691;
  assign n6738 = n3691 & n4692;
  assign n6739 = ~preset & ~n6738;
  assign n3121 = ~n6737 & n6739;
  assign n6741 = ~\[13460]  & ~n3717_1;
  assign n6742 = n3717_1 & ~n4376;
  assign n6743 = ~preset & ~n6742;
  assign n3126 = ~n6741 & n6743;
  assign n6745 = ~\[13475]  & ~n3720;
  assign n6746 = n3720 & n4955;
  assign n6747 = ~preset & ~n6746;
  assign n3131 = ~n6745 & n6747;
  assign n6749 = \[13490]  & n4097_1;
  assign n6750 = n4091 & ~n4365;
  assign n3136 = n6749 | n6750;
  assign n6752 = n4399 & n6333;
  assign n6753 = \[13505]  & n6335;
  assign n3141 = n6752 | n6753;
  assign n6755 = ppeakb_5_5_ & ~n2989;
  assign n6756 = \[5240]  & n3081_1;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = \[13955]  & n2912_1;
  assign n6759 = \[8330]  & n2931;
  assign n6760 = \[6485]  & n2936;
  assign n6761 = \[9245]  & n2964;
  assign n6762 = \[5885]  & n2955_1;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = \[7235]  & n2959;
  assign n6765 = \[7910]  & n2916_1;
  assign n6766 = ~n6764 & ~n6765;
  assign n6767 = \[14075]  & n2939;
  assign n6768 = \[7790]  & n2961;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = n6766 & n6769;
  assign n6771 = n6763 & n6770;
  assign n6772 = n2907_1 & ~n6771;
  assign n6773 = ~n6760 & ~n6772;
  assign n6774 = ~n6759 & n6773;
  assign n6775 = ~n6758 & n6774;
  assign n6776 = ~n2906 & ~n6775;
  assign n6777 = ppeaka_5_5_ & n4124;
  assign n6778 = ~n6776 & ~n6777;
  assign n3146 = ~n6757 | ~n6778;
  assign n6780 = \[13550]  & ~n3065;
  assign n6781 = \[9890]  & n3068;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = \[10355]  & n2931;
  assign n6784 = \[6650]  & n2917;
  assign n6785 = ~n6783 & ~n6784;
  assign n3150 = ~n6782 | ~n6785;
  assign n6787 = ppeakp_6_6_ & ~n3147;
  assign n6788 = ppeaka_6_6_ & ~n3156;
  assign n6789 = \[9575]  & n3021;
  assign n6790 = ~n6788 & ~n6789;
  assign n6791 = ~n6787 & n6790;
  assign n6792 = \[14705]  & n3095;
  assign n6793 = ppeakb_6_6_ & n2917;
  assign n6794 = \[10085]  & ~n2927;
  assign n6795 = ~n6793 & ~n6794;
  assign n6796 = ~n6792 & n6795;
  assign n3155 = ~n6791 | ~n6796;
  assign n6798 = ~\[13580]  & ~n3162;
  assign n6799 = ~pdata_15_15_ & n3162;
  assign n6800 = ~preset & ~n6799;
  assign n3159 = ~n6798 & n6800;
  assign n6802 = ~pdata_13_13_ & n3175;
  assign n6803 = ~\[13595]  & ~n3175;
  assign n6804 = ~preset & ~n6803;
  assign n3164 = ~n6802 & n6804;
  assign n6806 = ~\[13610]  & ~n3181;
  assign n6807 = ~pdata_10_10_ & n3181;
  assign n6808 = ~preset & ~n6807;
  assign n3169 = ~n6806 & n6808;
  assign n6810 = \[13625]  & n3194_1;
  assign n3174 = n4849 | n6810;
  assign n6812 = ~\[13640]  & ~n3218;
  assign n6813 = ~pdata_2_2_ & n3218;
  assign n6814 = ~preset & ~n6813;
  assign n3179 = ~n6812 & n6814;
  assign n6816 = \[13655]  & n3225;
  assign n6817 = pdata_0_0_ & n3963;
  assign n3184 = n6816 | n6817;
  assign n6819 = \[13670]  & n3225;
  assign n6820 = pdata_13_13_ & n3963;
  assign n3189 = n6819 | n6820;
  assign n6822 = ~\[13685]  & ~n3231;
  assign n6823 = ~pdata_6_6_ & n3231;
  assign n6824 = ~preset & ~n6823;
  assign n3194 = ~n6822 & n6824;
  assign n6826 = n4161 & n3556;
  assign n6827 = \[13700]  & n3312;
  assign n3199 = n6826 | n6827;
  assign n6829 = n3660 & n4428;
  assign n6830 = \[13715]  & n3178;
  assign n3204 = n6829 | n6830;
  assign n6832 = ~n3646 & n4428;
  assign n6833 = \[13730]  & n3178;
  assign n3209 = n6832 | n6833;
  assign n6835 = ~\[13745]  & ~n3265;
  assign n6836 = n3265 & ~n3675;
  assign n6837 = ~preset & ~n6836;
  assign n3214 = ~n6835 & n6837;
  assign n6839 = n3963 & n3541;
  assign n6840 = \[13775]  & n3225;
  assign n3219 = n6839 | n6840;
  assign n6842 = ~\[13790]  & ~n3231;
  assign n6843 = n3231 & ~n3572_1;
  assign n6844 = ~preset & ~n6843;
  assign n3224 = ~n6842 & n6844;
  assign n6846 = ~\[13805]  & ~n3691;
  assign n6847 = n3691 & n4392;
  assign n6848 = ~preset & ~n6847;
  assign n3229 = ~n6846 & n6848;
  assign n6850 = ~\[13820]  & ~n3717_1;
  assign n6851 = n3717_1 & ~n4087_1;
  assign n6852 = ~preset & ~n6851;
  assign n3234 = ~n6850 & n6852;
  assign n6854 = ~\[13835]  & ~n3720;
  assign n6855 = n3720 & ~n4104;
  assign n6856 = ~preset & ~n6855;
  assign n3239 = ~n6854 & n6856;
  assign n6858 = ~n3958_1 & n4091;
  assign n6859 = \[13850]  & n4097_1;
  assign n3244 = n6858 | n6859;
  assign n6861 = ~n3866 & n6333;
  assign n6862 = \[13865]  & n6335;
  assign n3249 = n6861 | n6862;
  assign n6864 = \[13880]  & n6335;
  assign n6865 = ~n4080 & n6333;
  assign n3254 = n6864 | n6865;
  assign n6867 = ~\[13895]  & ~n2843;
  assign n6868 = ~pdata_8_8_ & n2843;
  assign n6869 = ~preset & ~n6868;
  assign n3259 = ~n6867 & n6869;
  assign n6871 = ppeakb_11_11_ & ppeaka_11_11_;
  assign n6872 = n2912_1 & ~n6871;
  assign n6873 = ~n5558 & ~n6872;
  assign n6874 = \[15335]  & n2936;
  assign n6875 = \[5120]  & n3021;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = ppeakp_11_11_ & ~n3035;
  assign n6878 = n6876 & ~n6877;
  assign n6879 = n6873 & n6878;
  assign n6880 = ~n2906 & ~n6879;
  assign n6881 = ppeaka_12_12_ & n2975_1;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ppeaka_11_11_ & ~n3042_1;
  assign n6884 = ppeakb_11_11_ & ~n3050;
  assign n6885 = \[7820]  & n3030;
  assign n6886 = \[7145]  & n2961;
  assign n6887 = \[11735]  & n3044;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = ~n6885 & n6888;
  assign n6890 = \[4295]  & ~n3047;
  assign n6891 = \[9650]  & n2964;
  assign n6892 = ~n6890 & ~n6891;
  assign n6893 = n6889 & n6892;
  assign n6894 = ~n6884 & n6893;
  assign n6895 = n2907_1 & ~n6894;
  assign n6896 = ~n6883 & ~n6895;
  assign n3264 = ~n6882 | ~n6896;
  assign n6898 = ppeakp_0_0_ & ~n3035;
  assign n6899 = ppeaka_0_0_ & ~n3042_1;
  assign n6900 = ppeakb_0_0_ & ppeaka_0_0_;
  assign n6901 = n2912_1 & ~n6900;
  assign n6902 = \[14840]  & n2961;
  assign n6903 = \[4310]  & ~n3047;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = \[9110]  & n3030;
  assign n6906 = \[13970]  & n3020;
  assign n6907 = ppeakb_0_0_ & ~n3050;
  assign n6908 = ~n6906 & ~n6907;
  assign n6909 = ~n6905 & n6908;
  assign n6910 = \[11255]  & n3044;
  assign n6911 = \[11480]  & n2964;
  assign n6912 = ~n6910 & ~n6911;
  assign n6913 = n6909 & n6912;
  assign n6914 = n6904 & n6913;
  assign n6915 = n2907_1 & ~n6914;
  assign n6916 = ppeaka_1_1_ & n2975_1;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = \[8240]  & n3024;
  assign n6919 = \[16025]  & n2936;
  assign n6920 = ~n6918 & ~n6919;
  assign n6921 = n6917 & n6920;
  assign n6922 = ~n6901 & n6921;
  assign n6923 = ~n6899 & n6922;
  assign n3268 = n6898 | ~n6923;
  assign n6925 = ppeakp_5_5_ & ~n3147;
  assign n6926 = ppeaka_5_5_ & ~n3156;
  assign n6927 = \[11660]  & n3021;
  assign n6928 = ~n6926 & ~n6927;
  assign n6929 = ~n6925 & n6928;
  assign n6930 = \[15080]  & n3095;
  assign n6931 = ppeakb_5_5_ & n2917;
  assign n6932 = \[8840]  & ~n2927;
  assign n6933 = ~n6931 & ~n6932;
  assign n6934 = ~n6930 & n6933;
  assign n3272 = ~n6929 | ~n6934;
  assign n6936 = ~\[13955]  & ~n3162;
  assign n6937 = ~pdata_5_5_ & n3162;
  assign n6938 = ~preset & ~n6937;
  assign n3276 = ~n6936 & n6938;
  assign n6940 = ~\[13970]  & ~n3181;
  assign n6941 = ~pdata_0_0_ & n3181;
  assign n6942 = ~preset & ~n6941;
  assign n3281 = ~n6940 & n6942;
  assign n6944 = ~\[13985]  & ~n3181;
  assign n6945 = ~pdata_7_7_ & n3181;
  assign n6946 = ~preset & ~n6945;
  assign n3286 = ~n6944 & n6946;
  assign n6948 = \[14000]  & n3194_1;
  assign n3291 = n3197 | n6948;
  assign n6950 = ~\[14015]  & ~n3203;
  assign n6951 = ~pdata_13_13_ & n3203;
  assign n6952 = ~preset & ~n6951;
  assign n3296 = ~n6950 & n6952;
  assign n6954 = ~pdata_8_8_ & n3208;
  assign n6955 = ~\[14030]  & ~n3208;
  assign n6956 = ~preset & ~n6955;
  assign n3301 = ~n6954 & n6956;
  assign n6958 = \[14045]  & n3225;
  assign n6959 = pdata_3_3_ & n3963;
  assign n3306 = n6958 | n6959;
  assign n6961 = \[14060]  & n3225;
  assign n6962 = pdata_10_10_ & n3963;
  assign n3311 = n6961 | n6962;
  assign n6964 = ~\[14075]  & ~n3231;
  assign n6965 = ~pdata_5_5_ & n3231;
  assign n6966 = ~preset & ~n6965;
  assign n3316 = ~n6964 & n6966;
  assign n6968 = ~\[14090]  & ~n3249_1;
  assign n6969 = ~pdata_11_11_ & n3249_1;
  assign n6970 = ~preset & ~n6969;
  assign n3321 = ~n6968 & n6970;
  assign n6972 = n3556 & n4428;
  assign n6973 = \[14105]  & n3178;
  assign n3326 = n6972 | n6973;
  assign n6975 = n3541 & n4428;
  assign n6976 = \[14120]  & n3178;
  assign n3331 = n6975 | n6976;
  assign n6978 = ~\[14135]  & ~n3265;
  assign n6979 = n3265 & n4344_1;
  assign n6980 = ~preset & ~n6979;
  assign n3336 = ~n6978 & n6980;
  assign n6982 = n3963 & n3660;
  assign n6983 = \[14150]  & n3225;
  assign n3341 = n6982 | n6983;
  assign n6985 = n3963 & n3653_1;
  assign n6986 = \[14165]  & n3225;
  assign n3346 = n6985 | n6986;
  assign n6988 = ~\[14180]  & ~n3231;
  assign n6989 = n3231 & ~n4605;
  assign n6990 = ~preset & ~n6989;
  assign n3351 = ~n6988 & n6990;
  assign n6992 = ~\[14210]  & ~n3717_1;
  assign n6993 = n3717_1 & n3866;
  assign n6994 = ~preset & ~n6993;
  assign n3356 = ~n6992 & n6994;
  assign n6996 = ~\[14225]  & ~n3720;
  assign n6997 = n3720 & ~n4672;
  assign n6998 = ~preset & ~n6997;
  assign n3361 = ~n6996 & n6998;
  assign n7000 = \[14240]  & n4097_1;
  assign n7001 = n4091 & ~n4392;
  assign n3366 = n7000 | n7001;
  assign n7003 = n4095 & n6333;
  assign n7004 = \[14255]  & n6335;
  assign n3371 = n7003 | n7004;
  assign n7006 = ~n4692 & n6333;
  assign n7007 = \[14270]  & n6335;
  assign n3376 = n7006 | n7007;
  assign n7009 = ~\[14285]  & ~n2843;
  assign n7010 = ~pdata_7_7_ & n2843;
  assign n7011 = ~preset & ~n7010;
  assign n3381 = ~n7009 & n7011;
  assign n7013 = ppeakb_3_3_ & ~n2989;
  assign n7014 = \[6530]  & n2961;
  assign n7015 = \[14045]  & n2952;
  assign n7016 = \[14915]  & n2939;
  assign n7017 = \[7940]  & n2964;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = \[4490]  & n2955_1;
  assign n7020 = n7018 & ~n7019;
  assign n7021 = ~n7015 & n7020;
  assign n7022 = ppeaka_3_3_ & ~n2950_1;
  assign n7023 = \[8510]  & n2959;
  assign n7024 = \[9215]  & n2916_1;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = ~n7022 & n7025;
  assign n7027 = n7021 & n7026;
  assign n7028 = ~n7014 & n7027;
  assign n7029 = n2907_1 & ~n7028;
  assign n7030 = \[7760]  & n2936;
  assign n7031 = \[13220]  & n2912_1;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = \[15860]  & n2931;
  assign n7034 = n7032 & ~n7033;
  assign n7035 = ~n7029 & n7034;
  assign n3386 = n7013 | ~n7035;
  assign n7037 = ppeakp_10_10_ & ~n3035;
  assign n7038 = ppeaka_10_10_ & ~n3042_1;
  assign n7039 = ppeakb_10_10_ & ppeaka_10_10_;
  assign n7040 = n2912_1 & ~n7039;
  assign n7041 = ppeaka_11_11_ & n2975_1;
  assign n7042 = \[13850]  & n3024;
  assign n7043 = \[14960]  & n2936;
  assign n7044 = \[11705]  & n2964;
  assign n7045 = ppeakb_10_10_ & ~n3050;
  assign n7046 = \[11015]  & n3044;
  assign n7047 = \[5015]  & ~n3047;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n7045 & n7048;
  assign n7050 = \[13610]  & n3020;
  assign n7051 = \[8465]  & n3030;
  assign n7052 = \[6515]  & n2961;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = ~n7050 & n7053;
  assign n7055 = n7049 & n7054;
  assign n7056 = ~n7044 & n7055;
  assign n7057 = n2907_1 & ~n7056;
  assign n7058 = ~n7043 & ~n7057;
  assign n7059 = ~n7042 & n7058;
  assign n7060 = ~n7041 & n7059;
  assign n7061 = ~n7040 & n7060;
  assign n7062 = ~n7038 & n7061;
  assign n3390 = n7037 | ~n7062;
  assign n7064 = ppeakp_1_1_ & ~n3035;
  assign n7065 = ppeaka_1_1_ & ~n3042_1;
  assign n7066 = ppeakb_1_1_ & ppeaka_1_1_;
  assign n7067 = n2912_1 & ~n7066;
  assign n7068 = \[7175]  & n3030;
  assign n7069 = \[14420]  & n2961;
  assign n7070 = ~n7068 & ~n7069;
  assign n7071 = \[11495]  & n3044;
  assign n7072 = \[4925]  & n2964;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = ppeakb_1_1_ & ~n3050;
  assign n7075 = \[5030]  & ~n3047;
  assign n7076 = ~n7074 & ~n7075;
  assign n7077 = n7073 & n7076;
  assign n7078 = n7070 & n7077;
  assign n7079 = n2907_1 & ~n7078;
  assign n7080 = \[4400]  & n3021;
  assign n7081 = ~n5009 & ~n7080;
  assign n7082 = ~n7079 & n7081;
  assign n7083 = \[15680]  & n2936;
  assign n7084 = ppeaka_2_2_ & n2975_1;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = n7082 & n7085;
  assign n7087 = ~n7067 & n7086;
  assign n7088 = ~n7065 & n7087;
  assign n3394 = n7064 | ~n7088;
  assign n7090 = ppeakp_4_4_ & ~n3147;
  assign n7091 = ppeaka_4_4_ & ~n3156;
  assign n7092 = \[11435]  & n3021;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = ~n7090 & n7093;
  assign n7095 = \[15440]  & n3095;
  assign n7096 = ppeakb_4_4_ & n2917;
  assign n7097 = \[9515]  & ~n2927;
  assign n7098 = ~n7096 & ~n7097;
  assign n7099 = ~n7095 & n7098;
  assign n3398 = ~n7094 | ~n7099;
  assign n7101 = ~\[14360]  & ~n3162;
  assign n7102 = ~pdata_4_4_ & n3162;
  assign n7103 = ~preset & ~n7102;
  assign n3402 = ~n7101 & n7103;
  assign n7105 = ~\[14375]  & ~n3162;
  assign n7106 = ~pdata_13_13_ & n3162;
  assign n7107 = ~preset & ~n7106;
  assign n3407 = ~n7105 & n7107;
  assign n7109 = ~pdata_15_15_ & n3175;
  assign n7110 = ~\[14390]  & ~n3175;
  assign n7111 = ~preset & ~n7110;
  assign n3412 = ~n7109 & n7111;
  assign n7113 = ~\[14405]  & ~n3181;
  assign n7114 = ~pdata_8_8_ & n3181;
  assign n7115 = ~preset & ~n7114;
  assign n3417 = ~n7113 & n7115;
  assign n7117 = \[14420]  & n3194_1;
  assign n3422 = n4254 | n7117;
  assign n7119 = ~\[14435]  & ~n3203;
  assign n7120 = ~pdata_14_14_ & n3203;
  assign n7121 = ~preset & ~n7120;
  assign n3427 = ~n7119 & n7121;
  assign n7123 = ~pdata_7_7_ & n3208;
  assign n7124 = ~\[14450]  & ~n3208;
  assign n7125 = ~preset & ~n7124;
  assign n3432 = ~n7123 & n7125;
  assign n7127 = \[14465]  & n3225;
  assign n7128 = pdata_2_2_ & n3963;
  assign n3437 = n7127 | n7128;
  assign n7130 = \[14480]  & n3225;
  assign n7131 = pdata_11_11_ & n3963;
  assign n3442 = n7130 | n7131;
  assign n7133 = ~\[14495]  & ~n3231;
  assign n7134 = ~pdata_4_4_ & n3231;
  assign n7135 = ~preset & ~n7134;
  assign n3447 = ~n7133 & n7135;
  assign n7137 = ~\[14510]  & ~n3249_1;
  assign n7138 = ~pdata_1_1_ & n3249_1;
  assign n7139 = ~preset & ~n7138;
  assign n3452 = ~n7137 & n7139;
  assign n7141 = n3572_1 & n4428;
  assign n7142 = \[14525]  & n3178;
  assign n3457 = n7141 | n7142;
  assign n7144 = ~n3667_1 & n4428;
  assign n7145 = \[14540]  & n3178;
  assign n3462 = n7144 | n7145;
  assign n7147 = ~\[14555]  & ~n3265;
  assign n7148 = n3265 & ~n3556;
  assign n7149 = ~preset & ~n7148;
  assign n3467 = ~n7147 & n7149;
  assign n7151 = n3963 & ~n3310;
  assign n7152 = \[14570]  & n3225;
  assign n3472 = n7151 | n7152;
  assign n7154 = n3963 & n3564;
  assign n7155 = \[14585]  & n3225;
  assign n3477 = n7154 | n7155;
  assign n7157 = ~\[14600]  & ~n3231;
  assign n7158 = n3231 & ~n3660;
  assign n7159 = ~preset & ~n7158;
  assign n3482 = ~n7157 & n7159;
  assign n7161 = ~\[14615]  & ~n3691;
  assign n7162 = n3691 & n4080;
  assign n7163 = ~preset & ~n7162;
  assign n3487 = ~n7161 & n7163;
  assign n7165 = ~\[14630]  & ~n3717_1;
  assign n7166 = n3717_1 & ~n4357;
  assign n7167 = ~preset & ~n7166;
  assign n3492 = ~n7165 & n7167;
  assign n7169 = \[14660]  & n4097_1;
  assign n7170 = n4091 & n4111;
  assign n3497 = n7169 | n7170;
  assign n7172 = n3966 & n6333;
  assign n7173 = \[14675]  & n6335;
  assign n3502 = n7172 | n7173;
  assign n7175 = ~n4392 & n6333;
  assign n7176 = \[14690]  & n6335;
  assign n3507 = n7175 | n7176;
  assign n7178 = ~\[14705]  & ~n2843;
  assign n7179 = ~pdata_6_6_ & n2843;
  assign n7180 = ~preset & ~n7179;
  assign n3512 = ~n7178 & n7180;
  assign n7182 = \[6410]  & n2931;
  assign n7183 = ppeakb_8_8_ & ~n2989;
  assign n7184 = \[5810]  & n2936;
  assign n7185 = \[9050]  & n2912_1;
  assign n7186 = ppeaka_8_8_ & ~n2950_1;
  assign n7187 = \[14900]  & n2952;
  assign n7188 = \[13010]  & n2939;
  assign n7189 = \[6005]  & n2964;
  assign n7190 = ~n7188 & ~n7189;
  assign n7191 = ~n7187 & n7190;
  assign n7192 = \[6665]  & n2916_1;
  assign n7193 = \[8435]  & n2961;
  assign n7194 = \[14030]  & n2955_1;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = ~n7192 & n7195;
  assign n7197 = \[6605]  & n2959;
  assign n7198 = n7196 & ~n7197;
  assign n7199 = n7191 & n7198;
  assign n7200 = ~n7186 & n7199;
  assign n7201 = n2907_1 & ~n7200;
  assign n7202 = ~n7185 & ~n7201;
  assign n7203 = ~n7184 & n7202;
  assign n7204 = ~n7183 & n7203;
  assign n3517 = n7182 | ~n7204;
  assign n7206 = ppeakb_13_13_ & ppeaka_13_13_;
  assign n7207 = n2912_1 & ~n7206;
  assign n7208 = ~n5208 & ~n7207;
  assign n7209 = \[14540]  & n2936;
  assign n7210 = \[15920]  & n3021;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = ppeakp_13_13_ & ~n3035;
  assign n7213 = n7211 & ~n7212;
  assign n7214 = n7208 & n7213;
  assign n7215 = ~n2906 & ~n7214;
  assign n7216 = ppeaka_14_14_ & n2975_1;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = ppeaka_13_13_ & ~n3042_1;
  assign n7219 = \[15500]  & ~n3047;
  assign n7220 = \[10190]  & n3044;
  assign n7221 = \[8420]  & n2961;
  assign n7222 = \[14015]  & n3030;
  assign n7223 = ~n7221 & ~n7222;
  assign n7224 = ~n7220 & n7223;
  assign n7225 = ppeakb_13_13_ & ~n3050;
  assign n7226 = \[5645]  & n2964;
  assign n7227 = ~n7225 & ~n7226;
  assign n7228 = n7224 & n7227;
  assign n7229 = ~n7219 & n7228;
  assign n7230 = n2907_1 & ~n7229;
  assign n7231 = ~n7218 & ~n7230;
  assign n3521 = ~n7217 | ~n7231;
  assign n7233 = ppeakp_2_2_ & ~n3035;
  assign n7234 = ppeaka_2_2_ & ~n3042_1;
  assign n7235 = \[13715]  & n2936;
  assign n7236 = ppeakb_2_2_ & ppeaka_2_2_;
  assign n7237 = n2912_1 & ~n7236;
  assign n7238 = ppeaka_3_3_ & n2975_1;
  assign n7239 = \[9635]  & n2964;
  assign n7240 = \[15515]  & ~n3047;
  assign n7241 = ~n7239 & ~n7240;
  assign n7242 = \[7805]  & n3030;
  assign n7243 = \[5105]  & n3020;
  assign n7244 = ppeakb_2_2_ & ~n3050;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n7242 & n7245;
  assign n7247 = \[11720]  & n3044;
  assign n7248 = \[14000]  & n2961;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = n7246 & n7249;
  assign n7251 = n7241 & n7250;
  assign n7252 = n2907_1 & ~n7251;
  assign n7253 = ~n5588 & ~n7252;
  assign n7254 = ~n7238 & n7253;
  assign n7255 = ~n7237 & n7254;
  assign n7256 = ~n7235 & n7255;
  assign n7257 = ~n7234 & n7256;
  assign n3525 = n7233 | ~n7257;
  assign n7259 = \[14765]  & ~n3065;
  assign n7260 = \[5270]  & n2917;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = \[12875]  & n2931;
  assign n7263 = \[9875]  & n3068;
  assign n7264 = ~n7262 & ~n7263;
  assign n3529 = ~n7261 | ~n7264;
  assign n7266 = ppeaks_9_9_ & ~n3090;
  assign n7267 = \[14165]  & n3081_1;
  assign n7268 = \[13820]  & n2931;
  assign n7269 = \[13040]  & n2936;
  assign n7270 = \[8780]  & n2917;
  assign n7271 = \[10685]  & n3021;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = \[7970]  & n2912_1;
  assign n7274 = n7272 & ~n7273;
  assign n7275 = ~n7269 & n7274;
  assign n7276 = \[11045]  & n3095;
  assign n7277 = ~n6672 & ~n7276;
  assign n7278 = \[9590]  & n3068;
  assign n7279 = \[12440]  & n2949;
  assign n7280 = \[9470]  & n2964;
  assign n7281 = \[4745]  & n2959;
  assign n7282 = \[5405]  & n2961;
  assign n7283 = \[11135]  & n2955_1;
  assign n7284 = ~n7282 & ~n7283;
  assign n7285 = ~n7281 & n7284;
  assign n7286 = ~n7280 & n7285;
  assign n7287 = ~n7279 & n7286;
  assign n7288 = \[5465]  & n2939;
  assign n7289 = n7287 & ~n7288;
  assign n7290 = n2907_1 & ~n7289;
  assign n7291 = ~n7278 & ~n7290;
  assign n7292 = n7277 & n7291;
  assign n7293 = n7275 & n7292;
  assign n7294 = ~n7268 & n7293;
  assign n7295 = ~n2906 & ~n7294;
  assign n7296 = ~n7267 & ~n7295;
  assign n3534 = n7266 | ~n7296;
  assign n7298 = ppeakp_14_14_ & ~n3147;
  assign n7299 = ppeaka_14_14_ & ~n3156;
  assign n7300 = \[11675]  & n3021;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~n7298 & n7301;
  assign n7303 = \[11525]  & n3095;
  assign n7304 = ppeakb_14_14_ & n2917;
  assign n7305 = \[7580]  & ~n2927;
  assign n7306 = ~n7304 & ~n7305;
  assign n7307 = ~n7303 & n7306;
  assign n3538 = ~n7302 | ~n7307;
  assign n7309 = ~pdata_10_10_ & n3175;
  assign n7310 = ~\[14810]  & ~n3175;
  assign n7311 = ~preset & ~n7310;
  assign n3542 = ~n7309 & n7311;
  assign n7313 = ~\[14825]  & ~n3181;
  assign n7314 = ~pdata_5_5_ & n3181;
  assign n7315 = ~preset & ~n7314;
  assign n3547 = ~n7313 & n7315;
  assign n7317 = pdata_0_0_ & n3192;
  assign n7318 = \[14840]  & n3194_1;
  assign n3552 = n7317 | n7318;
  assign n7320 = \[14855]  & n3194_1;
  assign n3557 = n4556 | n7320;
  assign n7322 = ~\[14870]  & ~n3203;
  assign n7323 = ~pdata_4_4_ & n3203;
  assign n7324 = ~preset & ~n7323;
  assign n3562 = ~n7322 & n7324;
  assign n7326 = ~\[14885]  & ~n3218;
  assign n7327 = ~pdata_13_13_ & n3218;
  assign n7328 = ~preset & ~n7327;
  assign n3567 = ~n7326 & n7328;
  assign n7330 = pdata_8_8_ & n3963;
  assign n7331 = \[14900]  & n3225;
  assign n3572 = n7330 | n7331;
  assign n7333 = ~\[14915]  & ~n3231;
  assign n7334 = ~pdata_3_3_ & n3231;
  assign n7335 = ~preset & ~n7334;
  assign n3577 = ~n7333 & n7335;
  assign n7337 = \[14930]  & n3240;
  assign n3582 = n4589 | n7337;
  assign n7339 = n3564 & n4428;
  assign n7340 = \[14960]  & n3178;
  assign n3587 = n7339 | n7340;
  assign n7342 = ~\[14975]  & ~n3265;
  assign n7343 = n3265 & ~n3572_1;
  assign n7344 = ~preset & ~n7343;
  assign n3592 = ~n7342 & n7344;
  assign n7346 = ~\[14990]  & ~n3218;
  assign n7347 = n3218 & n3667_1;
  assign n7348 = ~preset & ~n7347;
  assign n3597 = ~n7346 & n7348;
  assign n7350 = n3963 & n3675;
  assign n7351 = \[15005]  & n3225;
  assign n3602 = n7350 | n7351;
  assign n7353 = ~\[15020]  & ~n3231;
  assign n7354 = n3231 & n3310;
  assign n7355 = ~preset & ~n7354;
  assign n3607 = ~n7353 & n7355;
  assign n7357 = ~\[15035]  & ~n3717_1;
  assign n7358 = n3717_1 & ~n3966;
  assign n7359 = ~preset & ~n7358;
  assign n3612 = ~n7357 & n7359;
  assign n7361 = ~\[15050]  & ~n3717_1;
  assign n7362 = n3717_1 & n4080;
  assign n7363 = ~preset & ~n7362;
  assign n3617 = ~n7361 & n7363;
  assign n7365 = n4111 & n6333;
  assign n7366 = \[15065]  & n6335;
  assign n3622 = n7365 | n7366;
  assign n7368 = ~\[15080]  & ~n2843;
  assign n7369 = ~pdata_5_5_ & n2843;
  assign n7370 = ~preset & ~n7369;
  assign n3627 = ~n7368 & n7370;
  assign n7372 = ppeakb_9_9_ & ~n2989;
  assign n7373 = \[5720]  & n2931;
  assign n7374 = \[15185]  & n2936;
  assign n7375 = \[8390]  & n2912_1;
  assign n7376 = ppeaka_9_9_ & ~n2950_1;
  assign n7377 = \[4520]  & n2959;
  assign n7378 = \[15275]  & n2952;
  assign n7379 = ~n7377 & ~n7378;
  assign n7380 = \[6680]  & n2964;
  assign n7381 = \[14855]  & n2961;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = \[7850]  & n2955_1;
  assign n7384 = n7382 & ~n7383;
  assign n7385 = \[16010]  & n2939;
  assign n7386 = \[5990]  & n2916_1;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = n7384 & n7387;
  assign n7389 = n7379 & n7388;
  assign n7390 = ~n7376 & n7389;
  assign n7391 = n2907_1 & ~n7390;
  assign n7392 = ~n7375 & ~n7391;
  assign n7393 = ~n7374 & n7392;
  assign n7394 = ~n7373 & n7393;
  assign n3632 = n7372 | ~n7394;
  assign n7396 = ppeakp_12_12_ & ~n3035;
  assign n7397 = \[14120]  & n2936;
  assign n7398 = \[4940]  & n2964;
  assign n7399 = \[11510]  & n3044;
  assign n7400 = \[7775]  & n2961;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = \[4415]  & n3020;
  assign n7403 = \[7190]  & n3030;
  assign n7404 = ~n7402 & ~n7403;
  assign n7405 = n7401 & n7404;
  assign n7406 = ~n7398 & n7405;
  assign n7407 = n2907_1 & ~n7406;
  assign n7408 = ~n7397 & ~n7407;
  assign n7409 = ppeakb_12_12_ & ppeaka_12_12_;
  assign n7410 = n2912_1 & ~n7409;
  assign n7411 = n7408 & ~n7410;
  assign n7412 = ~n4977 & n7411;
  assign n7413 = ~n7396 & n7412;
  assign n7414 = ~n2906 & ~n7413;
  assign n7415 = ppeaka_13_13_ & n2975_1;
  assign n7416 = \[15845]  & n4453_1;
  assign n7417 = ~n7415 & ~n7416;
  assign n7418 = ~n7414 & n7417;
  assign n7419 = ppeaka_12_12_ & ~n3042_1;
  assign n7420 = ppeakb_12_12_ & n4451;
  assign n7421 = ~n7419 & ~n7420;
  assign n3636 = ~n7418 | ~n7421;
  assign n7423 = ppeakp_3_3_ & ~n3035;
  assign n7424 = ppeaka_3_3_ & ~n3042_1;
  assign n7425 = ppeaka_4_4_ & n2975_1;
  assign n7426 = \[13355]  & n2936;
  assign n7427 = ppeakb_3_3_ & ppeaka_3_3_;
  assign n7428 = n2912_1 & ~n7427;
  assign n7429 = ~n7426 & ~n7428;
  assign n7430 = ~n7425 & n7429;
  assign n7431 = \[15560]  & n3021;
  assign n7432 = \[13625]  & n2961;
  assign n7433 = \[9920]  & n3044;
  assign n7434 = ~n7432 & ~n7433;
  assign n7435 = ppeakb_3_3_ & ~n3050;
  assign n7436 = \[15245]  & n3030;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = \[15860]  & ~n3047;
  assign n7439 = \[8960]  & n2964;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = n7437 & n7440;
  assign n7442 = n7434 & n7441;
  assign n7443 = n2907_1 & ~n7442;
  assign n7444 = ~n7431 & ~n7443;
  assign n7445 = ~n5374 & n7444;
  assign n7446 = n7430 & n7445;
  assign n7447 = ~n7424 & n7446;
  assign n3640 = n7423 | ~n7447;
  assign n7449 = \[15140]  & ~n3065;
  assign n7450 = \[10730]  & n3068;
  assign n7451 = ~n7449 & ~n7450;
  assign n7452 = \[10070]  & n2931;
  assign n7453 = \[5975]  & n2917;
  assign n7454 = ~n7452 & ~n7453;
  assign n3644 = ~n7451 | ~n7454;
  assign n7456 = ppeaks_8_8_ & ~n3090;
  assign n7457 = \[15365]  & n3081_1;
  assign n7458 = \[9440]  & n2917;
  assign n7459 = \[7595]  & n3021;
  assign n7460 = ~n7458 & ~n7459;
  assign n7461 = \[10775]  & n3095;
  assign n7462 = \[7340]  & n2912_1;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = \[13385]  & n2936;
  assign n7465 = \[8915]  & n3068;
  assign n7466 = \[13160]  & n2949;
  assign n7467 = \[7520]  & n2964;
  assign n7468 = \[12590]  & n2939;
  assign n7469 = ~n7467 & ~n7468;
  assign n7470 = \[6815]  & n2959;
  assign n7471 = \[10865]  & n2955_1;
  assign n7472 = \[6095]  & n2961;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = ~n7470 & n7473;
  assign n7475 = n7469 & n7474;
  assign n7476 = ~n7466 & n7475;
  assign n7477 = n2907_1 & ~n7476;
  assign n7478 = ~n7465 & ~n7477;
  assign n7479 = ~n7464 & n7478;
  assign n7480 = n7463 & n7479;
  assign n7481 = \[13460]  & n2931;
  assign n7482 = n7480 & ~n7481;
  assign n7483 = n7460 & n7482;
  assign n7484 = ~n4445 & n7483;
  assign n7485 = ~n2906 & ~n7484;
  assign n7486 = ~n7457 & ~n7485;
  assign n3649 = n7456 | ~n7486;
  assign n7488 = ppeakp_15_15_ & ~n3147;
  assign n7489 = ppeaka_15_15_ & ~n3156;
  assign n7490 = \[11450]  & n3021;
  assign n7491 = ~n7489 & ~n7490;
  assign n7492 = ~n7488 & n7491;
  assign n7493 = \[11285]  & n3095;
  assign n7494 = ppeakb_15_15_ & n2917;
  assign n7495 = \[8210]  & ~n2927;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7493 & n7496;
  assign n3653 = ~n7492 | ~n7497;
  assign n7499 = ~pdata_9_9_ & n3175;
  assign n7500 = ~\[15185]  & ~n3175;
  assign n7501 = ~preset & ~n7500;
  assign n3657 = ~n7499 & n7501;
  assign n7503 = ~\[15200]  & ~n3181;
  assign n7504 = ~pdata_6_6_ & n3181;
  assign n7505 = ~preset & ~n7504;
  assign n3662 = ~n7503 & n7505;
  assign n7507 = ~\[15215]  & ~n3181;
  assign n7508 = ~pdata_15_15_ & n3181;
  assign n7509 = ~preset & ~n7508;
  assign n3667 = ~n7507 & n7509;
  assign n7511 = \[15230]  & n3194_1;
  assign n3672 = n4846 | n7511;
  assign n7513 = ~\[15245]  & ~n3203;
  assign n7514 = ~pdata_3_3_ & n3203;
  assign n7515 = ~preset & ~n7514;
  assign n3677 = ~n7513 & n7515;
  assign n7517 = ~\[15260]  & ~n3218;
  assign n7518 = ~pdata_12_12_ & n3218;
  assign n7519 = ~preset & ~n7518;
  assign n3682 = ~n7517 & n7519;
  assign n7521 = \[15275]  & n3225;
  assign n7522 = pdata_9_9_ & n3963;
  assign n3687 = n7521 | n7522;
  assign n7524 = ~\[15290]  & ~n3231;
  assign n7525 = ~pdata_2_2_ & n3231;
  assign n7526 = ~preset & ~n7525;
  assign n3692 = ~n7524 & n7526;
  assign n7528 = \[15305]  & n3240;
  assign n3697 = n5464 | n7528;
  assign n7530 = n4161 & ~n3646;
  assign n7531 = \[15320]  & n3312;
  assign n3702 = n7530 | n7531;
  assign n7533 = ~n3549 & n4428;
  assign n7534 = \[15335]  & n3178;
  assign n3707 = n7533 | n7534;
  assign n7536 = ~\[15350]  & ~n3265;
  assign n7537 = n3265 & ~n4605;
  assign n7538 = ~preset & ~n7537;
  assign n3712 = ~n7536 & n7538;
  assign n7540 = n3963 & ~n4626;
  assign n7541 = \[15365]  & n3225;
  assign n3717 = n7540 | n7541;
  assign n7543 = ~\[15380]  & ~n3231;
  assign n7544 = n3231 & n4298;
  assign n7545 = ~preset & ~n7544;
  assign n3722 = ~n7543 & n7545;
  assign n7547 = ~\[15395]  & ~n3717_1;
  assign n7548 = n3717_1 & ~n4399;
  assign n7549 = ~preset & ~n7548;
  assign n3727 = ~n7547 & n7549;
  assign n7551 = ~\[15410]  & ~n3717_1;
  assign n7552 = n3717_1 & n4692;
  assign n7553 = ~preset & ~n7552;
  assign n3732 = ~n7551 & n7553;
  assign n7555 = ~n4955 & n6333;
  assign n7556 = \[15425]  & n6335;
  assign n3737 = n7555 | n7556;
  assign n7558 = ~\[15440]  & ~n2843;
  assign n7559 = ~pdata_4_4_ & n2843;
  assign n7560 = ~preset & ~n7559;
  assign n3742 = ~n7558 & n7560;
  assign n7562 = ppeakb_6_6_ & ~n2989;
  assign n7563 = \[7685]  & n2931;
  assign n7564 = \[4385]  & n2936;
  assign n7565 = \[7745]  & n2912_1;
  assign n7566 = ppeaka_6_6_ & ~n2950_1;
  assign n7567 = \[7865]  & n2959;
  assign n7568 = \[7160]  & n2961;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = \[6575]  & n2955_1;
  assign n7571 = \[10265]  & n2916_1;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = \[13685]  & n2939;
  assign n7574 = n7572 & ~n7573;
  assign n7575 = \[4610]  & n2964;
  assign n7576 = \[15635]  & n2952;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = n7574 & n7577;
  assign n7579 = n7569 & n7578;
  assign n7580 = ~n7566 & n7579;
  assign n7581 = n2907_1 & ~n7580;
  assign n7582 = ~n7565 & ~n7581;
  assign n7583 = ~n7564 & n7582;
  assign n7584 = ~n7563 & n7583;
  assign n3747 = n7562 | ~n7584;
  assign n7586 = ppeakp_15_15_ & ~n3035;
  assign n7587 = ppeaka_15_15_ & ~n3042_1;
  assign n7588 = ppeakb_15_15_ & ppeaka_15_15_;
  assign n7589 = n2912_1 & ~n7588;
  assign n7590 = \[13730]  & n2936;
  assign n7591 = ppeakb_15_15_ & n4451;
  assign n7592 = \[15215]  & n3020;
  assign n7593 = \[13550]  & ~n3047;
  assign n7594 = \[7205]  & n3030;
  assign n7595 = \[6365]  & n3044;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7593 & n7596;
  assign n7598 = \[15950]  & n2961;
  assign n7599 = \[7010]  & n2964;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = n7597 & n7600;
  assign n7602 = ~n7592 & n7601;
  assign n7603 = n2907_1 & ~n7602;
  assign n7604 = ~n4760 & ~n7603;
  assign n7605 = ~n7591 & n7604;
  assign n7606 = ~n7590 & n7605;
  assign n7607 = ~n7589 & n7606;
  assign n7608 = ~n7587 & n7607;
  assign n3751 = n7586 | ~n7608;
  assign n7610 = ppeakp_4_4_ & ~n3035;
  assign n7611 = ppeaka_4_4_ & ~n3042_1;
  assign n7612 = ppeaka_5_5_ & n2975_1;
  assign n7613 = \[14525]  & n2936;
  assign n7614 = ppeakb_4_4_ & ppeaka_4_4_;
  assign n7615 = n2912_1 & ~n7614;
  assign n7616 = ~n7613 & ~n7615;
  assign n7617 = ~n7612 & n7616;
  assign n7618 = ppeakb_4_4_ & n4451;
  assign n7619 = \[15905]  & n3020;
  assign n7620 = \[14765]  & ~n3047;
  assign n7621 = \[14870]  & n3030;
  assign n7622 = \[8300]  & n2964;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = ~n7620 & n7623;
  assign n7625 = \[8975]  & n3044;
  assign n7626 = \[13280]  & n2961;
  assign n7627 = ~n7625 & ~n7626;
  assign n7628 = n7624 & n7627;
  assign n7629 = ~n7619 & n7628;
  assign n7630 = n2907_1 & ~n7629;
  assign n7631 = ~n4197 & ~n7630;
  assign n7632 = ~n7618 & n7631;
  assign n7633 = n7617 & n7632;
  assign n7634 = ~n7611 & n7633;
  assign n3755 = n7610 | ~n7634;
  assign n7636 = \[15500]  & ~n3065;
  assign n7637 = \[15305]  & n2917;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = \[9800]  & n2931;
  assign n7640 = \[10445]  & n3068;
  assign n7641 = ~n7639 & ~n7640;
  assign n3759 = ~n7638 | ~n7641;
  assign n7643 = \[15515]  & ~n3065;
  assign n7644 = \[8930]  & n3068;
  assign n7645 = ~n7643 & ~n7644;
  assign n7646 = \[13475]  & n2931;
  assign n7647 = \[9710]  & n2917;
  assign n7648 = ~n7646 & ~n7647;
  assign n3764 = ~n7645 | ~n7648;
  assign n7650 = \[10670]  & n3020;
  assign n7651 = \[6125]  & n2959;
  assign n7652 = \[12890]  & n2949;
  assign n7653 = \[5390]  & n2961;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~n7651 & n7654;
  assign n7656 = \[9455]  & n2964;
  assign n7657 = \[7415]  & n2955_1;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = n7655 & n7658;
  assign n7660 = ~n7650 & n7659;
  assign n7661 = n2907_1 & ~n7660;
  assign n7662 = \[15380]  & n2940_1;
  assign n7663 = \[9935]  & n3095;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = ~n7661 & n7664;
  assign n7666 = \[5330]  & n2912_1;
  assign n7667 = \[13175]  & n3068;
  assign n7668 = \[7490]  & n2917;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = \[13025]  & n2936;
  assign n7671 = n7669 & ~n7670;
  assign n7672 = ~n7666 & n7671;
  assign n7673 = \[12605]  & n2931;
  assign n7674 = n7672 & ~n7673;
  assign n7675 = n7665 & n7674;
  assign n7676 = ~n6918 & n7675;
  assign n7677 = ~n2906 & ~n7676;
  assign n7678 = ppeaks_0_0_ & ~n3090;
  assign n7679 = \[13400]  & n3081_1;
  assign n7680 = ~n7678 & ~n7679;
  assign n3769 = n7677 | ~n7680;
  assign n7682 = ~pdata_12_12_ & n3175;
  assign n7683 = ~\[15545]  & ~n3175;
  assign n7684 = ~preset & ~n7683;
  assign n3773 = ~n7682 & n7684;
  assign n7686 = ~\[15560]  & ~n3181;
  assign n7687 = ~pdata_3_3_ & n3181;
  assign n7688 = ~preset & ~n7687;
  assign n3778 = ~n7686 & n7688;
  assign n7690 = ~\[15575]  & ~n3181;
  assign n7691 = ~pdata_14_14_ & n3181;
  assign n7692 = ~preset & ~n7691;
  assign n3783 = ~n7690 & n7692;
  assign n7694 = \[15590]  & n3194_1;
  assign n3788 = n5249 | n7694;
  assign n7696 = \[15605]  & n3194_1;
  assign n3793 = n7317 | n7696;
  assign n7698 = ~\[15620]  & ~n3218;
  assign n7699 = ~pdata_15_15_ & n3218;
  assign n7700 = ~preset & ~n7699;
  assign n3798 = ~n7698 & n7700;
  assign n7702 = \[15635]  & n3225;
  assign n7703 = n3177 & n3224_1;
  assign n3803 = n7702 | n7703;
  assign n7705 = ~\[15650]  & ~n3231;
  assign n7706 = ~pdata_1_1_ & n3231;
  assign n7707 = ~preset & ~n7706;
  assign n3808 = ~n7705 & n7707;
  assign n7709 = \[15665]  & n3240;
  assign n3813 = n5679 | n7709;
  assign n7711 = ~n3310 & n4428;
  assign n7712 = \[15680]  & n3178;
  assign n3818 = n7711 | n7712;
  assign n7714 = ~n4626 & n4428;
  assign n7715 = \[15695]  & n3178;
  assign n3823 = n7714 | n7715;
  assign n7717 = ~\[15710]  & ~n3265;
  assign n7718 = n3265 & ~n3660;
  assign n7719 = ~preset & ~n7718;
  assign n3828 = ~n7717 & n7719;
  assign n7721 = ~\[15725]  & ~n3218;
  assign n7722 = n3218 & n3646;
  assign n7723 = ~preset & ~n7722;
  assign n3833 = ~n7721 & n7723;
  assign n7725 = ~\[15755]  & ~n3691;
  assign n7726 = n3691 & ~n4111;
  assign n7727 = ~preset & ~n7726;
  assign n3838 = ~n7725 & n7727;
  assign n7729 = n4087_1 & n4091;
  assign n7730 = \[15770]  & n4097_1;
  assign n3843 = n7729 | n7730;
  assign n7732 = ~\[15785]  & ~n2843;
  assign n7733 = ~pdata_3_3_ & n2843;
  assign n7734 = ~preset & ~n7733;
  assign n3848 = ~n7732 & n7734;
  assign n7736 = ppeakb_7_7_ & ~n2989;
  assign n7737 = \[15980]  & n3081_1;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = \[6500]  & n2936;
  assign n7740 = \[7055]  & n2931;
  assign n7741 = \[7115]  & n2912_1;
  assign n7742 = \[5915]  & n2959;
  assign n7743 = \[9095]  & n2961;
  assign n7744 = \[13340]  & n2939;
  assign n7745 = \[14450]  & n2955_1;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = ~n7743 & n7746;
  assign n7748 = \[5315]  & n2964;
  assign n7749 = \[14930]  & n2916_1;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = n7747 & n7750;
  assign n7752 = ~n7742 & n7751;
  assign n7753 = n2907_1 & ~n7752;
  assign n7754 = ~n7741 & ~n7753;
  assign n7755 = ~n7740 & n7754;
  assign n7756 = ~n7739 & n7755;
  assign n7757 = ~n2906 & ~n7756;
  assign n7758 = ppeaka_7_7_ & n4124;
  assign n7759 = ~n7757 & ~n7758;
  assign n3853 = ~n7738 | ~n7759;
  assign n7761 = ppeakb_14_14_ & ppeaka_14_14_;
  assign n7762 = n2912_1 & ~n7761;
  assign n7763 = \[15575]  & n3021;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = ppeakp_14_14_ & ~n3035;
  assign n7766 = \[9080]  & n2961;
  assign n7767 = \[14435]  & n3030;
  assign n7768 = \[6335]  & n2964;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = \[8315]  & n3044;
  assign n7771 = n7769 & ~n7770;
  assign n7772 = ~n7766 & n7771;
  assign n7773 = n2907_1 & ~n7772;
  assign n7774 = \[13370]  & n2936;
  assign n7775 = ~n4493 & ~n7774;
  assign n7776 = ~n7773 & n7775;
  assign n7777 = ~n7765 & n7776;
  assign n7778 = n7764 & n7777;
  assign n7779 = ~n2906 & ~n7778;
  assign n7780 = ppeaka_15_15_ & n2975_1;
  assign n7781 = \[15140]  & n4453_1;
  assign n7782 = ~n7780 & ~n7781;
  assign n7783 = ~n7779 & n7782;
  assign n7784 = ppeaka_14_14_ & ~n3042_1;
  assign n7785 = ppeakb_14_14_ & n4451;
  assign n7786 = ~n7784 & ~n7785;
  assign n3857 = ~n7783 | ~n7786;
  assign n7788 = ppeakp_5_5_ & ~n3035;
  assign n7789 = ppeaka_5_5_ & ~n3042_1;
  assign n7790 = ppeakb_5_5_ & ppeaka_5_5_;
  assign n7791 = n2912_1 & ~n7790;
  assign n7792 = \[14105]  & n2936;
  assign n7793 = ppeaka_6_6_ & n2975_1;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = ~n7791 & n7794;
  assign n7796 = \[14825]  & n3021;
  assign n7797 = \[8330]  & ~n3047;
  assign n7798 = \[6560]  & n3030;
  assign n7799 = \[7670]  & n2964;
  assign n7800 = \[15590]  & n2961;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7798 & n7801;
  assign n7803 = ppeakb_5_5_ & ~n3050;
  assign n7804 = \[5660]  & n3044;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = n7802 & n7805;
  assign n7807 = ~n7797 & n7806;
  assign n7808 = n2907_1 & ~n7807;
  assign n7809 = ~n3093 & ~n7808;
  assign n7810 = ~n7796 & n7809;
  assign n7811 = n7795 & n7810;
  assign n7812 = ~n7789 & n7811;
  assign n3861 = n7788 | ~n7812;
  assign n7814 = \[15845]  & ~n3065;
  assign n7815 = \[8285]  & n3068;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = \[9500]  & n2931;
  assign n7818 = \[9980]  & n2917;
  assign n7819 = ~n7817 & ~n7818;
  assign n3865 = ~n7816 | ~n7819;
  assign n7821 = \[15860]  & ~n3065;
  assign n7822 = \[15665]  & n2917;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = \[13130]  & n2931;
  assign n7825 = \[10145]  & n3068;
  assign n7826 = ~n7824 & ~n7825;
  assign n3870 = ~n7823 | ~n7826;
  assign n7828 = ppeaks_10_10_ & ~n3090;
  assign n7829 = \[14585]  & n3081_1;
  assign n7830 = \[9860]  & n3068;
  assign n7831 = \[10205]  & n3095;
  assign n7832 = \[10400]  & n3021;
  assign n7833 = ~n7042 & ~n7832;
  assign n7834 = ~n7831 & n7833;
  assign n7835 = ~n7830 & n7834;
  assign n7836 = \[6155]  & n2940_1;
  assign n7837 = \[12800]  & n2936;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = \[6035]  & n2912_1;
  assign n7840 = n7838 & ~n7839;
  assign n7841 = \[12860]  & n2931;
  assign n7842 = \[4700]  & n2961;
  assign n7843 = \[8810]  & n2964;
  assign n7844 = \[12665]  & n2949;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = \[5450]  & n2959;
  assign n7847 = \[8135]  & n2916_1;
  assign n7848 = \[8060]  & n2955_1;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7846 & n7849;
  assign n7851 = n7845 & n7850;
  assign n7852 = ~n7842 & n7851;
  assign n7853 = n2907_1 & ~n7852;
  assign n7854 = ~n7841 & ~n7853;
  assign n7855 = n7840 & n7854;
  assign n7856 = n7835 & n7855;
  assign n7857 = ~n2906 & ~n7856;
  assign n7858 = ~n7829 & ~n7857;
  assign n3875 = n7828 | ~n7858;
  assign n7860 = ~pdata_11_11_ & n3175;
  assign n7861 = ~\[15890]  & ~n3175;
  assign n7862 = ~preset & ~n7861;
  assign n3879 = ~n7860 & n7862;
  assign n7864 = ~\[15905]  & ~n3181;
  assign n7865 = ~pdata_4_4_ & n3181;
  assign n7866 = ~preset & ~n7865;
  assign n3884 = ~n7864 & n7866;
  assign n7868 = ~\[15920]  & ~n3181;
  assign n7869 = ~pdata_13_13_ & n3181;
  assign n7870 = ~preset & ~n7869;
  assign n3889 = ~n7868 & n7870;
  assign n7872 = \[15935]  & n3194_1;
  assign n3894 = n5061 | n7872;
  assign n7874 = \[15950]  & n3194_1;
  assign n3899 = n5438 | n7874;
  assign n7876 = ~\[15965]  & ~n3218;
  assign n7877 = ~pdata_14_14_ & n3218;
  assign n7878 = ~preset & ~n7877;
  assign n3904 = ~n7876 & n7878;
  assign n7880 = pdata_7_7_ & n3963;
  assign n7881 = \[15980]  & n3225;
  assign n3909 = n7880 | n7881;
  assign n7883 = ~\[15995]  & ~n3231;
  assign n7884 = ~pdata_0_0_ & n3231;
  assign n7885 = ~preset & ~n7884;
  assign n3914 = ~n7883 & n7885;
  assign n7887 = ~\[16010]  & ~n3231;
  assign n7888 = ~pdata_9_9_ & n3231;
  assign n7889 = ~preset & ~n7888;
  assign n3919 = ~n7887 & n7889;
  assign n7891 = \[16025]  & n3178;
  assign n7892 = ~n4298 & n4428;
  assign n3924 = n7891 | n7892;
  assign n7894 = n3653_1 & n4428;
  assign n7895 = \[16040]  & n3178;
  assign n3929 = n7894 | n7895;
  assign n7897 = ~\[16055]  & ~n3265;
  assign n7898 = n3265 & n3310;
  assign n7899 = ~preset & ~n7898;
  assign n3934 = ~n7897 & n7899;
  assign n7901 = ~\[16070]  & ~n3218;
  assign n7902 = n3218 & n4326;
  assign n7903 = ~preset & ~n7902;
  assign n3939 = ~n7901 & n7903;
  assign n7905 = n3963 & ~n4344_1;
  assign n7906 = \[16085]  & n3225;
  assign n3944 = n7905 | n7906;
  assign n7908 = ~\[16100]  & ~n3691;
  assign n7909 = n3691 & n4365;
  assign n7910 = ~preset & ~n7909;
  assign n3949 = ~n7908 & n7910;
  assign n7912 = ~pdn & n2923;
  assign n7913 = ~\[17791]  & n7912;
  assign n7914 = ~\[18467]  & ~n3688;
  assign n7915 = ~n3689 & ~n7914;
  assign n7916 = ~\[17570]  & n7915;
  assign n7917 = \[17999]  & ~\[18220] ;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = ~n7913 & n7918;
  assign n7920 = ~\[17167]  & n3030;
  assign n7921 = n2880 & n7920;
  assign n7922 = n7919 & ~n7921;
  assign n7923 = ~n3175 & n7922;
  assign n7924 = ~\[17583]  & \[17648] ;
  assign n7925 = ~n3273 & ~n7924;
  assign n7926 = \[16933]  & ~\[17388] ;
  assign n7927 = \[18363]  & ~\[18415] ;
  assign n7928 = ~n7926 & ~n7927;
  assign n7929 = ~\[17414]  & \[17843] ;
  assign n7930 = \[18311]  & ~\[18389] ;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = n7928 & n7931;
  assign n7933 = \[17037]  & ~\[17102] ;
  assign n7934 = ~n3208 & ~n7933;
  assign n7935 = ~\[17050]  & \[17115] ;
  assign n7936 = \[17206]  & ~\[17271] ;
  assign n7937 = ~n3724 & ~n7936;
  assign n7938 = ~\[17518]  & \[17817] ;
  assign n7939 = ~n3706 & ~n7938;
  assign n7940 = n7937 & n7939;
  assign n7941 = ~n7935 & n7940;
  assign n7942 = n7934 & n7941;
  assign n7943 = n7932 & n7942;
  assign n7944 = n7925 & n7943;
  assign n7945 = n7923 & n7944;
  assign n7946 = n3264_1 & n7945;
  assign n7947 = n3568 & ~n7946;
  assign n7948 = ppeakb_8_8_ & n7947;
  assign n7949 = n7938 & ~n7946;
  assign n7950 = ~preset & n7949;
  assign n7951 = \[11420]  & n7950;
  assign n7952 = ~n7948 & ~n7951;
  assign n4032 = ~preset & n7933;
  assign n7954 = n2986 & n7916;
  assign n7955 = ~n4032 & ~n7954;
  assign n7956 = ~n7946 & ~n7955;
  assign n7957 = ppeakp_8_8_ & n7956;
  assign n7958 = ~preset & n7924;
  assign n7959 = \[13460]  & n7958;
  assign n7960 = ~n7957 & ~n7959;
  assign n4097 = ~preset & n7936;
  assign n7962 = ~n7946 & n4097;
  assign n7963 = \[11225]  & n7962;
  assign n4519 = ~preset & n7927;
  assign n7965 = ~n7946 & n4519;
  assign n7966 = \[8000]  & n7965;
  assign n7967 = ~n7963 & ~n7966;
  assign n7968 = n7960 & n7967;
  assign n7969 = n7952 & n7968;
  assign n7970 = n3706 & ~n7946;
  assign n7971 = \[7595]  & n7970;
  assign n7972 = n7916 & ~n7946;
  assign n7973 = n3908 & n7972;
  assign n7974 = paddress_8_8_ & n7946;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = ~n3391 & n7975;
  assign n7977 = ~n7971 & n7976;
  assign n7978 = ~preset & ~n7977;
  assign n4057 = n3255 & n7920;
  assign n7980 = ~n7946 & n4057;
  assign n7981 = ~n3192 & ~n7980;
  assign n7982 = ppeaka_8_8_ & ~n7981;
  assign n7983 = ~preset & ~\[17050] ;
  assign n4012 = \[17115]  & n7983;
  assign n7985 = ~n7946 & n4012;
  assign n7986 = \[13160]  & n7985;
  assign n4510 = ~preset & n7930;
  assign n7988 = ~n7946 & n4510;
  assign n7989 = \[8750]  & n7988;
  assign n7990 = ~n7986 & ~n7989;
  assign n7991 = ~n7982 & n7990;
  assign n7992 = n4082 & ~n7946;
  assign n7993 = \[8915]  & n7992;
  assign n4548 = n3217 & n3255;
  assign n4142 = ~preset & n7926;
  assign n7996 = ~n4548 & ~n4142;
  assign n7997 = ~n3963 & n7996;
  assign n7998 = ~n4161 & n7997;
  assign n4107 = n3230 & n3255;
  assign n4505 = ~preset & n3208;
  assign n8001 = ~n4107 & ~n4505;
  assign n8002 = ~n4428 & n8001;
  assign n8003 = n7998 & n8002;
  assign n8004 = ~n7946 & ~n8003;
  assign n8005 = ppeaks_8_8_ & n8004;
  assign n8006 = ~n7993 & ~n8005;
  assign n8007 = n7991 & n8006;
  assign n8008 = ~n7978 & n8007;
  assign n3954 = ~n7969 | ~n8008;
  assign n8010 = ppeaka_7_7_ & ~n7925;
  assign n8011 = n3700 & n7939;
  assign n8012 = ppeakb_7_7_ & ~n8011;
  assign n8013 = n7925 & n8011;
  assign n8014 = \[16907]  & n8013;
  assign n8015 = ~n8012 & ~n8014;
  assign n8016 = ~n8010 & n8015;
  assign n3958 = ~preset & ~n8016;
  assign n8018 = ~preset & ~\[17388] ;
  assign n8019 = ~\[16933]  & ~n3274;
  assign n3968 = n8018 & ~n8019;
  assign n8021 = ppeaks_9_9_ & n8004;
  assign n8022 = \[10040]  & n7988;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = ppeaka_9_9_ & ~n7981;
  assign n8025 = ppeakb_9_9_ & n7947;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = \[9590]  & n7992;
  assign n8028 = n8026 & ~n8027;
  assign n8029 = n8023 & n8028;
  assign n8030 = \[10685]  & n7970;
  assign n8031 = paddress_9_9_ & n7946;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = n3896 & n7972;
  assign n8034 = ~n3374 & ~n8033;
  assign n8035 = n8032 & n8034;
  assign n8036 = ~preset & ~n8035;
  assign n8037 = \[13820]  & n7958;
  assign n8038 = \[11645]  & n7950;
  assign n8039 = \[15770]  & n7962;
  assign n8040 = ~n8038 & ~n8039;
  assign n8041 = \[12440]  & n7985;
  assign n8042 = \[7370]  & n7965;
  assign n8043 = ppeakp_9_9_ & n7956;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = ~n8041 & n8044;
  assign n8046 = n8040 & n8045;
  assign n8047 = ~n8037 & n8046;
  assign n8048 = ~n8036 & n8047;
  assign n3973 = ~n8029 | ~n8048;
  assign n8050 = ppeaka_8_8_ & ~n7925;
  assign n8051 = \[16959]  & n8013;
  assign n8052 = ppeakb_8_8_ & ~n8011;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = ~n8050 & n8053;
  assign n3977 = ~preset & ~n8054;
  assign n8056 = ~\[16920]  & \[16972] ;
  assign n3982 = ~preset & n8056;
  assign n8058 = ~preset & ~\[18389] ;
  assign n3987 = \[16985]  & n8058;
  assign n8060 = \[16998]  & n8013;
  assign n8061 = ppeaka_5_5_ & ~n7925;
  assign n8062 = ppeakb_5_5_ & ~n8011;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n8060 & n8063;
  assign n3992 = ~preset & ~n8064;
  assign n8066 = ~\[17011]  & n8013;
  assign n3997 = ~preset & ~n8066;
  assign n4002 = ~preset & ~pdn;
  assign n8069 = ~preset & ~\[17102] ;
  assign n8070 = ~\[17037]  & ~\[18025] ;
  assign n4007 = n8069 & ~n8070;
  assign n8072 = ppeakb_6_6_ & ~n8011;
  assign n8073 = ppeaka_6_6_ & ~n7925;
  assign n8074 = \[17063]  & n8013;
  assign n8075 = ~n8073 & ~n8074;
  assign n8076 = ~n8072 & n8075;
  assign n4017 = ~preset & ~n8076;
  assign n8078 = \[17076]  & n8013;
  assign n8079 = ppeakb_15_15_ & ~n8011;
  assign n8080 = ppeaka_15_15_ & ~n7925;
  assign n8081 = ~n8079 & ~n8080;
  assign n8082 = ~n8078 & n8081;
  assign n4022 = ~preset & ~n8082;
  assign n4027 = \[17089]  & n4002;
  assign n8085 = n3697_1 & n7983;
  assign n4037 = n4012 | n8085;
  assign n8087 = \[17128]  & n8013;
  assign n8088 = ppeakb_3_3_ & ~n8011;
  assign n8089 = ppeaka_3_3_ & ~n7925;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = ~n8087 & n8090;
  assign n4042 = ~preset & ~n8091;
  assign n8093 = ~\[17141]  & n8013;
  assign n4047 = ~preset & ~n8093;
  assign n4052 = \[17154]  & n8069;
  assign n8096 = ~preset & ~\[17232] ;
  assign n8097 = ~\[17180]  & ~n3695;
  assign n4062 = n8096 & ~n8097;
  assign n8099 = \[17193]  & n8013;
  assign n8100 = ppeakb_4_4_ & ~n8011;
  assign n8101 = ppeaka_4_4_ & ~n7925;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n8099 & n8102;
  assign n4067 = ~preset & ~n8103;
  assign n8105 = ~preset & ~\[17271] ;
  assign n8106 = ~\[17206]  & ~n3693;
  assign n4072 = n8105 & ~n8106;
  assign n4077 = \[17219]  & n7983;
  assign n8109 = \[17245]  & ~n3711;
  assign n4087 = ~preset & n8109;
  assign n8111 = ppeakb_1_1_ & ~n8011;
  assign n8112 = ppeaka_1_1_ & ~n7925;
  assign n8113 = \[17258]  & n8013;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = ~n8111 & n8114;
  assign n4092 = ~preset & ~n8115;
  assign n8117 = ~\[18376]  & n2955_1;
  assign n8118 = n3255 & n8117;
  assign n4102 = n4505 | n8118;
  assign n4112 = \[17310]  & n8018;
  assign n8121 = ppeakb_2_2_ & ~n8011;
  assign n8122 = ppeaka_2_2_ & ~n7925;
  assign n8123 = \[17323]  & n8013;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~n8121 & n8124;
  assign n4117 = ~preset & ~n8125;
  assign n8127 = ~\[17336]  & n8013;
  assign n4122 = ~preset & ~n8127;
  assign n4127 = \[17349]  & n8105;
  assign n8130 = ~\[17167]  & \[17362] ;
  assign n4132 = ~preset & n8130;
  assign n8132 = ~\[17297]  & \[17375] ;
  assign n4137 = ~preset & n8132;
  assign n8134 = \[16100]  & n7950;
  assign n8135 = \[8645]  & n7965;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = ppeakp_11_11_ & n7956;
  assign n8138 = ppeaks_11_11_ & n8004;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ppeakb_11_11_ & n7947;
  assign n8141 = \[10130]  & n7992;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = n8139 & n8142;
  assign n8144 = n8136 & n8143;
  assign n8145 = \[10115]  & n7970;
  assign n8146 = n4044 & n7972;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = \[13115]  & n7924;
  assign n8149 = paddress_11_11_ & n7946;
  assign n8150 = ~n8148 & ~n8149;
  assign n8151 = n8147 & n8150;
  assign n8152 = ~n3355 & n8151;
  assign n8153 = ~preset & ~n8152;
  assign n8154 = ppeaka_11_11_ & ~n7981;
  assign n8155 = \[10595]  & n7988;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = \[13490]  & n7962;
  assign n8158 = \[12125]  & n7985;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = n8156 & n8159;
  assign n8161 = ~n8153 & n8160;
  assign n4147 = ~n8144 | ~n8161;
  assign n8163 = ~preset & ~\[17414] ;
  assign n4151 = \[17843]  & n8163;
  assign n8165 = ~preset & ~\[17700] ;
  assign n8166 = ~\[17427]  & ~\[17518] ;
  assign n4156 = n8165 & ~n8166;
  assign n8168 = \[10925]  & n7950;
  assign n8169 = ppeakp_10_10_ & n7956;
  assign n8170 = \[13850]  & n7962;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = ~n8168 & n8171;
  assign n8173 = \[9305]  & n7965;
  assign n8174 = \[9860]  & n7992;
  assign n8175 = ppeakb_10_10_ & n7947;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8173 & n8176;
  assign n8178 = n8172 & n8177;
  assign n8179 = n3873 & n7972;
  assign n8180 = \[10400]  & n7970;
  assign n8181 = paddress_10_10_ & n7946;
  assign n8182 = \[12860]  & n7924;
  assign n8183 = ~n3525_1 & ~n8182;
  assign n8184 = ~n8181 & n8183;
  assign n8185 = ~n8180 & n8184;
  assign n8186 = ~n8179 & n8185;
  assign n8187 = ~preset & ~n8186;
  assign n8188 = ppeaks_10_10_ & n8004;
  assign n8189 = \[12665]  & n7985;
  assign n8190 = \[9770]  & n7988;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = ~n8188 & n8191;
  assign n8193 = ppeaka_10_10_ & ~n7981;
  assign n8194 = n8192 & ~n8193;
  assign n8195 = ~n8187 & n8194;
  assign n4166 = ~n8178 | ~n8195;
  assign n8197 = ~\[17479]  & n8013;
  assign n4170 = ~preset & ~n8197;
  assign n8199 = ppeaka_13_13_ & ~n7925;
  assign n8200 = \[17492]  & n8013;
  assign n8201 = ppeakb_13_13_ & ~n8011;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = ~n8199 & n8202;
  assign n4175 = ~preset & ~n8203;
  assign n4180 = \[17505]  & n8163;
  assign n8206 = ~\[17518]  & ~\[17817] ;
  assign n4185 = n8165 & ~n8206;
  assign n8208 = ~preset & ~n2882_1;
  assign n8209 = \[17531]  & n8208;
  assign n4190 = n3255 | n8209;
  assign n8211 = ~\[17752]  & n3174_1;
  assign n8212 = ~preset & \[17544] ;
  assign n8213 = ~n8211 & n8212;
  assign n8214 = n6364 & n8211;
  assign n4195 = n8213 | n8214;
  assign n8216 = \[4775]  & n7988;
  assign n8217 = \[9740]  & n7965;
  assign n8218 = ~n8216 & ~n8217;
  assign n8219 = \[14240]  & n7962;
  assign n8220 = n8218 & ~n8219;
  assign n8221 = ppeakb_13_13_ & n7947;
  assign n8222 = ppeaks_13_13_ & n8004;
  assign n8223 = ppeakp_13_13_ & n7956;
  assign n8224 = ~n8222 & ~n8223;
  assign n8225 = ~n8221 & n8224;
  assign n8226 = n8220 & n8225;
  assign n8227 = \[8885]  & n7970;
  assign n8228 = n4010 & n7972;
  assign n8229 = paddress_13_13_ & n7946;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = ~n3630 & n8230;
  assign n8232 = ~n8227 & n8231;
  assign n8233 = ~preset & ~n8232;
  assign n8234 = ppeaka_13_13_ & ~n7981;
  assign n8235 = \[14690]  & n7985;
  assign n8236 = \[12620]  & n7958;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = ~n8234 & n8237;
  assign n8239 = \[13805]  & n7950;
  assign n8240 = \[10700]  & n7992;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = n8238 & n8241;
  assign n8243 = ~n8233 & n8242;
  assign n4200 = ~n8226 | ~n8243;
  assign n8245 = ~\[17570]  & ~n7915;
  assign n8246 = n2882_1 & n5965;
  assign n8247 = n5905 & n6361;
  assign n8248 = n6431 & n8247;
  assign n8249 = n8246 & n8248;
  assign n8250 = n6534 & n6588;
  assign n8251 = n5789 & n6482;
  assign n8252 = ~n6527 & ~n6579;
  assign n8253 = ~n6258 & ~n6304;
  assign n8254 = n8252 & n8253;
  assign n8255 = n8251 & n8254;
  assign n8256 = n8250 & n8255;
  assign n8257 = n8249 & n8256;
  assign n8258 = \[17596]  & n8257;
  assign n8259 = ~\[18597]  & ~n8258;
  assign n8260 = n2901 & n8259;
  assign n8261 = \[17986]  & ~n8260;
  assign n8262 = ~\[17804]  & ~n8261;
  assign n8263 = ~preset & n8262;
  assign n4204 = ~n8245 & n8263;
  assign n8265 = ~\[17583]  & ~\[17648] ;
  assign n4209 = n8165 & ~n8265;
  assign n8267 = n2876 & ~n8257;
  assign n8268 = ~preset & n8267;
  assign n8269 = n2920_1 & n8262;
  assign n4214 = n8268 | n8269;
  assign n8271 = ~preset & \[17609] ;
  assign n8272 = ~n8211 & n8271;
  assign n8273 = n5792 & n8211;
  assign n4219 = n8272 | n8273;
  assign n8275 = \[10010]  & n7965;
  assign n8276 = \[15755]  & n7950;
  assign n8277 = ppeakb_12_12_ & n7947;
  assign n8278 = ppeaks_12_12_ & n8004;
  assign n8279 = ppeakp_12_12_ & n7956;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = ~n8277 & n8280;
  assign n8282 = ~n8276 & n8281;
  assign n8283 = ~n8275 & n8282;
  assign n8284 = \[9845]  & n7970;
  assign n8285 = n4035 & n7972;
  assign n8286 = paddress_12_12_ & n7946;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~n3316_1 & n8287;
  assign n8289 = ~n8284 & n8288;
  assign n8290 = ~preset & ~n8289;
  assign n8291 = \[14660]  & n7962;
  assign n8292 = \[6860]  & n7988;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = \[12395]  & n7958;
  assign n8295 = n8293 & ~n8294;
  assign n8296 = ppeaka_12_12_ & ~n7981;
  assign n8297 = \[15065]  & n7985;
  assign n8298 = ~n8296 & ~n8297;
  assign n8299 = \[10415]  & n7992;
  assign n8300 = n8298 & ~n8299;
  assign n8301 = n8295 & n8300;
  assign n8302 = ~n8290 & n8301;
  assign n4224 = ~n8283 | ~n8302;
  assign n8304 = ~\[17570]  & ~\[17635] ;
  assign n4228 = n8263 & ~n8304;
  assign n8306 = ~\[17427]  & ~\[17648] ;
  assign n4233 = n8165 & ~n8306;
  assign n4238 = ~preset & n8257;
  assign n8309 = ~preset & \[17674] ;
  assign n8310 = ~n8211 & n8309;
  assign n8311 = n5968 & n8211;
  assign n4243 = n8310 | n8311;
  assign n8313 = ppeakb_15_15_ & n7947;
  assign n8314 = \[8765]  & n7988;
  assign n8315 = \[6320]  & n7992;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = ~n8313 & n8316;
  assign n8318 = \[14615]  & n7950;
  assign n8319 = \[12425]  & n7962;
  assign n8320 = ~n8318 & ~n8319;
  assign n8321 = n8317 & n8320;
  assign n8322 = n3975 & n7972;
  assign n8323 = \[4880]  & n7970;
  assign n8324 = paddress_15_15_ & n7946;
  assign n8325 = \[15050]  & n7924;
  assign n8326 = ~n3579 & ~n8325;
  assign n8327 = ~n8324 & n8326;
  assign n8328 = ~n8323 & n8327;
  assign n8329 = ~n8322 & n8328;
  assign n8330 = ~preset & ~n8329;
  assign n8331 = ppeaka_15_15_ & ~n7981;
  assign n8332 = \[13880]  & n7985;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = ppeakp_15_15_ & n7956;
  assign n8335 = \[6755]  & n7965;
  assign n8336 = ppeaks_15_15_ & n8004;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~n8334 & n8337;
  assign n8339 = n8333 & n8338;
  assign n8340 = ~n8330 & n8339;
  assign n4248 = ~n8321 | ~n8340;
  assign n4252 = \[18142]  & n8165;
  assign n8343 = ~\[17713]  & ~n8211;
  assign n8344 = ~ppeaki_4_4_ & n8211;
  assign n8345 = ~preset & ~n8344;
  assign n4257 = ~n8343 & n8345;
  assign n8347 = ppeaka_14_14_ & ~n7981;
  assign n8348 = ~preset & n7970;
  assign n8349 = \[9560]  & n8348;
  assign n8350 = ~n8347 & ~n8349;
  assign n8351 = \[14270]  & n7985;
  assign n8352 = ppeaks_14_14_ & n8004;
  assign n8353 = ~n8351 & ~n8352;
  assign n8354 = ppeakp_14_14_ & n7956;
  assign n8355 = \[12650]  & n7962;
  assign n8356 = ~n8354 & ~n8355;
  assign n8357 = n8353 & n8356;
  assign n8358 = n8350 & n8357;
  assign n8359 = n4001 & n7972;
  assign n8360 = paddress_14_14_ & n7946;
  assign n8361 = \[15410]  & n7924;
  assign n8362 = ~n3611 & ~n8361;
  assign n8363 = ~n8360 & n8362;
  assign n8364 = ~n8359 & n8363;
  assign n8365 = ~preset & ~n8364;
  assign n8366 = \[6080]  & n7965;
  assign n8367 = ppeakb_14_14_ & n7947;
  assign n8368 = \[10985]  & n7992;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = ~n8366 & n8369;
  assign n8371 = \[13445]  & n7950;
  assign n8372 = \[5480]  & n7988;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = n8370 & n8373;
  assign n8375 = ~n8365 & n8374;
  assign n4262 = ~n8358 | ~n8375;
  assign n4266 = \[17739]  & n8165;
  assign n8378 = ~\[17752]  & ~n3174_1;
  assign n4271 = n8208 & ~n8378;
  assign n8380 = ppeakb_9_9_ & ~n8011;
  assign n8381 = \[17765]  & n8013;
  assign n8382 = ppeaka_9_9_ & ~n7925;
  assign n8383 = ~n8381 & ~n8382;
  assign n8384 = ~n8380 & n8383;
  assign n4276 = ~preset & ~n8384;
  assign n8386 = \[17778]  & n8013;
  assign n8387 = ppeakb_14_14_ & ~n8011;
  assign n8388 = ppeaka_14_14_ & ~n7925;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = ~n8386 & n8389;
  assign n4281 = ~preset & ~n8390;
  assign n8392 = ~\[17791]  & ~n7912;
  assign n4286 = n8163 & ~n8392;
  assign n4291 = n4002 & ~n8262;
  assign n8395 = ~\[17817]  & ~n3690;
  assign n4296 = n8165 & ~n8395;
  assign n8397 = \[17050]  & ~\[17219] ;
  assign n8398 = \[17232]  & ~\[18441] ;
  assign n8399 = pwr_0_0_ & ~n8398;
  assign n8400 = ~n8397 & n8399;
  assign n8401 = ~\[17427]  & \[17518] ;
  assign n8402 = \[17271]  & ~\[17349] ;
  assign n8403 = \[17583]  & ~\[18077] ;
  assign n8404 = ~n8402 & ~n8403;
  assign n8405 = ~n8401 & n8404;
  assign n8406 = n8400 & n8405;
  assign n8407 = n7934 & n8406;
  assign n8408 = n7941 & ~n8407;
  assign n8409 = n7925 & n8408;
  assign n4301 = ~preset & ~n8409;
  assign n8411 = ~\[17791]  & ~\[17843] ;
  assign n4305 = n8163 & ~n8411;
  assign n8413 = ~\[17856]  & ~n2903;
  assign n4310 = ~preset & ~n8413;
  assign n8415 = ~\[17869]  & n8013;
  assign n4315 = ~preset & ~n8415;
  assign n8417 = ~\[17882]  & n8013;
  assign n4320 = ~preset & ~n8417;
  assign n8419 = ~\[16985]  & \[18389] ;
  assign n8420 = ~n6026 & ~n8419;
  assign n8421 = \[18415]  & ~\[18480] ;
  assign n8422 = ~n5842 & ~n8421;
  assign n8423 = \[17297]  & ~\[17375] ;
  assign n8424 = \[16920]  & ~\[16972] ;
  assign n8425 = ~n8423 & ~n8424;
  assign n8426 = n8422 & n8425;
  assign n8427 = n8420 & n8426;
  assign n8428 = ~\[18298]  & \[18376] ;
  assign n8429 = ~n3162 & ~n8428;
  assign n8430 = ~\[18428]  & \[18493] ;
  assign n8431 = ~n2843 & ~n8430;
  assign n8432 = n8429 & n8431;
  assign n8433 = ~n3181 & ~n5777;
  assign n8434 = n7934 & n8433;
  assign n8435 = n8432 & n8434;
  assign n8436 = ~n3249_1 & n7932;
  assign n8437 = n8435 & n8436;
  assign n8438 = ~n3203 & n8437;
  assign n8439 = n7923 & n8438;
  assign n8440 = n8427 & n8439;
  assign n8441 = n3270 & n8440;
  assign n8442 = ~n3192 & ~n3238;
  assign n8443 = ~n4032 & ~n4519;
  assign n8444 = ~n4151 & n8443;
  assign n8445 = ~n4510 & n8444;
  assign n8446 = ~n4057 & n8445;
  assign n8447 = n8003 & n8446;
  assign n8448 = n8442 & n8447;
  assign n8449 = ~n8441 & ~n8448;
  assign n8450 = n7919 & ~n8441;
  assign n8451 = ~prd_0_0_ & n8441;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = ~preset & n8452;
  assign n4325 = n8449 | n8453;
  assign n8455 = ~\[17908]  & n8013;
  assign n4329 = ~preset & ~n8455;
  assign n8457 = \[17921]  & n8013;
  assign n8458 = ppeaka_10_10_ & ~n7925;
  assign n8459 = ppeakb_10_10_ & ~n8011;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = ~n8457 & n8460;
  assign n4334 = ~preset & ~n8461;
  assign n8463 = ~\[17934]  & n8013;
  assign n4339 = ~preset & ~n8463;
  assign n8465 = ~\[17947]  & n8013;
  assign n4344 = ~preset & ~n8465;
  assign n8467 = ~\[17960]  & n8013;
  assign n4349 = ~preset & ~n8467;
  assign n8469 = \[17973]  & n8013;
  assign n8470 = ppeakb_12_12_ & ~n8011;
  assign n8471 = ppeaka_12_12_ & ~n7925;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = ~n8469 & n8472;
  assign n4354 = ~preset & ~n8473;
  assign n8475 = ~\[17635]  & ~\[17986] ;
  assign n4359 = n8263 & ~n8475;
  assign n8477 = ~\[17999]  & ~\[18077] ;
  assign n4364 = n8165 & ~n8477;
  assign n8479 = ~\[17531]  & n2880;
  assign n8480 = ~preset & \[18012] ;
  assign n8481 = ~n8479 & n8480;
  assign n8482 = n6434 & n8479;
  assign n4369 = n8481 | n8482;
  assign n8484 = ~\[18025]  & ~n3701;
  assign n4374 = n8069 & ~n8484;
  assign n8486 = ~\[18038]  & n8013;
  assign n4379 = ~preset & ~n8486;
  assign n8488 = ~\[17414]  & n8262;
  assign n4384 = n4002 & ~n8488;
  assign n8490 = ~preset & n3690;
  assign n8491 = \[18064]  & n4002;
  assign n4388 = n8490 | n8491;
  assign n8493 = ~\[17583]  & ~\[18077] ;
  assign n4393 = n8165 & ~n8493;
  assign n8495 = n2852 & n3255;
  assign n8496 = ~preset & \[18090] ;
  assign n8497 = ~n8479 & n8496;
  assign n4398 = n8495 | n8497;
  assign n8499 = \[18103]  & ~\[18168] ;
  assign n4403 = ~preset & n8499;
  assign n8501 = ~\[18116]  & n8013;
  assign n4408 = ~preset & ~n8501;
  assign n8503 = ~preset & \[18129] ;
  assign n4413 = n8490 | n8503;
  assign n8505 = ~\[18142]  & ~\[18220] ;
  assign n4418 = n8165 & ~n8505;
  assign n8507 = n2849_1 & n3255;
  assign n8508 = ~preset & \[18155] ;
  assign n8509 = ~n8479 & n8508;
  assign n4423 = n8507 | n8509;
  assign n8511 = ~\[18181]  & n8013;
  assign n4433 = ~preset & ~n8511;
  assign n8513 = \[18194]  & n8013;
  assign n8514 = ppeaka_11_11_ & ~n7925;
  assign n8515 = ppeakb_11_11_ & ~n8011;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = ~n8513 & n8516;
  assign n4438 = ~preset & ~n8517;
  assign n8519 = ~\[18207]  & ~n2903;
  assign n4443 = n4002 & ~n8519;
  assign n8521 = ~\[17999]  & ~\[18220] ;
  assign n4448 = n8165 & ~n8521;
  assign n8523 = n2859 & n3255;
  assign n8524 = ~preset & \[18233] ;
  assign n8525 = ~n8479 & n8524;
  assign n4453 = n8523 | n8525;
  assign n8527 = ~\[17453]  & \[18246] ;
  assign n4458 = ~preset & n8527;
  assign n8529 = \[10670]  & n7970;
  assign n8530 = n3817 & n7972;
  assign n8531 = \[12605]  & n7924;
  assign n8532 = ~n8530 & ~n8531;
  assign n8533 = paddress_0_0_ & n7946;
  assign n8534 = ~n3280 & ~n8533;
  assign n8535 = n8532 & n8534;
  assign n8536 = ~n8529 & n8535;
  assign n8537 = ~preset & ~n8536;
  assign n8538 = \[12890]  & n4012;
  assign n8539 = \[8240]  & n4097;
  assign n8540 = ~n4151 & ~n8539;
  assign n8541 = ppeakb_0_0_ & n3568;
  assign n8542 = n8540 & ~n8541;
  assign n8543 = ~n8538 & n8542;
  assign n8544 = \[10025]  & n4510;
  assign n8545 = n8543 & ~n8544;
  assign n8546 = \[13175]  & n4082;
  assign n8547 = n8545 & ~n8546;
  assign n8548 = ppeaks_0_0_ & ~n8003;
  assign n8549 = n8547 & ~n8548;
  assign n8550 = ~n7946 & ~n8549;
  assign n8551 = \[8630]  & n7965;
  assign n8552 = ppeaka_0_0_ & ~n7981;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 = ppeakp_0_0_ & n7956;
  assign n8555 = \[11630]  & n7950;
  assign n8556 = ~n8554 & ~n8555;
  assign n8557 = n8553 & n8556;
  assign n8558 = ~n8550 & n8557;
  assign n4463 = n8537 | ~n8558;
  assign n8560 = \[17700]  & ~\[17739] ;
  assign n8561 = ~preset & piack_0_0_;
  assign n8562 = ~n8560 & n8561;
  assign n4467 = n4252 | n8562;
  assign n8564 = ~preset & ~\[18415] ;
  assign n8565 = ~\[18285]  & ~n3190;
  assign n4471 = n8564 & ~n8565;
  assign n8567 = \[18298]  & ~\[18376] ;
  assign n4476 = ~preset & n8567;
  assign n8569 = ~\[18311]  & ~\[18506] ;
  assign n4481 = n8058 & ~n8569;
  assign n8571 = ppeakb_1_1_ & n7947;
  assign n8572 = \[6305]  & n7962;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = \[9830]  & n8348;
  assign n8575 = \[10310]  & n7988;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = n8573 & n8576;
  assign n8578 = ppeaks_1_1_ & n8004;
  assign n8579 = \[9290]  & n7965;
  assign n8580 = ~n8578 & ~n8579;
  assign n8581 = \[12005]  & n7985;
  assign n8582 = n8580 & ~n8581;
  assign n8583 = n8577 & n8582;
  assign n8584 = ppeaka_1_1_ & ~n7981;
  assign n8585 = \[9485]  & n7950;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = ppeakp_1_1_ & n7956;
  assign n8588 = \[12920]  & n7992;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = \[12380]  & n7924;
  assign n8591 = ~n3294 & ~n8590;
  assign n8592 = paddress_1_1_ & n7946;
  assign n8593 = ~n3799 & ~n7917;
  assign n8594 = ~n7918 & ~n8593;
  assign n8595 = ~n7946 & n8594;
  assign n8596 = ~n8592 & ~n8595;
  assign n8597 = n8591 & n8596;
  assign n8598 = ~preset & ~n8597;
  assign n8599 = n8589 & ~n8598;
  assign n8600 = n8586 & n8599;
  assign n4486 = ~n8583 | ~n8600;
  assign n8602 = \[18337]  & n8013;
  assign n8603 = ppeaka_0_0_ & ~n7925;
  assign n8604 = ppeakb_0_0_ & ~n8011;
  assign n8605 = ~n8603 & ~n8604;
  assign n8606 = ~n8602 & n8605;
  assign n4490 = ~preset & ~n8606;
  assign n8608 = ~\[18350]  & n8013;
  assign n4495 = ~preset & ~n8608;
  assign n8610 = ~\[18285]  & ~\[18363] ;
  assign n4500 = n8564 & ~n8610;
  assign n8612 = ppeakp_2_2_ & n7956;
  assign n8613 = \[13100]  & n7958;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = \[4760]  & n7988;
  assign n8616 = \[15425]  & n7985;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = n8614 & n8617;
  assign n8619 = ppeaka_2_2_ & ~n7981;
  assign n8620 = \[9725]  & n7965;
  assign n8621 = \[6980]  & n7962;
  assign n8622 = ~n8620 & ~n8621;
  assign n8623 = ~n8619 & n8622;
  assign n8624 = n8618 & n8623;
  assign n8625 = \[10100]  & n7970;
  assign n8626 = paddress_2_2_ & n7946;
  assign n8627 = ~n8625 & ~n8626;
  assign n8628 = n3785 & n7972;
  assign n8629 = ~n3477_1 & ~n8628;
  assign n8630 = n8627 & n8629;
  assign n8631 = ~preset & ~n8630;
  assign n8632 = \[7535]  & n7950;
  assign n8633 = ppeaks_2_2_ & n8004;
  assign n8634 = \[12680]  & n7992;
  assign n8635 = ~n8633 & ~n8634;
  assign n8636 = ~n8632 & n8635;
  assign n8637 = ppeakb_2_2_ & n7947;
  assign n8638 = n8636 & ~n8637;
  assign n8639 = ~n8631 & n8638;
  assign n4515 = ~n8624 | ~n8639;
  assign n8641 = \[18428]  & ~\[18493] ;
  assign n4524 = ~preset & n8641;
  assign n4529 = \[18441]  & n8096;
  assign n8644 = ppeaka_3_3_ & ~n7981;
  assign n8645 = \[6845]  & n7988;
  assign n8646 = \[12455]  & n7992;
  assign n8647 = ~n8645 & ~n8646;
  assign n8648 = ~n8644 & n8647;
  assign n8649 = \[8165]  & n7950;
  assign n8650 = \[4910]  & n7962;
  assign n8651 = \[14255]  & n7985;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = ~n8649 & n8652;
  assign n8654 = n8648 & n8653;
  assign n8655 = n3765 & n7972;
  assign n8656 = \[5570]  & n7970;
  assign n8657 = paddress_3_3_ & n7946;
  assign n8658 = \[12845]  & n7924;
  assign n8659 = ~n3454 & ~n8658;
  assign n8660 = ~n8657 & n8659;
  assign n8661 = ~n8656 & n8660;
  assign n8662 = ~n8655 & n8661;
  assign n8663 = ~preset & ~n8662;
  assign n8664 = ppeakp_3_3_ & n7956;
  assign n8665 = ppeaks_3_3_ & n8004;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = \[9995]  & n7965;
  assign n8668 = ppeakb_3_3_ & n7947;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = n8666 & n8669;
  assign n8671 = ~n8663 & n8670;
  assign n4534 = ~n8654 | ~n8671;
  assign n8673 = ~\[17700]  & n3689;
  assign n8674 = n4002 & ~n8673;
  assign n4538 = ~n7914 & n8674;
  assign n4543 = \[18480]  & n8564;
  assign n8677 = ~\[18506]  & ~n3236;
  assign n4553 = n8058 & ~n8677;
  assign n8679 = ppeaka_4_4_ & ~n7981;
  assign n8680 = \[5615]  & n7962;
  assign n8681 = ~n8679 & ~n8680;
  assign n8682 = ppeakp_4_4_ & n7956;
  assign n8683 = \[5375]  & n7965;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = \[14675]  & n7985;
  assign n8686 = ppeaks_4_4_ & n8004;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = n8684 & n8687;
  assign n8689 = n8681 & n8688;
  assign n8690 = n3756 & n7972;
  assign n8691 = paddress_4_4_ & n7946;
  assign n8692 = \[15035]  & n7924;
  assign n8693 = ~n3496 & ~n8692;
  assign n8694 = ~n8691 & n8693;
  assign n8695 = ~n8690 & n8694;
  assign n8696 = ~preset & ~n8695;
  assign n8697 = \[4865]  & n8348;
  assign n8698 = \[12245]  & n7992;
  assign n8699 = \[6170]  & n7988;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = ~n8697 & n8700;
  assign n8702 = \[6230]  & n7950;
  assign n8703 = ppeakb_4_4_ & n7947;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8701 & n8704;
  assign n8706 = ~n8696 & n8705;
  assign n4558 = ~n8689 | ~n8706;
  assign n8708 = ppeakb_5_5_ & n7947;
  assign n8709 = \[15395]  & n7958;
  assign n8710 = ~n8708 & ~n8709;
  assign n8711 = ppeakp_5_5_ & n7956;
  assign n8712 = \[4670]  & n7965;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = \[11465]  & n7962;
  assign n8715 = \[13505]  & n7985;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = n8713 & n8716;
  assign n8718 = n8710 & n8717;
  assign n8719 = \[9545]  & n7970;
  assign n8720 = paddress_5_5_ & n7946;
  assign n8721 = n3735 & n7972;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = ~n3437_1 & n8722;
  assign n8724 = ~n8719 & n8723;
  assign n8725 = ~preset & ~n8724;
  assign n8726 = ppeaka_5_5_ & ~n7981;
  assign n8727 = \[6995]  & n7992;
  assign n8728 = ppeaks_5_5_ & n8004;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = ~n8726 & n8729;
  assign n8731 = \[6905]  & n7950;
  assign n8732 = \[8105]  & n7988;
  assign n8733 = ~n8731 & ~n8732;
  assign n8734 = n8730 & n8733;
  assign n8735 = ~n8725 & n8734;
  assign n4562 = ~n8718 | ~n8735;
  assign n8737 = pdn & ~\[18545] ;
  assign n8738 = ~preset & ~n8737;
  assign n4566 = ~n3688 & n8738;
  assign n8740 = ppeakp_6_6_ & n7956;
  assign n8741 = \[6740]  & n7965;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = \[14210]  & n7958;
  assign n8744 = \[11690]  & n7962;
  assign n8745 = ppeakb_6_6_ & n7947;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = ~n8743 & n8746;
  assign n8748 = n8742 & n8747;
  assign n8749 = ppeaka_6_6_ & ~n7981;
  assign n8750 = \[7625]  & n7992;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = \[4835]  & n7950;
  assign n8753 = n8751 & ~n8752;
  assign n8754 = n8748 & n8753;
  assign n8755 = \[8870]  & n7970;
  assign n8756 = paddress_6_6_ & n7946;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = n3715 & n7972;
  assign n8759 = ~n3419 & ~n8758;
  assign n8760 = n8757 & n8759;
  assign n8761 = ~preset & ~n8760;
  assign n8762 = ppeaks_6_6_ & n8004;
  assign n8763 = \[7475]  & n7988;
  assign n8764 = ~n8762 & ~n8763;
  assign n8765 = \[13865]  & n7985;
  assign n8766 = n8764 & ~n8765;
  assign n8767 = ~n8761 & n8766;
  assign n4571 = ~n8754 | ~n8767;
  assign n8769 = ~\[18571]  & n8013;
  assign n4575 = ~preset & ~n8769;
  assign n8771 = ~\[18584]  & n8013;
  assign n4580 = ~preset & ~n8771;
  assign n4585 = n4002 & ~n8259;
  assign n8774 = \[18610]  & n8208;
  assign n8775 = ~\[17453]  & ~\[18168] ;
  assign n8776 = n3174_1 & n8775;
  assign n8777 = n3256 & ~n8776;
  assign n4590 = n8774 | n8777;
  assign n8779 = ppeaks_7_7_ & n8004;
  assign n8780 = \[5540]  & n7950;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = \[12905]  & n7985;
  assign n8783 = \[6065]  & n7965;
  assign n8784 = \[8255]  & n7992;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = ~n8782 & n8785;
  assign n8787 = n8781 & n8786;
  assign n8788 = \[8225]  & n7970;
  assign n8789 = n3922 & n7972;
  assign n8790 = \[14630]  & n7924;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = paddress_7_7_ & n7946;
  assign n8793 = ~n3408 & ~n8792;
  assign n8794 = n8791 & n8793;
  assign n8795 = ~n8788 & n8794;
  assign n8796 = ~preset & ~n8795;
  assign n8797 = ppeakb_7_7_ & n7947;
  assign n8798 = ppeakp_7_7_ & n7956;
  assign n8799 = \[9410]  & n7988;
  assign n8800 = ~n8798 & ~n8799;
  assign n8801 = ~n8797 & n8800;
  assign n8802 = ppeaka_7_7_ & ~n7981;
  assign n8803 = \[10970]  & n7962;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = n8801 & n8804;
  assign n8806 = ~n8796 & n8805;
  assign n4595 = ~n8787 | ~n8806;
  assign n8808 = n2880 & n4590;
  assign n8809 = ~\[17232]  & ~\[17271] ;
  assign n8810 = ~\[17297]  & n8809;
  assign n8811 = ~\[17050]  & ~\[17102] ;
  assign n8812 = ~\[16920]  & n8811;
  assign n8813 = n8810 & n8812;
  assign n8814 = ~\[18376]  & ~\[18415] ;
  assign n8815 = ~\[18493]  & n8814;
  assign n8816 = ~\[17388]  & ~\[18389] ;
  assign n8817 = n8815 & n8816;
  assign n8818 = ~\[17167]  & n8817;
  assign n8819 = n8813 & n8818;
  assign n8820 = ~n3044 & n8819;
  assign n8821 = n3255 & ~n8820;
  assign n4599 = n8808 | n8821;
  always @ (posedge clock) begin
    ndout <= n274;
    ppeakb_12_12_ <= n279;
    ppeakb_1_1_ <= n283;
    ppeaka_6_6_ <= n287;
    \[4295]  <= n291;
    \[4310]  <= n296;
    ppeaks_5_5_ <= n301;
    ppeakp_10_10_ <= n305;
    \[4355]  <= n309;
    \[4370]  <= n314;
    \[4385]  <= n319;
    \[4400]  <= n324;
    \[4415]  <= n329;
    \[4430]  <= n334;
    \[4445]  <= n339;
    \[4460]  <= n344;
    \[4475]  <= n349;
    \[4490]  <= n354;
    \[4505]  <= n359;
    \[4520]  <= n364;
    \[4535]  <= n369;
    \[4550]  <= n374;
    \[4565]  <= n379;
    \[4580]  <= n384;
    \[4595]  <= n389;
    \[4610]  <= n394;
    \[4625]  <= n399;
    \[4640]  <= n404;
    \[4655]  <= n409;
    \[4670]  <= n414;
    \[4700]  <= n419;
    \[4715]  <= n424;
    \[4730]  <= n429;
    \[4745]  <= n434;
    \[4760]  <= n439;
    \[4775]  <= n444;
    \[4790]  <= n449;
    \[4805]  <= n454;
    \[4820]  <= n459;
    \[4835]  <= n464;
    \[4850]  <= n469;
    \[4865]  <= n474;
    \[4880]  <= n479;
    \[4895]  <= n484;
    \[4910]  <= n489;
    \[4925]  <= n494;
    \[4940]  <= n499;
    \[4955]  <= n504;
    \[4970]  <= n509;
    ppeakb_0_0_ <= n514;
    ppeaka_7_7_ <= n518;
    \[5015]  <= n522;
    \[5030]  <= n527;
    ppeaks_4_4_ <= n532;
    ppeakp_11_11_ <= n536;
    \[5075]  <= n540;
    \[5090]  <= n545;
    \[5105]  <= n550;
    \[5120]  <= n555;
    \[5135]  <= n560;
    \[5150]  <= n565;
    \[5165]  <= n570;
    \[5180]  <= n575;
    \[5195]  <= n580;
    \[5210]  <= n585;
    \[5225]  <= n590;
    \[5240]  <= n595;
    \[5255]  <= n600;
    \[5270]  <= n605;
    \[5285]  <= n610;
    \[5300]  <= n615;
    \[5315]  <= n620;
    \[5330]  <= n625;
    \[5345]  <= n630;
    \[5360]  <= n635;
    \[5375]  <= n640;
    \[5390]  <= n645;
    \[5405]  <= n650;
    \[5420]  <= n655;
    \[5435]  <= n660;
    \[5450]  <= n665;
    \[5465]  <= n670;
    \[5480]  <= n675;
    \[5495]  <= n680;
    \[5510]  <= n685;
    \[5525]  <= n690;
    \[5540]  <= n695;
    \[5555]  <= n700;
    \[5570]  <= n705;
    \[5600]  <= n710;
    \[5615]  <= n715;
    \[5630]  <= n720;
    \[5645]  <= n725;
    \[5660]  <= n730;
    \[5675]  <= n735;
    ppeakb_10_10_ <= n740;
    ppeaka_8_8_ <= n744;
    \[5720]  <= n748;
    ppeaks_14_14_ <= n753;
    ppeaks_7_7_ <= n757;
    ppeakp_12_12_ <= n761;
    \[5780]  <= n765;
    \[5795]  <= n770;
    \[5810]  <= n775;
    \[5825]  <= n780;
    \[5840]  <= n785;
    \[5855]  <= n790;
    \[5870]  <= n795;
    \[5885]  <= n800;
    \[5900]  <= n805;
    \[5915]  <= n810;
    \[5930]  <= n815;
    \[5945]  <= n820;
    \[5960]  <= n825;
    \[5975]  <= n830;
    \[5990]  <= n835;
    \[6005]  <= n840;
    \[6020]  <= n845;
    \[6035]  <= n850;
    \[6050]  <= n855;
    \[6065]  <= n860;
    \[6080]  <= n865;
    \[6095]  <= n870;
    \[6110]  <= n875;
    \[6125]  <= n880;
    \[6140]  <= n885;
    \[6155]  <= n890;
    \[6170]  <= n895;
    \[6185]  <= n900;
    \[6200]  <= n905;
    \[6215]  <= n910;
    \[6230]  <= n915;
    \[6245]  <= n920;
    \[6260]  <= n925;
    \[6275]  <= n930;
    \[6290]  <= n935;
    \[6305]  <= n940;
    \[6320]  <= n945;
    \[6335]  <= n950;
    \[6350]  <= n955;
    \[6365]  <= n960;
    ppeakb_11_11_ <= n965;
    ppeakb_2_2_ <= n969;
    \[6410]  <= n973;
    ppeaks_15_15_ <= n978;
    ppeaks_6_6_ <= n982;
    ppeakp_13_13_ <= n986;
    \[6470]  <= n990;
    \[6485]  <= n995;
    \[6500]  <= n1000;
    \[6515]  <= n1005;
    \[6530]  <= n1010;
    \[6545]  <= n1015;
    \[6560]  <= n1020;
    \[6575]  <= n1025;
    \[6590]  <= n1030;
    \[6605]  <= n1035;
    \[6620]  <= n1040;
    \[6635]  <= n1045;
    \[6650]  <= n1050;
    \[6665]  <= n1055;
    \[6680]  <= n1060;
    \[6695]  <= n1065;
    \[6710]  <= n1070;
    \[6725]  <= n1075;
    \[6740]  <= n1080;
    \[6755]  <= n1085;
    \[6770]  <= n1090;
    \[6785]  <= n1095;
    \[6815]  <= n1100;
    \[6830]  <= n1105;
    \[6845]  <= n1110;
    \[6860]  <= n1115;
    \[6875]  <= n1120;
    \[6890]  <= n1125;
    \[6905]  <= n1130;
    \[6920]  <= n1135;
    \[6935]  <= n1140;
    \[6950]  <= n1145;
    \[6965]  <= n1150;
    \[6980]  <= n1155;
    \[6995]  <= n1160;
    \[7010]  <= n1165;
    \[7025]  <= n1170;
    \[7055]  <= n1175;
    ppeaks_12_12_ <= n1180;
    ppeaks_1_1_ <= n1184;
    ppeakp_3_3_ <= n1188;
    \[7115]  <= n1192;
    \[7130]  <= n1197;
    \[7145]  <= n1202;
    \[7160]  <= n1207;
    \[7175]  <= n1212;
    \[7190]  <= n1217;
    \[7205]  <= n1222;
    \[7220]  <= n1227;
    \[7235]  <= n1232;
    \[7250]  <= n1237;
    \[7265]  <= n1242;
    \[7280]  <= n1247;
    \[7295]  <= n1252;
    \[7310]  <= n1257;
    \[7325]  <= n1262;
    \[7340]  <= n1267;
    \[7355]  <= n1272;
    \[7370]  <= n1277;
    \[7385]  <= n1282;
    \[7400]  <= n1287;
    \[7415]  <= n1292;
    \[7430]  <= n1297;
    \[7445]  <= n1302;
    \[7460]  <= n1307;
    \[7475]  <= n1312;
    \[7490]  <= n1317;
    \[7505]  <= n1322;
    \[7520]  <= n1327;
    \[7535]  <= n1332;
    \[7550]  <= n1337;
    \[7565]  <= n1342;
    \[7580]  <= n1347;
    \[7595]  <= n1352;
    \[7625]  <= n1357;
    \[7640]  <= n1362;
    \[7655]  <= n1367;
    \[7670]  <= n1372;
    \[7685]  <= n1377;
    ppeaks_13_13_ <= n1382;
    ppeakp_7_7_ <= n1386;
    ppeakp_2_2_ <= n1390;
    \[7745]  <= n1394;
    \[7760]  <= n1399;
    \[7775]  <= n1404;
    \[7790]  <= n1409;
    \[7805]  <= n1414;
    \[7820]  <= n1419;
    \[7835]  <= n1424;
    \[7850]  <= n1429;
    \[7865]  <= n1434;
    \[7880]  <= n1439;
    \[7895]  <= n1444;
    \[7910]  <= n1449;
    \[7925]  <= n1454;
    \[7940]  <= n1459;
    \[7955]  <= n1464;
    \[7970]  <= n1469;
    \[8000]  <= n1474;
    \[8015]  <= n1479;
    \[8030]  <= n1484;
    \[8045]  <= n1489;
    \[8060]  <= n1494;
    \[8075]  <= n1499;
    \[8090]  <= n1504;
    \[8105]  <= n1509;
    \[8120]  <= n1514;
    \[8135]  <= n1519;
    \[8150]  <= n1524;
    \[8165]  <= n1529;
    \[8180]  <= n1534;
    \[8195]  <= n1539;
    \[8210]  <= n1544;
    \[8225]  <= n1549;
    \[8240]  <= n1554;
    \[8255]  <= n1559;
    \[8285]  <= n1564;
    \[8300]  <= n1569;
    \[8315]  <= n1574;
    \[8330]  <= n1579;
    ppeaks_3_3_ <= n1584;
    ppeakp_8_8_ <= n1588;
    ppeakp_1_1_ <= n1592;
    \[8390]  <= n1596;
    \[8405]  <= n1601;
    \[8420]  <= n1606;
    \[8435]  <= n1611;
    \[8450]  <= n1616;
    \[8465]  <= n1621;
    \[8480]  <= n1626;
    \[8495]  <= n1631;
    \[8510]  <= n1636;
    \[8525]  <= n1641;
    \[8540]  <= n1646;
    \[8555]  <= n1651;
    \[8570]  <= n1656;
    \[8585]  <= n1661;
    \[8600]  <= n1666;
    \[8615]  <= n1671;
    \[8630]  <= n1676;
    \[8645]  <= n1681;
    \[8660]  <= n1686;
    \[8675]  <= n1691;
    \[8690]  <= n1696;
    \[8705]  <= n1701;
    \[8720]  <= n1706;
    \[8735]  <= n1711;
    \[8750]  <= n1716;
    \[8765]  <= n1721;
    \[8780]  <= n1726;
    \[8810]  <= n1731;
    \[8825]  <= n1736;
    \[8840]  <= n1741;
    \[8855]  <= n1746;
    \[8870]  <= n1751;
    \[8885]  <= n1756;
    \[8900]  <= n1761;
    \[8915]  <= n1766;
    \[8930]  <= n1771;
    \[8945]  <= n1776;
    \[8960]  <= n1781;
    \[8975]  <= n1786;
    ppeaks_11_11_ <= n1791;
    ppeaks_2_2_ <= n1795;
    ppeakp_9_9_ <= n1799;
    ppeakp_0_0_ <= n1803;
    \[9050]  <= n1807;
    \[9065]  <= n1812;
    \[9080]  <= n1817;
    \[9095]  <= n1822;
    \[9110]  <= n1827;
    \[9125]  <= n1832;
    \[9140]  <= n1837;
    \[9155]  <= n1842;
    \[9170]  <= n1847;
    \[9185]  <= n1852;
    \[9200]  <= n1857;
    \[9215]  <= n1862;
    \[9230]  <= n1867;
    \[9245]  <= n1872;
    \[9260]  <= n1877;
    \[9275]  <= n1882;
    \[9290]  <= n1887;
    \[9305]  <= n1892;
    \[9320]  <= n1897;
    \[9335]  <= n1902;
    \[9350]  <= n1907;
    \[9365]  <= n1912;
    \[9380]  <= n1917;
    \[9395]  <= n1922;
    \[9410]  <= n1927;
    \[9440]  <= n1932;
    \[9455]  <= n1937;
    \[9470]  <= n1942;
    \[9485]  <= n1947;
    \[9500]  <= n1952;
    \[9515]  <= n1957;
    \[9530]  <= n1962;
    \[9545]  <= n1967;
    \[9560]  <= n1972;
    \[9575]  <= n1977;
    \[9590]  <= n1982;
    \[9605]  <= n1987;
    \[9620]  <= n1992;
    \[9635]  <= n1997;
    \[9650]  <= n2002;
    \[9665]  <= n2007;
    \[9680]  <= n2012;
    ppeaki_6_6_ <= n2017;
    \[9710]  <= n2021;
    \[9725]  <= n2026;
    \[9740]  <= n2031;
    \[9770]  <= n2036;
    \[9785]  <= n2041;
    \[9800]  <= n2046;
    \[9815]  <= n2051;
    \[9830]  <= n2056;
    \[9845]  <= n2061;
    \[9860]  <= n2066;
    \[9875]  <= n2071;
    \[9890]  <= n2076;
    \[9905]  <= n2081;
    \[9920]  <= n2086;
    \[9935]  <= n2091;
    \[9950]  <= n2096;
    \[9980]  <= n2101;
    \[9995]  <= n2106;
    \[10010]  <= n2111;
    \[10025]  <= n2116;
    \[10040]  <= n2121;
    \[10055]  <= n2126;
    \[10070]  <= n2131;
    \[10085]  <= n2136;
    \[10100]  <= n2141;
    \[10115]  <= n2146;
    \[10130]  <= n2151;
    \[10145]  <= n2156;
    \[10175]  <= n2161;
    \[10190]  <= n2166;
    \[10205]  <= n2171;
    \[10220]  <= n2176;
    ppeaki_15_15_ <= n2181;
    ppeaki_4_4_ <= n2185;
    \[10265]  <= n2189;
    \[10280]  <= n2194;
    \[10310]  <= n2199;
    \[10325]  <= n2204;
    \[10340]  <= n2209;
    \[10355]  <= n2214;
    \[10370]  <= n2219;
    \[10400]  <= n2224;
    \[10415]  <= n2229;
    \[10430]  <= n2234;
    \[10445]  <= n2239;
    \[10460]  <= n2244;
    \[10475]  <= n2249;
    \[10490]  <= n2254;
    \[10505]  <= n2259;
    ppeaki_14_14_ <= n2264;
    ppeaki_5_5_ <= n2268;
    \[10550]  <= n2272;
    \[10565]  <= n2277;
    \[10580]  <= n2282;
    \[10595]  <= n2287;
    \[10610]  <= n2292;
    \[10625]  <= n2297;
    \[10655]  <= n2302;
    \[10670]  <= n2307;
    \[10685]  <= n2312;
    \[10700]  <= n2317;
    \[10715]  <= n2322;
    \[10730]  <= n2327;
    \[10745]  <= n2332;
    \[10760]  <= n2337;
    \[10775]  <= n2342;
    \[10790]  <= n2347;
    \[10805]  <= n2352;
    \[10820]  <= n2357;
    \[10850]  <= n2362;
    \[10865]  <= n2367;
    \[10880]  <= n2372;
    \[10895]  <= n2377;
    \[10925]  <= n2382;
    \[10940]  <= n2387;
    \[10955]  <= n2392;
    \[10970]  <= n2397;
    \[10985]  <= n2402;
    \[11015]  <= n2407;
    \[11030]  <= n2412;
    \[11045]  <= n2417;
    \[11060]  <= n2422;
    \[11075]  <= n2427;
    \[11090]  <= n2432;
    \[11120]  <= n2437;
    \[11135]  <= n2442;
    \[11150]  <= n2447;
    \[11165]  <= n2452;
    \[11180]  <= n2457;
    \[11195]  <= n2462;
    \[11210]  <= n2467;
    \[11225]  <= n2472;
    \[11240]  <= n2477;
    \[11255]  <= n2482;
    \[11270]  <= n2487;
    \[11285]  <= n2492;
    \[11300]  <= n2497;
    \[11315]  <= n2502;
    \[11330]  <= n2507;
    \[11345]  <= n2512;
    \[11375]  <= n2517;
    \[11390]  <= n2522;
    \[11405]  <= n2527;
    \[11420]  <= n2532;
    \[11435]  <= n2537;
    \[11450]  <= n2542;
    \[11465]  <= n2547;
    \[11480]  <= n2552;
    \[11495]  <= n2557;
    \[11510]  <= n2562;
    \[11525]  <= n2567;
    \[11540]  <= n2572;
    \[11555]  <= n2577;
    \[11570]  <= n2582;
    \[11585]  <= n2587;
    \[11600]  <= n2592;
    \[11615]  <= n2597;
    \[11630]  <= n2602;
    \[11645]  <= n2607;
    \[11660]  <= n2612;
    \[11675]  <= n2617;
    \[11690]  <= n2622;
    \[11705]  <= n2627;
    \[11720]  <= n2632;
    \[11735]  <= n2637;
    \[11750]  <= n2642;
    \[11765]  <= n2647;
    \[11780]  <= n2652;
    \[11795]  <= n2657;
    \[11810]  <= n2662;
    ppeaki_9_9_ <= n2667;
    ppeakb_14_14_ <= n2671;
    \[11885]  <= n2675;
    \[11900]  <= n2680;
    \[11915]  <= n2685;
    \[11930]  <= n2690;
    ppeaki_8_8_ <= n2695;
    ppeakb_15_15_ <= n2699;
    \[12005]  <= n2703;
    \[12020]  <= n2708;
    \[12035]  <= n2713;
    \[12050]  <= n2718;
    \[12065]  <= n2723;
    \[12080]  <= n2728;
    ppeaki_7_7_ <= n2733;
    \[12125]  <= n2737;
    \[12140]  <= n2742;
    \[12155]  <= n2747;
    \[12170]  <= n2752;
    \[12185]  <= n2757;
    \[12200]  <= n2762;
    ppeakb_13_13_ <= n2767;
    \[12245]  <= n2771;
    \[12260]  <= n2776;
    \[12275]  <= n2781;
    ppeaki_13_13_ <= n2786;
    ppeaki_2_2_ <= n2790;
    \[12335]  <= n2794;
    \[12350]  <= n2799;
    \[12365]  <= n2804;
    \[12380]  <= n2809;
    \[12395]  <= n2814;
    \[12410]  <= n2819;
    \[12425]  <= n2824;
    \[12440]  <= n2829;
    \[12455]  <= n2834;
    \[12470]  <= n2839;
    \[12485]  <= n2844;
    ppeaki_12_12_ <= n2849;
    ppeaki_3_3_ <= n2853;
    \[12545]  <= n2857;
    \[12560]  <= n2862;
    \[12575]  <= n2867;
    \[12590]  <= n2872;
    \[12605]  <= n2877;
    \[12620]  <= n2882;
    \[12635]  <= n2887;
    \[12650]  <= n2892;
    \[12665]  <= n2897;
    \[12680]  <= n2902;
    \[12695]  <= n2907;
    ppeaki_11_11_ <= n2912;
    ppeaki_0_0_ <= n2916;
    \[12770]  <= n2920;
    \[12800]  <= n2925;
    \[12815]  <= n2930;
    \[12830]  <= n2935;
    \[12845]  <= n2940;
    \[12860]  <= n2945;
    \[12875]  <= n2950;
    \[12890]  <= n2955;
    \[12905]  <= n2960;
    \[12920]  <= n2965;
    \[12935]  <= n2970;
    ppeaki_10_10_ <= n2975;
    ppeaki_1_1_ <= n2979;
    \[13010]  <= n2983;
    \[13025]  <= n2988;
    \[13040]  <= n2993;
    \[13055]  <= n2998;
    \[13070]  <= n3003;
    \[13085]  <= n3008;
    \[13100]  <= n3013;
    \[13115]  <= n3018;
    \[13130]  <= n3023;
    \[13160]  <= n3028;
    \[13175]  <= n3033;
    ppeakb_4_4_ <= n3038;
    ppeaka_9_9_ <= n3042;
    \[13220]  <= n3046;
    \[13235]  <= n3051;
    \[13250]  <= n3056;
    \[13265]  <= n3061;
    \[13280]  <= n3066;
    \[13295]  <= n3071;
    \[13310]  <= n3076;
    \[13325]  <= n3081;
    \[13340]  <= n3086;
    \[13355]  <= n3091;
    \[13370]  <= n3096;
    \[13385]  <= n3101;
    \[13400]  <= n3106;
    \[13415]  <= n3111;
    \[13430]  <= n3116;
    \[13445]  <= n3121;
    \[13460]  <= n3126;
    \[13475]  <= n3131;
    \[13490]  <= n3136;
    \[13505]  <= n3141;
    ppeakb_5_5_ <= n3146;
    \[13550]  <= n3150;
    ppeakp_6_6_ <= n3155;
    \[13580]  <= n3159;
    \[13595]  <= n3164;
    \[13610]  <= n3169;
    \[13625]  <= n3174;
    \[13640]  <= n3179;
    \[13655]  <= n3184;
    \[13670]  <= n3189;
    \[13685]  <= n3194;
    \[13700]  <= n3199;
    \[13715]  <= n3204;
    \[13730]  <= n3209;
    \[13745]  <= n3214;
    \[13775]  <= n3219;
    \[13790]  <= n3224;
    \[13805]  <= n3229;
    \[13820]  <= n3234;
    \[13835]  <= n3239;
    \[13850]  <= n3244;
    \[13865]  <= n3249;
    \[13880]  <= n3254;
    \[13895]  <= n3259;
    ppeaka_11_11_ <= n3264;
    ppeaka_0_0_ <= n3268;
    ppeakp_5_5_ <= n3272;
    \[13955]  <= n3276;
    \[13970]  <= n3281;
    \[13985]  <= n3286;
    \[14000]  <= n3291;
    \[14015]  <= n3296;
    \[14030]  <= n3301;
    \[14045]  <= n3306;
    \[14060]  <= n3311;
    \[14075]  <= n3316;
    \[14090]  <= n3321;
    \[14105]  <= n3326;
    \[14120]  <= n3331;
    \[14135]  <= n3336;
    \[14150]  <= n3341;
    \[14165]  <= n3346;
    \[14180]  <= n3351;
    \[14210]  <= n3356;
    \[14225]  <= n3361;
    \[14240]  <= n3366;
    \[14255]  <= n3371;
    \[14270]  <= n3376;
    \[14285]  <= n3381;
    ppeakb_3_3_ <= n3386;
    ppeaka_10_10_ <= n3390;
    ppeaka_1_1_ <= n3394;
    ppeakp_4_4_ <= n3398;
    \[14360]  <= n3402;
    \[14375]  <= n3407;
    \[14390]  <= n3412;
    \[14405]  <= n3417;
    \[14420]  <= n3422;
    \[14435]  <= n3427;
    \[14450]  <= n3432;
    \[14465]  <= n3437;
    \[14480]  <= n3442;
    \[14495]  <= n3447;
    \[14510]  <= n3452;
    \[14525]  <= n3457;
    \[14540]  <= n3462;
    \[14555]  <= n3467;
    \[14570]  <= n3472;
    \[14585]  <= n3477;
    \[14600]  <= n3482;
    \[14615]  <= n3487;
    \[14630]  <= n3492;
    \[14660]  <= n3497;
    \[14675]  <= n3502;
    \[14690]  <= n3507;
    \[14705]  <= n3512;
    ppeakb_8_8_ <= n3517;
    ppeaka_13_13_ <= n3521;
    ppeaka_2_2_ <= n3525;
    \[14765]  <= n3529;
    ppeaks_9_9_ <= n3534;
    ppeakp_14_14_ <= n3538;
    \[14810]  <= n3542;
    \[14825]  <= n3547;
    \[14840]  <= n3552;
    \[14855]  <= n3557;
    \[14870]  <= n3562;
    \[14885]  <= n3567;
    \[14900]  <= n3572;
    \[14915]  <= n3577;
    \[14930]  <= n3582;
    \[14960]  <= n3587;
    \[14975]  <= n3592;
    \[14990]  <= n3597;
    \[15005]  <= n3602;
    \[15020]  <= n3607;
    \[15035]  <= n3612;
    \[15050]  <= n3617;
    \[15065]  <= n3622;
    \[15080]  <= n3627;
    ppeakb_9_9_ <= n3632;
    ppeaka_12_12_ <= n3636;
    ppeaka_3_3_ <= n3640;
    \[15140]  <= n3644;
    ppeaks_8_8_ <= n3649;
    ppeakp_15_15_ <= n3653;
    \[15185]  <= n3657;
    \[15200]  <= n3662;
    \[15215]  <= n3667;
    \[15230]  <= n3672;
    \[15245]  <= n3677;
    \[15260]  <= n3682;
    \[15275]  <= n3687;
    \[15290]  <= n3692;
    \[15305]  <= n3697;
    \[15320]  <= n3702;
    \[15335]  <= n3707;
    \[15350]  <= n3712;
    \[15365]  <= n3717;
    \[15380]  <= n3722;
    \[15395]  <= n3727;
    \[15410]  <= n3732;
    \[15425]  <= n3737;
    \[15440]  <= n3742;
    ppeakb_6_6_ <= n3747;
    ppeaka_15_15_ <= n3751;
    ppeaka_4_4_ <= n3755;
    \[15500]  <= n3759;
    \[15515]  <= n3764;
    ppeaks_0_0_ <= n3769;
    \[15545]  <= n3773;
    \[15560]  <= n3778;
    \[15575]  <= n3783;
    \[15590]  <= n3788;
    \[15605]  <= n3793;
    \[15620]  <= n3798;
    \[15635]  <= n3803;
    \[15650]  <= n3808;
    \[15665]  <= n3813;
    \[15680]  <= n3818;
    \[15695]  <= n3823;
    \[15710]  <= n3828;
    \[15725]  <= n3833;
    \[15755]  <= n3838;
    \[15770]  <= n3843;
    \[15785]  <= n3848;
    ppeakb_7_7_ <= n3853;
    ppeaka_14_14_ <= n3857;
    ppeaka_5_5_ <= n3861;
    \[15845]  <= n3865;
    \[15860]  <= n3870;
    ppeaks_10_10_ <= n3875;
    \[15890]  <= n3879;
    \[15905]  <= n3884;
    \[15920]  <= n3889;
    \[15935]  <= n3894;
    \[15950]  <= n3899;
    \[15965]  <= n3904;
    \[15980]  <= n3909;
    \[15995]  <= n3914;
    \[16010]  <= n3919;
    \[16025]  <= n3924;
    \[16040]  <= n3929;
    \[16055]  <= n3934;
    \[16070]  <= n3939;
    \[16085]  <= n3944;
    \[16100]  <= n3949;
    paddress_8_8_ <= n3954;
    \[16907]  <= n3958;
    \[16920]  <= n3963;
    \[16933]  <= n3968;
    paddress_9_9_ <= n3973;
    \[16959]  <= n3977;
    \[16972]  <= n3982;
    \[16985]  <= n3987;
    \[16998]  <= n3992;
    \[17011]  <= n3997;
    \[17024]  <= n4002;
    \[17037]  <= n4007;
    \[17050]  <= n4012;
    \[17063]  <= n4017;
    \[17076]  <= n4022;
    \[17089]  <= n4027;
    \[17102]  <= n4032;
    \[17115]  <= n4037;
    \[17128]  <= n4042;
    \[17141]  <= n4047;
    \[17154]  <= n4052;
    \[17167]  <= n4057;
    \[17180]  <= n4062;
    \[17193]  <= n4067;
    \[17206]  <= n4072;
    \[17219]  <= n4077;
    \[17232]  <= n4082;
    \[17245]  <= n4087;
    \[17258]  <= n4092;
    \[17271]  <= n4097;
    \[17284]  <= n4102;
    \[17297]  <= n4107;
    \[17310]  <= n4112;
    \[17323]  <= n4117;
    \[17336]  <= n4122;
    \[17349]  <= n4127;
    \[17362]  <= n4132;
    \[17375]  <= n4137;
    \[17388]  <= n4142;
    paddress_11_11_ <= n4147;
    \[17414]  <= n4151;
    \[17427]  <= n4156;
    \[17453]  <= n4161;
    paddress_10_10_ <= n4166;
    \[17479]  <= n4170;
    \[17492]  <= n4175;
    \[17505]  <= n4180;
    \[17518]  <= n4185;
    \[17531]  <= n4190;
    \[17544]  <= n4195;
    paddress_13_13_ <= n4200;
    \[17570]  <= n4204;
    \[17583]  <= n4209;
    \[17596]  <= n4214;
    \[17609]  <= n4219;
    paddress_12_12_ <= n4224;
    \[17635]  <= n4228;
    \[17648]  <= n4233;
    \[17661]  <= n4238;
    \[17674]  <= n4243;
    paddress_15_15_ <= n4248;
    \[17700]  <= n4252;
    \[17713]  <= n4257;
    paddress_14_14_ <= n4262;
    \[17739]  <= n4266;
    \[17752]  <= n4271;
    \[17765]  <= n4276;
    \[17778]  <= n4281;
    \[17791]  <= n4286;
    \[17804]  <= n4291;
    \[17817]  <= n4296;
    pwr_0_0_ <= n4301;
    \[17843]  <= n4305;
    \[17856]  <= n4310;
    \[17869]  <= n4315;
    \[17882]  <= n4320;
    prd_0_0_ <= n4325;
    \[17908]  <= n4329;
    \[17921]  <= n4334;
    \[17934]  <= n4339;
    \[17947]  <= n4344;
    \[17960]  <= n4349;
    \[17973]  <= n4354;
    \[17986]  <= n4359;
    \[17999]  <= n4364;
    \[18012]  <= n4369;
    \[18025]  <= n4374;
    \[18038]  <= n4379;
    pdn <= n4384;
    \[18064]  <= n4388;
    \[18077]  <= n4393;
    \[18090]  <= n4398;
    \[18103]  <= n4403;
    \[18116]  <= n4408;
    \[18129]  <= n4413;
    \[18142]  <= n4418;
    \[18155]  <= n4423;
    \[18168]  <= n4428;
    \[18181]  <= n4433;
    \[18194]  <= n4438;
    \[18207]  <= n4443;
    \[18220]  <= n4448;
    \[18233]  <= n4453;
    \[18246]  <= n4458;
    paddress_0_0_ <= n4463;
    piack_0_0_ <= n4467;
    \[18285]  <= n4471;
    \[18298]  <= n4476;
    \[18311]  <= n4481;
    paddress_1_1_ <= n4486;
    \[18337]  <= n4490;
    \[18350]  <= n4495;
    \[18363]  <= n4500;
    \[18376]  <= n4505;
    \[18389]  <= n4510;
    paddress_2_2_ <= n4515;
    \[18415]  <= n4519;
    \[18428]  <= n4524;
    \[18441]  <= n4529;
    paddress_3_3_ <= n4534;
    \[18467]  <= n4538;
    \[18480]  <= n4543;
    \[18493]  <= n4548;
    \[18506]  <= n4553;
    paddress_4_4_ <= n4558;
    paddress_5_5_ <= n4562;
    \[18545]  <= n4566;
    paddress_6_6_ <= n4571;
    \[18571]  <= n4575;
    \[18584]  <= n4580;
    \[18597]  <= n4585;
    \[18610]  <= n4590;
    paddress_7_7_ <= n4595;
    \[18636]  <= n4599;
  end
endmodule


