// Benchmark "i6" written by ABC on Tue May 16 16:07:50 2017

module i6 ( 
    \V138(0) , \V96(0) , \V96(1) , \V64(13) , \V96(2) , \V64(12) ,
    \V96(3) , \V64(15) , \V96(4) , \V64(14) , \V96(5) , \V96(6) , \V96(7) ,
    \V64(11) , \V96(8) , \V64(10) , \V96(9) , \V97(0) , \V64(17) ,
    \V64(16) , \V64(19) , \V64(18) , \V64(23) , \V64(22) , \V64(25) ,
    \V64(24) , \V98(0) , \V64(21) , \V64(20) , \V64(27) , \V64(26) ,
    \V64(29) , \V64(28) , \V99(0) , \V64(31) , \V64(30) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) ,
    \V32(15) , \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) ,
    \V32(11) , \V32(10) , \V32(17) , \V32(16) , \V32(19) , \V32(18) ,
    \V32(23) , \V32(22) , \V32(25) , \V32(24) , \V32(21) , \V32(20) ,
    \V131(27) , \V131(26) , \V32(27) , \V131(29) , \V96(13) , \V32(26) ,
    \V131(28) , \V96(12) , \V32(29) , \V96(15) , \V32(28) , \V96(14) ,
    \V96(11) , \V96(10) , \V131(21) , \V131(20) , \V32(31) , \V131(23) ,
    \V131(3) , \V32(30) , \V131(22) , \V131(2) , \V131(25) , \V131(5) ,
    \V96(17) , \V131(24) , \V131(4) , \V96(16) , \V131(17) , \V96(19) ,
    \V131(16) , \V96(18) , \V131(19) , \V131(1) , \V96(23) , \V131(18) ,
    \V131(0) , \V96(22) , \V96(25) , \V96(24) , \V131(7) , \V96(21) ,
    \V131(6) , \V96(20) , \V131(11) , \V131(9) , \V131(10) , \V131(8) ,
    \V131(13) , \V131(12) , \V131(15) , \V96(27) , \V131(14) , \V96(26) ,
    \V96(29) , \V96(28) , \V64(0) , \V96(31) , \V133(1) , \V64(1) ,
    \V96(30) , \V133(0) , \V64(2) , \V64(3) , \V64(4) , \V64(5) , \V64(6) ,
    \V64(7) , \V64(8) , \V64(9) , \V134(0) , \V131(31) , \V131(30) ,
    \V138(3) , \V138(2) , \V138(4) ,
    \V198(11) , \V198(10) , \V198(13) , \V198(12) , \V198(15) , \V198(14) ,
    \V166(3) , \V166(2) , \V166(5) , \V166(4) , \V166(1) , \V166(0) ,
    \V166(7) , \V166(6) , \V166(9) , \V166(8) , \V198(31) , \V198(30) ,
    \V205(3) , \V205(2) , \V205(5) , \V205(4) , \V166(27) , \V166(26) ,
    \V198(3) , \V198(2) , \V205(1) , \V198(5) , \V205(0) , \V198(4) ,
    \V198(1) , \V198(0) , \V205(6) , \V166(21) , \V166(20) , \V166(23) ,
    \V166(22) , \V198(7) , \V166(25) , \V198(6) , \V166(24) , \V198(9) ,
    \V166(17) , \V198(8) , \V166(16) , \V166(19) , \V166(18) , \V166(11) ,
    \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) , \V198(27) ,
    \V198(26) , \V198(29) , \V198(28) , \V198(21) , \V198(20) , \V198(23) ,
    \V198(22) , \V198(25) , \V198(24) , \V198(17) , \V198(16) , \V198(19) ,
    \V198(18)   );
  input  \V138(0) , \V96(0) , \V96(1) , \V64(13) , \V96(2) , \V64(12) ,
    \V96(3) , \V64(15) , \V96(4) , \V64(14) , \V96(5) , \V96(6) , \V96(7) ,
    \V64(11) , \V96(8) , \V64(10) , \V96(9) , \V97(0) , \V64(17) ,
    \V64(16) , \V64(19) , \V64(18) , \V64(23) , \V64(22) , \V64(25) ,
    \V64(24) , \V98(0) , \V64(21) , \V64(20) , \V64(27) , \V64(26) ,
    \V64(29) , \V64(28) , \V99(0) , \V64(31) , \V64(30) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) ,
    \V32(15) , \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) ,
    \V32(11) , \V32(10) , \V32(17) , \V32(16) , \V32(19) , \V32(18) ,
    \V32(23) , \V32(22) , \V32(25) , \V32(24) , \V32(21) , \V32(20) ,
    \V131(27) , \V131(26) , \V32(27) , \V131(29) , \V96(13) , \V32(26) ,
    \V131(28) , \V96(12) , \V32(29) , \V96(15) , \V32(28) , \V96(14) ,
    \V96(11) , \V96(10) , \V131(21) , \V131(20) , \V32(31) , \V131(23) ,
    \V131(3) , \V32(30) , \V131(22) , \V131(2) , \V131(25) , \V131(5) ,
    \V96(17) , \V131(24) , \V131(4) , \V96(16) , \V131(17) , \V96(19) ,
    \V131(16) , \V96(18) , \V131(19) , \V131(1) , \V96(23) , \V131(18) ,
    \V131(0) , \V96(22) , \V96(25) , \V96(24) , \V131(7) , \V96(21) ,
    \V131(6) , \V96(20) , \V131(11) , \V131(9) , \V131(10) , \V131(8) ,
    \V131(13) , \V131(12) , \V131(15) , \V96(27) , \V131(14) , \V96(26) ,
    \V96(29) , \V96(28) , \V64(0) , \V96(31) , \V133(1) , \V64(1) ,
    \V96(30) , \V133(0) , \V64(2) , \V64(3) , \V64(4) , \V64(5) , \V64(6) ,
    \V64(7) , \V64(8) , \V64(9) , \V134(0) , \V131(31) , \V131(30) ,
    \V138(3) , \V138(2) , \V138(4) ;
  output \V198(11) , \V198(10) , \V198(13) , \V198(12) , \V198(15) ,
    \V198(14) , \V166(3) , \V166(2) , \V166(5) , \V166(4) , \V166(1) ,
    \V166(0) , \V166(7) , \V166(6) , \V166(9) , \V166(8) , \V198(31) ,
    \V198(30) , \V205(3) , \V205(2) , \V205(5) , \V205(4) , \V166(27) ,
    \V166(26) , \V198(3) , \V198(2) , \V205(1) , \V198(5) , \V205(0) ,
    \V198(4) , \V198(1) , \V198(0) , \V205(6) , \V166(21) , \V166(20) ,
    \V166(23) , \V166(22) , \V198(7) , \V166(25) , \V198(6) , \V166(24) ,
    \V198(9) , \V166(17) , \V198(8) , \V166(16) , \V166(19) , \V166(18) ,
    \V166(11) , \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) ,
    \V198(27) , \V198(26) , \V198(29) , \V198(28) , \V198(21) , \V198(20) ,
    \V198(23) , \V198(22) , \V198(25) , \V198(24) , \V198(17) , \V198(16) ,
    \V198(19) , \V198(18) ;
  wire n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n279, n280, n281, n282,
    n283, n284, n285, n287, n288, n289, n290, n291, n292, n293, n295, n296,
    n297, n298, n299, n300, n301, n303, n304, n305, n306, n307, n308, n309,
    n311, n312, n313, n314, n315, n316, n317, n319, n320, n321, n322, n323,
    n324, n325, n327, n328, n329, n330, n331, n332, n333, n335, n336, n337,
    n338, n339, n340, n341, n343, n344, n345, n346, n347, n348, n349, n351,
    n352, n353, n354, n355, n356, n357, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n396, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n432, n433, n434, n435, n436, n437, n438, n440, n441, n442, n443,
    n444, n445, n446, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n554, n555, n556, n557, n558, n559, n560, n562,
    n563, n564, n565, n566, n567, n568, n570, n571, n572, n573, n574, n575,
    n576, n578, n579, n580, n581, n582, n583, n584, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n598, n599, n600, n601, n602,
    n603, n604, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n618, n619, n620, n621, n622, n623, n624, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642,
    n643, n644, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n658, n659, n660, n661, n662, n663, n664, n666, n667, n668, n669,
    n670, n671, n672, n674, n675, n676, n677, n678, n679, n680, n682, n683,
    n684, n685, n686, n687, n688, n690, n691, n692, n693, n694, n695, n696,
    n698, n699, n700, n701, n702, n703, n704, n706, n707, n708, n709, n710,
    n711, n712, n714, n715, n716, n717, n718, n719, n720, n722, n723, n724,
    n725, n726, n727, n728, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896;
  assign n206 = \V138(2)  & ~\V138(4) ;
  assign n207 = \V138(0)  & ~\V131(7) ;
  assign n208 = \V138(2)  & n207;
  assign n209 = \V138(4)  & n208;
  assign n210 = \V138(0)  & \V131(7) ;
  assign n211 = ~\V138(2)  & n210;
  assign n212 = \V138(4)  & n211;
  assign n213 = ~\V138(0)  & \V96(7) ;
  assign n214 = ~\V138(2)  & n213;
  assign n215 = \V138(4)  & n214;
  assign n216 = ~n212 & ~n215;
  assign n217 = ~n209 & n216;
  assign \V198(11)  = n206 | ~n217;
  assign n219 = \V138(0)  & ~\V131(6) ;
  assign n220 = \V138(2)  & n219;
  assign n221 = \V138(4)  & n220;
  assign n222 = \V138(0)  & \V131(6) ;
  assign n223 = ~\V138(2)  & n222;
  assign n224 = \V138(4)  & n223;
  assign n225 = ~\V138(0)  & \V96(6) ;
  assign n226 = ~\V138(2)  & n225;
  assign n227 = \V138(4)  & n226;
  assign n228 = ~n224 & ~n227;
  assign n229 = ~n221 & n228;
  assign \V198(10)  = n206 | ~n229;
  assign n231 = \V138(0)  & ~\V131(9) ;
  assign n232 = \V138(2)  & n231;
  assign n233 = \V138(4)  & n232;
  assign n234 = \V138(0)  & \V131(9) ;
  assign n235 = ~\V138(2)  & n234;
  assign n236 = \V138(4)  & n235;
  assign n237 = ~\V138(0)  & \V96(9) ;
  assign n238 = ~\V138(2)  & n237;
  assign n239 = \V138(4)  & n238;
  assign n240 = ~n236 & ~n239;
  assign n241 = ~n233 & n240;
  assign \V198(13)  = n206 | ~n241;
  assign n243 = \V138(0)  & ~\V131(8) ;
  assign n244 = \V138(2)  & n243;
  assign n245 = \V138(4)  & n244;
  assign n246 = \V138(0)  & \V131(8) ;
  assign n247 = ~\V138(2)  & n246;
  assign n248 = \V138(4)  & n247;
  assign n249 = ~\V138(0)  & \V96(8) ;
  assign n250 = ~\V138(2)  & n249;
  assign n251 = \V138(4)  & n250;
  assign n252 = ~n248 & ~n251;
  assign n253 = ~n245 & n252;
  assign \V198(12)  = n206 | ~n253;
  assign n255 = \V138(0)  & ~\V131(11) ;
  assign n256 = \V138(2)  & n255;
  assign n257 = \V138(4)  & n256;
  assign n258 = \V138(0)  & \V131(11) ;
  assign n259 = ~\V138(2)  & n258;
  assign n260 = \V138(4)  & n259;
  assign n261 = ~\V138(0)  & \V96(11) ;
  assign n262 = ~\V138(2)  & n261;
  assign n263 = \V138(4)  & n262;
  assign n264 = ~n260 & ~n263;
  assign n265 = ~n257 & n264;
  assign \V198(15)  = n206 | ~n265;
  assign n267 = \V138(0)  & ~\V131(10) ;
  assign n268 = \V138(2)  & n267;
  assign n269 = \V138(4)  & n268;
  assign n270 = \V138(0)  & \V131(10) ;
  assign n271 = ~\V138(2)  & n270;
  assign n272 = \V138(4)  & n271;
  assign n273 = ~\V138(0)  & \V96(10) ;
  assign n274 = ~\V138(2)  & n273;
  assign n275 = \V138(4)  & n274;
  assign n276 = ~n272 & ~n275;
  assign n277 = ~n269 & n276;
  assign \V198(14)  = n206 | ~n277;
  assign n279 = ~\V64(3)  & \V138(2) ;
  assign n280 = \V138(0)  & n279;
  assign n281 = \V64(3)  & ~\V138(2) ;
  assign n282 = \V138(0)  & n281;
  assign n283 = \V32(3)  & ~\V138(2) ;
  assign n284 = ~\V138(0)  & n283;
  assign n285 = ~n282 & ~n284;
  assign \V166(3)  = n280 | ~n285;
  assign n287 = ~\V64(2)  & \V138(2) ;
  assign n288 = \V138(0)  & n287;
  assign n289 = \V64(2)  & ~\V138(2) ;
  assign n290 = \V138(0)  & n289;
  assign n291 = \V32(2)  & ~\V138(2) ;
  assign n292 = ~\V138(0)  & n291;
  assign n293 = ~n290 & ~n292;
  assign \V166(2)  = n288 | ~n293;
  assign n295 = ~\V64(5)  & \V138(2) ;
  assign n296 = \V138(0)  & n295;
  assign n297 = \V64(5)  & ~\V138(2) ;
  assign n298 = \V138(0)  & n297;
  assign n299 = \V32(5)  & ~\V138(2) ;
  assign n300 = ~\V138(0)  & n299;
  assign n301 = ~n298 & ~n300;
  assign \V166(5)  = n296 | ~n301;
  assign n303 = ~\V64(4)  & \V138(2) ;
  assign n304 = \V138(0)  & n303;
  assign n305 = \V64(4)  & ~\V138(2) ;
  assign n306 = \V138(0)  & n305;
  assign n307 = \V32(4)  & ~\V138(2) ;
  assign n308 = ~\V138(0)  & n307;
  assign n309 = ~n306 & ~n308;
  assign \V166(4)  = n304 | ~n309;
  assign n311 = ~\V64(1)  & \V138(2) ;
  assign n312 = \V138(0)  & n311;
  assign n313 = \V64(1)  & ~\V138(2) ;
  assign n314 = \V138(0)  & n313;
  assign n315 = \V32(1)  & ~\V138(2) ;
  assign n316 = ~\V138(0)  & n315;
  assign n317 = ~n314 & ~n316;
  assign \V166(1)  = n312 | ~n317;
  assign n319 = ~\V64(0)  & \V138(2) ;
  assign n320 = \V138(0)  & n319;
  assign n321 = \V64(0)  & ~\V138(2) ;
  assign n322 = \V138(0)  & n321;
  assign n323 = \V32(0)  & ~\V138(2) ;
  assign n324 = ~\V138(0)  & n323;
  assign n325 = ~n322 & ~n324;
  assign \V166(0)  = n320 | ~n325;
  assign n327 = ~\V64(7)  & \V138(2) ;
  assign n328 = \V138(0)  & n327;
  assign n329 = \V64(7)  & ~\V138(2) ;
  assign n330 = \V138(0)  & n329;
  assign n331 = \V32(7)  & ~\V138(2) ;
  assign n332 = ~\V138(0)  & n331;
  assign n333 = ~n330 & ~n332;
  assign \V166(7)  = n328 | ~n333;
  assign n335 = ~\V64(6)  & \V138(2) ;
  assign n336 = \V138(0)  & n335;
  assign n337 = \V64(6)  & ~\V138(2) ;
  assign n338 = \V138(0)  & n337;
  assign n339 = \V32(6)  & ~\V138(2) ;
  assign n340 = ~\V138(0)  & n339;
  assign n341 = ~n338 & ~n340;
  assign \V166(6)  = n336 | ~n341;
  assign n343 = ~\V64(9)  & \V138(2) ;
  assign n344 = \V138(0)  & n343;
  assign n345 = \V64(9)  & ~\V138(2) ;
  assign n346 = \V138(0)  & n345;
  assign n347 = \V32(9)  & ~\V138(2) ;
  assign n348 = ~\V138(0)  & n347;
  assign n349 = ~n346 & ~n348;
  assign \V166(9)  = n344 | ~n349;
  assign n351 = ~\V64(8)  & \V138(2) ;
  assign n352 = \V138(0)  & n351;
  assign n353 = \V64(8)  & ~\V138(2) ;
  assign n354 = \V138(0)  & n353;
  assign n355 = \V32(8)  & ~\V138(2) ;
  assign n356 = ~\V138(0)  & n355;
  assign n357 = ~n354 & ~n356;
  assign \V166(8)  = n352 | ~n357;
  assign n359 = \V138(0)  & ~\V131(27) ;
  assign n360 = \V138(2)  & n359;
  assign n361 = \V138(4)  & n360;
  assign n362 = \V138(0)  & \V131(27) ;
  assign n363 = ~\V138(2)  & n362;
  assign n364 = \V138(4)  & n363;
  assign n365 = ~\V138(0)  & \V96(27) ;
  assign n366 = ~\V138(2)  & n365;
  assign n367 = \V138(4)  & n366;
  assign n368 = ~n364 & ~n367;
  assign n369 = ~n361 & n368;
  assign \V198(31)  = n206 | ~n369;
  assign n371 = \V138(0)  & ~\V131(26) ;
  assign n372 = \V138(2)  & n371;
  assign n373 = \V138(4)  & n372;
  assign n374 = \V138(0)  & \V131(26) ;
  assign n375 = ~\V138(2)  & n374;
  assign n376 = \V138(4)  & n375;
  assign n377 = ~\V138(0)  & \V96(26) ;
  assign n378 = ~\V138(2)  & n377;
  assign n379 = \V138(4)  & n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~n373 & n380;
  assign \V198(30)  = n206 | ~n381;
  assign n383 = ~\V138(3)  & \V138(2) ;
  assign n384 = \V138(0)  & ~\V131(31) ;
  assign n385 = \V138(2)  & n384;
  assign n386 = \V138(3)  & n385;
  assign n387 = \V138(0)  & \V131(31) ;
  assign n388 = ~\V138(2)  & n387;
  assign n389 = \V138(3)  & n388;
  assign n390 = ~\V138(0)  & \V96(31) ;
  assign n391 = ~\V138(2)  & n390;
  assign n392 = \V138(3)  & n391;
  assign n393 = ~n389 & ~n392;
  assign n394 = ~n386 & n393;
  assign \V205(3)  = n383 | ~n394;
  assign n396 = \V138(0)  & ~\V131(30) ;
  assign n397 = \V138(2)  & n396;
  assign n398 = \V138(3)  & n397;
  assign n399 = \V138(0)  & \V131(30) ;
  assign n400 = ~\V138(2)  & n399;
  assign n401 = \V138(3)  & n400;
  assign n402 = ~\V138(0)  & \V96(30) ;
  assign n403 = ~\V138(2)  & n402;
  assign n404 = \V138(3)  & n403;
  assign n405 = ~n401 & ~n404;
  assign n406 = ~n398 & n405;
  assign \V205(2)  = n383 | ~n406;
  assign n408 = \V138(0)  & ~\V133(1) ;
  assign n409 = \V138(2)  & n408;
  assign n410 = \V138(3)  & n409;
  assign n411 = \V138(0)  & \V133(1) ;
  assign n412 = ~\V138(2)  & n411;
  assign n413 = \V138(3)  & n412;
  assign n414 = ~\V138(0)  & \V98(0) ;
  assign n415 = ~\V138(2)  & n414;
  assign n416 = \V138(3)  & n415;
  assign n417 = ~n413 & ~n416;
  assign n418 = ~n410 & n417;
  assign \V205(5)  = n383 | ~n418;
  assign n420 = \V138(0)  & ~\V133(0) ;
  assign n421 = \V138(2)  & n420;
  assign n422 = \V138(3)  & n421;
  assign n423 = \V138(0)  & \V133(0) ;
  assign n424 = ~\V138(2)  & n423;
  assign n425 = \V138(3)  & n424;
  assign n426 = ~\V138(0)  & \V97(0) ;
  assign n427 = ~\V138(2)  & n426;
  assign n428 = \V138(3)  & n427;
  assign n429 = ~n425 & ~n428;
  assign n430 = ~n422 & n429;
  assign \V205(4)  = n383 | ~n430;
  assign n432 = ~\V64(27)  & \V138(2) ;
  assign n433 = \V138(0)  & n432;
  assign n434 = \V64(27)  & ~\V138(2) ;
  assign n435 = \V138(0)  & n434;
  assign n436 = \V32(27)  & ~\V138(2) ;
  assign n437 = ~\V138(0)  & n436;
  assign n438 = ~n435 & ~n437;
  assign \V166(27)  = n433 | ~n438;
  assign n440 = ~\V64(26)  & \V138(2) ;
  assign n441 = \V138(0)  & n440;
  assign n442 = \V64(26)  & ~\V138(2) ;
  assign n443 = \V138(0)  & n442;
  assign n444 = \V32(26)  & ~\V138(2) ;
  assign n445 = ~\V138(0)  & n444;
  assign n446 = ~n443 & ~n445;
  assign \V166(26)  = n441 | ~n446;
  assign n448 = \V138(0)  & ~\V64(31) ;
  assign n449 = \V138(2)  & n448;
  assign n450 = \V138(4)  & n449;
  assign n451 = \V138(0)  & \V64(31) ;
  assign n452 = ~\V138(2)  & n451;
  assign n453 = \V138(4)  & n452;
  assign n454 = ~\V138(0)  & \V32(31) ;
  assign n455 = ~\V138(2)  & n454;
  assign n456 = \V138(4)  & n455;
  assign n457 = ~n453 & ~n456;
  assign n458 = ~n450 & n457;
  assign \V198(3)  = n206 | ~n458;
  assign n460 = \V138(0)  & ~\V64(30) ;
  assign n461 = \V138(2)  & n460;
  assign n462 = \V138(4)  & n461;
  assign n463 = \V138(0)  & \V64(30) ;
  assign n464 = ~\V138(2)  & n463;
  assign n465 = \V138(4)  & n464;
  assign n466 = ~\V138(0)  & \V32(30) ;
  assign n467 = ~\V138(2)  & n466;
  assign n468 = \V138(4)  & n467;
  assign n469 = ~n465 & ~n468;
  assign n470 = ~n462 & n469;
  assign \V198(2)  = n206 | ~n470;
  assign n472 = \V138(0)  & ~\V131(29) ;
  assign n473 = \V138(2)  & n472;
  assign n474 = \V138(3)  & n473;
  assign n475 = \V138(0)  & \V131(29) ;
  assign n476 = ~\V138(2)  & n475;
  assign n477 = \V138(3)  & n476;
  assign n478 = ~\V138(0)  & \V96(29) ;
  assign n479 = ~\V138(2)  & n478;
  assign n480 = \V138(3)  & n479;
  assign n481 = ~n477 & ~n480;
  assign n482 = ~n474 & n481;
  assign \V205(1)  = n383 | ~n482;
  assign n484 = \V138(0)  & ~\V131(1) ;
  assign n485 = \V138(2)  & n484;
  assign n486 = \V138(4)  & n485;
  assign n487 = \V138(0)  & \V131(1) ;
  assign n488 = ~\V138(2)  & n487;
  assign n489 = \V138(4)  & n488;
  assign n490 = ~\V138(0)  & \V96(1) ;
  assign n491 = ~\V138(2)  & n490;
  assign n492 = \V138(4)  & n491;
  assign n493 = ~n489 & ~n492;
  assign n494 = ~n486 & n493;
  assign \V198(5)  = n206 | ~n494;
  assign n496 = \V138(0)  & ~\V131(28) ;
  assign n497 = \V138(2)  & n496;
  assign n498 = \V138(3)  & n497;
  assign n499 = \V138(0)  & \V131(28) ;
  assign n500 = ~\V138(2)  & n499;
  assign n501 = \V138(3)  & n500;
  assign n502 = ~\V138(0)  & \V96(28) ;
  assign n503 = ~\V138(2)  & n502;
  assign n504 = \V138(3)  & n503;
  assign n505 = ~n501 & ~n504;
  assign n506 = ~n498 & n505;
  assign \V205(0)  = n383 | ~n506;
  assign n508 = \V138(0)  & ~\V131(0) ;
  assign n509 = \V138(2)  & n508;
  assign n510 = \V138(4)  & n509;
  assign n511 = \V138(0)  & \V131(0) ;
  assign n512 = ~\V138(2)  & n511;
  assign n513 = \V138(4)  & n512;
  assign n514 = ~\V138(0)  & \V96(0) ;
  assign n515 = ~\V138(2)  & n514;
  assign n516 = \V138(4)  & n515;
  assign n517 = ~n513 & ~n516;
  assign n518 = ~n510 & n517;
  assign \V198(4)  = n206 | ~n518;
  assign n520 = \V138(0)  & ~\V64(29) ;
  assign n521 = \V138(2)  & n520;
  assign n522 = \V138(4)  & n521;
  assign n523 = \V138(0)  & \V64(29) ;
  assign n524 = ~\V138(2)  & n523;
  assign n525 = \V138(4)  & n524;
  assign n526 = ~\V138(0)  & \V32(29) ;
  assign n527 = ~\V138(2)  & n526;
  assign n528 = \V138(4)  & n527;
  assign n529 = ~n525 & ~n528;
  assign n530 = ~n522 & n529;
  assign \V198(1)  = n206 | ~n530;
  assign n532 = \V138(0)  & ~\V64(28) ;
  assign n533 = \V138(2)  & n532;
  assign n534 = \V138(4)  & n533;
  assign n535 = \V138(0)  & \V64(28) ;
  assign n536 = ~\V138(2)  & n535;
  assign n537 = \V138(4)  & n536;
  assign n538 = ~\V138(0)  & \V32(28) ;
  assign n539 = ~\V138(2)  & n538;
  assign n540 = \V138(4)  & n539;
  assign n541 = ~n537 & ~n540;
  assign n542 = ~n534 & n541;
  assign \V198(0)  = n206 | ~n542;
  assign n544 = \V138(0)  & \V134(0) ;
  assign n545 = \V138(2)  & n544;
  assign n546 = \V138(3)  & n545;
  assign n547 = ~\V138(2)  & n544;
  assign n548 = \V138(3)  & n547;
  assign n549 = ~\V138(0)  & \V99(0) ;
  assign n550 = ~\V138(2)  & n549;
  assign n551 = \V138(3)  & n550;
  assign n552 = ~n548 & ~n551;
  assign \V205(6)  = n546 | ~n552;
  assign n554 = ~\V64(21)  & \V138(2) ;
  assign n555 = \V138(0)  & n554;
  assign n556 = \V64(21)  & ~\V138(2) ;
  assign n557 = \V138(0)  & n556;
  assign n558 = \V32(21)  & ~\V138(2) ;
  assign n559 = ~\V138(0)  & n558;
  assign n560 = ~n557 & ~n559;
  assign \V166(21)  = n555 | ~n560;
  assign n562 = ~\V64(20)  & \V138(2) ;
  assign n563 = \V138(0)  & n562;
  assign n564 = \V64(20)  & ~\V138(2) ;
  assign n565 = \V138(0)  & n564;
  assign n566 = \V32(20)  & ~\V138(2) ;
  assign n567 = ~\V138(0)  & n566;
  assign n568 = ~n565 & ~n567;
  assign \V166(20)  = n563 | ~n568;
  assign n570 = ~\V64(23)  & \V138(2) ;
  assign n571 = \V138(0)  & n570;
  assign n572 = \V64(23)  & ~\V138(2) ;
  assign n573 = \V138(0)  & n572;
  assign n574 = \V32(23)  & ~\V138(2) ;
  assign n575 = ~\V138(0)  & n574;
  assign n576 = ~n573 & ~n575;
  assign \V166(23)  = n571 | ~n576;
  assign n578 = ~\V64(22)  & \V138(2) ;
  assign n579 = \V138(0)  & n578;
  assign n580 = \V64(22)  & ~\V138(2) ;
  assign n581 = \V138(0)  & n580;
  assign n582 = \V32(22)  & ~\V138(2) ;
  assign n583 = ~\V138(0)  & n582;
  assign n584 = ~n581 & ~n583;
  assign \V166(22)  = n579 | ~n584;
  assign n586 = \V138(0)  & ~\V131(3) ;
  assign n587 = \V138(2)  & n586;
  assign n588 = \V138(4)  & n587;
  assign n589 = \V138(0)  & \V131(3) ;
  assign n590 = ~\V138(2)  & n589;
  assign n591 = \V138(4)  & n590;
  assign n592 = ~\V138(0)  & \V96(3) ;
  assign n593 = ~\V138(2)  & n592;
  assign n594 = \V138(4)  & n593;
  assign n595 = ~n591 & ~n594;
  assign n596 = ~n588 & n595;
  assign \V198(7)  = n206 | ~n596;
  assign n598 = ~\V64(25)  & \V138(2) ;
  assign n599 = \V138(0)  & n598;
  assign n600 = \V64(25)  & ~\V138(2) ;
  assign n601 = \V138(0)  & n600;
  assign n602 = \V32(25)  & ~\V138(2) ;
  assign n603 = ~\V138(0)  & n602;
  assign n604 = ~n601 & ~n603;
  assign \V166(25)  = n599 | ~n604;
  assign n606 = \V138(0)  & ~\V131(2) ;
  assign n607 = \V138(2)  & n606;
  assign n608 = \V138(4)  & n607;
  assign n609 = \V138(0)  & \V131(2) ;
  assign n610 = ~\V138(2)  & n609;
  assign n611 = \V138(4)  & n610;
  assign n612 = ~\V138(0)  & \V96(2) ;
  assign n613 = ~\V138(2)  & n612;
  assign n614 = \V138(4)  & n613;
  assign n615 = ~n611 & ~n614;
  assign n616 = ~n608 & n615;
  assign \V198(6)  = n206 | ~n616;
  assign n618 = ~\V64(24)  & \V138(2) ;
  assign n619 = \V138(0)  & n618;
  assign n620 = \V64(24)  & ~\V138(2) ;
  assign n621 = \V138(0)  & n620;
  assign n622 = \V32(24)  & ~\V138(2) ;
  assign n623 = ~\V138(0)  & n622;
  assign n624 = ~n621 & ~n623;
  assign \V166(24)  = n619 | ~n624;
  assign n626 = \V138(0)  & ~\V131(5) ;
  assign n627 = \V138(2)  & n626;
  assign n628 = \V138(4)  & n627;
  assign n629 = \V138(0)  & \V131(5) ;
  assign n630 = ~\V138(2)  & n629;
  assign n631 = \V138(4)  & n630;
  assign n632 = ~\V138(0)  & \V96(5) ;
  assign n633 = ~\V138(2)  & n632;
  assign n634 = \V138(4)  & n633;
  assign n635 = ~n631 & ~n634;
  assign n636 = ~n628 & n635;
  assign \V198(9)  = n206 | ~n636;
  assign n638 = ~\V64(17)  & \V138(2) ;
  assign n639 = \V138(0)  & n638;
  assign n640 = \V64(17)  & ~\V138(2) ;
  assign n641 = \V138(0)  & n640;
  assign n642 = \V32(17)  & ~\V138(2) ;
  assign n643 = ~\V138(0)  & n642;
  assign n644 = ~n641 & ~n643;
  assign \V166(17)  = n639 | ~n644;
  assign n646 = \V138(0)  & ~\V131(4) ;
  assign n647 = \V138(2)  & n646;
  assign n648 = \V138(4)  & n647;
  assign n649 = \V138(0)  & \V131(4) ;
  assign n650 = ~\V138(2)  & n649;
  assign n651 = \V138(4)  & n650;
  assign n652 = ~\V138(0)  & \V96(4) ;
  assign n653 = ~\V138(2)  & n652;
  assign n654 = \V138(4)  & n653;
  assign n655 = ~n651 & ~n654;
  assign n656 = ~n648 & n655;
  assign \V198(8)  = n206 | ~n656;
  assign n658 = ~\V64(16)  & \V138(2) ;
  assign n659 = \V138(0)  & n658;
  assign n660 = \V64(16)  & ~\V138(2) ;
  assign n661 = \V138(0)  & n660;
  assign n662 = \V32(16)  & ~\V138(2) ;
  assign n663 = ~\V138(0)  & n662;
  assign n664 = ~n661 & ~n663;
  assign \V166(16)  = n659 | ~n664;
  assign n666 = ~\V64(19)  & \V138(2) ;
  assign n667 = \V138(0)  & n666;
  assign n668 = \V64(19)  & ~\V138(2) ;
  assign n669 = \V138(0)  & n668;
  assign n670 = \V32(19)  & ~\V138(2) ;
  assign n671 = ~\V138(0)  & n670;
  assign n672 = ~n669 & ~n671;
  assign \V166(19)  = n667 | ~n672;
  assign n674 = ~\V64(18)  & \V138(2) ;
  assign n675 = \V138(0)  & n674;
  assign n676 = \V64(18)  & ~\V138(2) ;
  assign n677 = \V138(0)  & n676;
  assign n678 = \V32(18)  & ~\V138(2) ;
  assign n679 = ~\V138(0)  & n678;
  assign n680 = ~n677 & ~n679;
  assign \V166(18)  = n675 | ~n680;
  assign n682 = ~\V64(11)  & \V138(2) ;
  assign n683 = \V138(0)  & n682;
  assign n684 = \V64(11)  & ~\V138(2) ;
  assign n685 = \V138(0)  & n684;
  assign n686 = \V32(11)  & ~\V138(2) ;
  assign n687 = ~\V138(0)  & n686;
  assign n688 = ~n685 & ~n687;
  assign \V166(11)  = n683 | ~n688;
  assign n690 = ~\V64(10)  & \V138(2) ;
  assign n691 = \V138(0)  & n690;
  assign n692 = \V64(10)  & ~\V138(2) ;
  assign n693 = \V138(0)  & n692;
  assign n694 = \V32(10)  & ~\V138(2) ;
  assign n695 = ~\V138(0)  & n694;
  assign n696 = ~n693 & ~n695;
  assign \V166(10)  = n691 | ~n696;
  assign n698 = ~\V64(13)  & \V138(2) ;
  assign n699 = \V138(0)  & n698;
  assign n700 = \V64(13)  & ~\V138(2) ;
  assign n701 = \V138(0)  & n700;
  assign n702 = \V32(13)  & ~\V138(2) ;
  assign n703 = ~\V138(0)  & n702;
  assign n704 = ~n701 & ~n703;
  assign \V166(13)  = n699 | ~n704;
  assign n706 = ~\V64(12)  & \V138(2) ;
  assign n707 = \V138(0)  & n706;
  assign n708 = \V64(12)  & ~\V138(2) ;
  assign n709 = \V138(0)  & n708;
  assign n710 = \V32(12)  & ~\V138(2) ;
  assign n711 = ~\V138(0)  & n710;
  assign n712 = ~n709 & ~n711;
  assign \V166(12)  = n707 | ~n712;
  assign n714 = ~\V64(15)  & \V138(2) ;
  assign n715 = \V138(0)  & n714;
  assign n716 = \V64(15)  & ~\V138(2) ;
  assign n717 = \V138(0)  & n716;
  assign n718 = \V32(15)  & ~\V138(2) ;
  assign n719 = ~\V138(0)  & n718;
  assign n720 = ~n717 & ~n719;
  assign \V166(15)  = n715 | ~n720;
  assign n722 = ~\V64(14)  & \V138(2) ;
  assign n723 = \V138(0)  & n722;
  assign n724 = \V64(14)  & ~\V138(2) ;
  assign n725 = \V138(0)  & n724;
  assign n726 = \V32(14)  & ~\V138(2) ;
  assign n727 = ~\V138(0)  & n726;
  assign n728 = ~n725 & ~n727;
  assign \V166(14)  = n723 | ~n728;
  assign n730 = \V138(0)  & ~\V131(23) ;
  assign n731 = \V138(2)  & n730;
  assign n732 = \V138(4)  & n731;
  assign n733 = \V138(0)  & \V131(23) ;
  assign n734 = ~\V138(2)  & n733;
  assign n735 = \V138(4)  & n734;
  assign n736 = ~\V138(0)  & \V96(23) ;
  assign n737 = ~\V138(2)  & n736;
  assign n738 = \V138(4)  & n737;
  assign n739 = ~n735 & ~n738;
  assign n740 = ~n732 & n739;
  assign \V198(27)  = n206 | ~n740;
  assign n742 = \V138(0)  & ~\V131(22) ;
  assign n743 = \V138(2)  & n742;
  assign n744 = \V138(4)  & n743;
  assign n745 = \V138(0)  & \V131(22) ;
  assign n746 = ~\V138(2)  & n745;
  assign n747 = \V138(4)  & n746;
  assign n748 = ~\V138(0)  & \V96(22) ;
  assign n749 = ~\V138(2)  & n748;
  assign n750 = \V138(4)  & n749;
  assign n751 = ~n747 & ~n750;
  assign n752 = ~n744 & n751;
  assign \V198(26)  = n206 | ~n752;
  assign n754 = \V138(0)  & ~\V131(25) ;
  assign n755 = \V138(2)  & n754;
  assign n756 = \V138(4)  & n755;
  assign n757 = \V138(0)  & \V131(25) ;
  assign n758 = ~\V138(2)  & n757;
  assign n759 = \V138(4)  & n758;
  assign n760 = ~\V138(0)  & \V96(25) ;
  assign n761 = ~\V138(2)  & n760;
  assign n762 = \V138(4)  & n761;
  assign n763 = ~n759 & ~n762;
  assign n764 = ~n756 & n763;
  assign \V198(29)  = n206 | ~n764;
  assign n766 = \V138(0)  & ~\V131(24) ;
  assign n767 = \V138(2)  & n766;
  assign n768 = \V138(4)  & n767;
  assign n769 = \V138(0)  & \V131(24) ;
  assign n770 = ~\V138(2)  & n769;
  assign n771 = \V138(4)  & n770;
  assign n772 = ~\V138(0)  & \V96(24) ;
  assign n773 = ~\V138(2)  & n772;
  assign n774 = \V138(4)  & n773;
  assign n775 = ~n771 & ~n774;
  assign n776 = ~n768 & n775;
  assign \V198(28)  = n206 | ~n776;
  assign n778 = \V138(0)  & ~\V131(17) ;
  assign n779 = \V138(2)  & n778;
  assign n780 = \V138(4)  & n779;
  assign n781 = \V138(0)  & \V131(17) ;
  assign n782 = ~\V138(2)  & n781;
  assign n783 = \V138(4)  & n782;
  assign n784 = ~\V138(0)  & \V96(17) ;
  assign n785 = ~\V138(2)  & n784;
  assign n786 = \V138(4)  & n785;
  assign n787 = ~n783 & ~n786;
  assign n788 = ~n780 & n787;
  assign \V198(21)  = n206 | ~n788;
  assign n790 = \V138(0)  & ~\V131(16) ;
  assign n791 = \V138(2)  & n790;
  assign n792 = \V138(4)  & n791;
  assign n793 = \V138(0)  & \V131(16) ;
  assign n794 = ~\V138(2)  & n793;
  assign n795 = \V138(4)  & n794;
  assign n796 = ~\V138(0)  & \V96(16) ;
  assign n797 = ~\V138(2)  & n796;
  assign n798 = \V138(4)  & n797;
  assign n799 = ~n795 & ~n798;
  assign n800 = ~n792 & n799;
  assign \V198(20)  = n206 | ~n800;
  assign n802 = \V138(0)  & ~\V131(19) ;
  assign n803 = \V138(2)  & n802;
  assign n804 = \V138(4)  & n803;
  assign n805 = \V138(0)  & \V131(19) ;
  assign n806 = ~\V138(2)  & n805;
  assign n807 = \V138(4)  & n806;
  assign n808 = ~\V138(0)  & \V96(19) ;
  assign n809 = ~\V138(2)  & n808;
  assign n810 = \V138(4)  & n809;
  assign n811 = ~n807 & ~n810;
  assign n812 = ~n804 & n811;
  assign \V198(23)  = n206 | ~n812;
  assign n814 = \V138(0)  & ~\V131(18) ;
  assign n815 = \V138(2)  & n814;
  assign n816 = \V138(4)  & n815;
  assign n817 = \V138(0)  & \V131(18) ;
  assign n818 = ~\V138(2)  & n817;
  assign n819 = \V138(4)  & n818;
  assign n820 = ~\V138(0)  & \V96(18) ;
  assign n821 = ~\V138(2)  & n820;
  assign n822 = \V138(4)  & n821;
  assign n823 = ~n819 & ~n822;
  assign n824 = ~n816 & n823;
  assign \V198(22)  = n206 | ~n824;
  assign n826 = \V138(0)  & ~\V131(21) ;
  assign n827 = \V138(2)  & n826;
  assign n828 = \V138(4)  & n827;
  assign n829 = \V138(0)  & \V131(21) ;
  assign n830 = ~\V138(2)  & n829;
  assign n831 = \V138(4)  & n830;
  assign n832 = ~\V138(0)  & \V96(21) ;
  assign n833 = ~\V138(2)  & n832;
  assign n834 = \V138(4)  & n833;
  assign n835 = ~n831 & ~n834;
  assign n836 = ~n828 & n835;
  assign \V198(25)  = n206 | ~n836;
  assign n838 = \V138(0)  & ~\V131(20) ;
  assign n839 = \V138(2)  & n838;
  assign n840 = \V138(4)  & n839;
  assign n841 = \V138(0)  & \V131(20) ;
  assign n842 = ~\V138(2)  & n841;
  assign n843 = \V138(4)  & n842;
  assign n844 = ~\V138(0)  & \V96(20) ;
  assign n845 = ~\V138(2)  & n844;
  assign n846 = \V138(4)  & n845;
  assign n847 = ~n843 & ~n846;
  assign n848 = ~n840 & n847;
  assign \V198(24)  = n206 | ~n848;
  assign n850 = \V138(0)  & ~\V131(13) ;
  assign n851 = \V138(2)  & n850;
  assign n852 = \V138(4)  & n851;
  assign n853 = \V138(0)  & \V131(13) ;
  assign n854 = ~\V138(2)  & n853;
  assign n855 = \V138(4)  & n854;
  assign n856 = ~\V138(0)  & \V96(13) ;
  assign n857 = ~\V138(2)  & n856;
  assign n858 = \V138(4)  & n857;
  assign n859 = ~n855 & ~n858;
  assign n860 = ~n852 & n859;
  assign \V198(17)  = n206 | ~n860;
  assign n862 = \V138(0)  & ~\V131(12) ;
  assign n863 = \V138(2)  & n862;
  assign n864 = \V138(4)  & n863;
  assign n865 = \V138(0)  & \V131(12) ;
  assign n866 = ~\V138(2)  & n865;
  assign n867 = \V138(4)  & n866;
  assign n868 = ~\V138(0)  & \V96(12) ;
  assign n869 = ~\V138(2)  & n868;
  assign n870 = \V138(4)  & n869;
  assign n871 = ~n867 & ~n870;
  assign n872 = ~n864 & n871;
  assign \V198(16)  = n206 | ~n872;
  assign n874 = \V138(0)  & ~\V131(15) ;
  assign n875 = \V138(2)  & n874;
  assign n876 = \V138(4)  & n875;
  assign n877 = \V138(0)  & \V131(15) ;
  assign n878 = ~\V138(2)  & n877;
  assign n879 = \V138(4)  & n878;
  assign n880 = ~\V138(0)  & \V96(15) ;
  assign n881 = ~\V138(2)  & n880;
  assign n882 = \V138(4)  & n881;
  assign n883 = ~n879 & ~n882;
  assign n884 = ~n876 & n883;
  assign \V198(19)  = n206 | ~n884;
  assign n886 = \V138(0)  & ~\V131(14) ;
  assign n887 = \V138(2)  & n886;
  assign n888 = \V138(4)  & n887;
  assign n889 = \V138(0)  & \V131(14) ;
  assign n890 = ~\V138(2)  & n889;
  assign n891 = \V138(4)  & n890;
  assign n892 = ~\V138(0)  & \V96(14) ;
  assign n893 = ~\V138(2)  & n892;
  assign n894 = \V138(4)  & n893;
  assign n895 = ~n891 & ~n894;
  assign n896 = ~n888 & n895;
  assign \V198(18)  = n206 | ~n896;
endmodule


