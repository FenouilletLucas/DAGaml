// Benchmark "i8" written by ABC on Tue May 16 16:07:50 2017

module i8 ( 
    \V116(12) , \V133(5) , \V116(15) , \V133(4) , \V116(14) , \V133(1) ,
    \V133(0) , \V133(7) , \V133(6) , \V116(3) , \V133(9) , \V116(2) ,
    \V133(8) , \V116(5) , \V116(4) , \V116(1) , \V116(0) , \V116(7) ,
    \V116(6) , \V116(9) , \V116(8) , \V116(31) , \V116(30) , \V118(1) ,
    \V118(0) , \V84(13) , \V84(12) , \V84(15) , \V84(14) , \V15(13) ,
    \V15(12) , \V84(11) , \V84(10) , \V15(14) , \V15(11) , \V15(10) ,
    \V84(17) , \V84(16) , \V84(19) , \V84(18) , \V84(23) , \V84(22) ,
    \V84(25) , \V84(24) , \V84(21) , \V84(20) , \V84(27) , \V84(26) ,
    \V84(29) , \V84(28) , \V47(13) , \V47(12) , \V47(15) , \V47(14) ,
    \V84(31) , \V84(30) , \V47(11) , \V47(10) , \V47(17) , \V47(16) ,
    \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V47(25) , \V47(24) ,
    \V122(0) , \V47(21) , \V47(20) , \V47(27) , \V47(26) , \V47(29) ,
    \V47(28) , \V84(0) , \V84(1) , \V47(31) , \V84(2) , \V47(30) ,
    \V84(3) , \V84(4) , \V84(5) , \V84(6) , \V84(7) , \V84(8) , \V84(9) ,
    \V48(0) , \V50(0) , \V52(0) , \V133(10) , \V119(0) , \V47(0) ,
    \V47(1) , \V47(2) , \V47(3) , \V47(4) , \V47(5) , \V47(6) , \V47(7) ,
    \V47(8) , \V47(9) , \V49(0) , \V121(17) , \V121(16) , \V51(0) ,
    \V116(27) , \V116(26) , \V116(29) , \V116(28) , \V15(0) , \V15(1) ,
    \V15(2) , \V15(3) , \V15(4) , \V15(5) , \V15(6) , \V116(21) , \V15(7) ,
    \V116(20) , \V15(8) , \V116(23) , \V15(9) , \V116(22) , \V116(25) ,
    \V116(24) , \V116(17) , \V116(16) , \V116(19) , \V116(18) , \V116(11) ,
    \V116(10) , \V133(3) , \V116(13) , \V133(2) ,
    \V212(3) , \V212(2) , \V212(5) , \V212(4) , \V212(1) , \V212(0) ,
    \V212(7) , \V212(6) , \V212(9) , \V212(8) , \V214(0) , \V143(0) ,
    \V145(1) , \V145(0) , \V149(2) , \V149(1) , \V149(0) , \V134(0) ,
    \V136(1) , \V136(0) , \V165(11) , \V197(3) , \V165(10) , \V197(2) ,
    \V165(13) , \V197(5) , \V165(12) , \V197(4) , \V197(27) , \V197(26) ,
    \V165(14) , \V197(29) , \V197(1) , \V197(28) , \V197(0) , \V197(7) ,
    \V197(6) , \V197(21) , \V197(9) , \V197(20) , \V197(8) , \V197(23) ,
    \V197(22) , \V197(25) , \V197(24) , \V213(0) , \V197(17) , \V197(16) ,
    \V197(19) , \V197(18) , \V197(11) , \V197(10) , \V197(13) , \V197(12) ,
    \V197(15) , \V197(14) , \V142(3) , \V142(2) , \V142(5) , \V142(4) ,
    \V197(31) , \V142(1) , \V197(30) , \V142(0) , \V165(3) , \V212(11) ,
    \V165(2) , \V212(10) , \V165(5) , \V212(13) , \V165(4) , \V212(12) ,
    \V146(0) , \V212(14) , \V165(1) , \V165(0) , \V165(7) , \V165(6) ,
    \V165(9) , \V165(8) , \V150(0)   );
  input  \V116(12) , \V133(5) , \V116(15) , \V133(4) , \V116(14) ,
    \V133(1) , \V133(0) , \V133(7) , \V133(6) , \V116(3) , \V133(9) ,
    \V116(2) , \V133(8) , \V116(5) , \V116(4) , \V116(1) , \V116(0) ,
    \V116(7) , \V116(6) , \V116(9) , \V116(8) , \V116(31) , \V116(30) ,
    \V118(1) , \V118(0) , \V84(13) , \V84(12) , \V84(15) , \V84(14) ,
    \V15(13) , \V15(12) , \V84(11) , \V84(10) , \V15(14) , \V15(11) ,
    \V15(10) , \V84(17) , \V84(16) , \V84(19) , \V84(18) , \V84(23) ,
    \V84(22) , \V84(25) , \V84(24) , \V84(21) , \V84(20) , \V84(27) ,
    \V84(26) , \V84(29) , \V84(28) , \V47(13) , \V47(12) , \V47(15) ,
    \V47(14) , \V84(31) , \V84(30) , \V47(11) , \V47(10) , \V47(17) ,
    \V47(16) , \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V47(25) ,
    \V47(24) , \V122(0) , \V47(21) , \V47(20) , \V47(27) , \V47(26) ,
    \V47(29) , \V47(28) , \V84(0) , \V84(1) , \V47(31) , \V84(2) ,
    \V47(30) , \V84(3) , \V84(4) , \V84(5) , \V84(6) , \V84(7) , \V84(8) ,
    \V84(9) , \V48(0) , \V50(0) , \V52(0) , \V133(10) , \V119(0) ,
    \V47(0) , \V47(1) , \V47(2) , \V47(3) , \V47(4) , \V47(5) , \V47(6) ,
    \V47(7) , \V47(8) , \V47(9) , \V49(0) , \V121(17) , \V121(16) ,
    \V51(0) , \V116(27) , \V116(26) , \V116(29) , \V116(28) , \V15(0) ,
    \V15(1) , \V15(2) , \V15(3) , \V15(4) , \V15(5) , \V15(6) , \V116(21) ,
    \V15(7) , \V116(20) , \V15(8) , \V116(23) , \V15(9) , \V116(22) ,
    \V116(25) , \V116(24) , \V116(17) , \V116(16) , \V116(19) , \V116(18) ,
    \V116(11) , \V116(10) , \V133(3) , \V116(13) , \V133(2) ;
  output \V212(3) , \V212(2) , \V212(5) , \V212(4) , \V212(1) , \V212(0) ,
    \V212(7) , \V212(6) , \V212(9) , \V212(8) , \V214(0) , \V143(0) ,
    \V145(1) , \V145(0) , \V149(2) , \V149(1) , \V149(0) , \V134(0) ,
    \V136(1) , \V136(0) , \V165(11) , \V197(3) , \V165(10) , \V197(2) ,
    \V165(13) , \V197(5) , \V165(12) , \V197(4) , \V197(27) , \V197(26) ,
    \V165(14) , \V197(29) , \V197(1) , \V197(28) , \V197(0) , \V197(7) ,
    \V197(6) , \V197(21) , \V197(9) , \V197(20) , \V197(8) , \V197(23) ,
    \V197(22) , \V197(25) , \V197(24) , \V213(0) , \V197(17) , \V197(16) ,
    \V197(19) , \V197(18) , \V197(11) , \V197(10) , \V197(13) , \V197(12) ,
    \V197(15) , \V197(14) , \V142(3) , \V142(2) , \V142(5) , \V142(4) ,
    \V197(31) , \V142(1) , \V197(30) , \V142(0) , \V165(3) , \V212(11) ,
    \V165(2) , \V212(10) , \V165(5) , \V212(13) , \V165(4) , \V212(12) ,
    \V146(0) , \V212(14) , \V165(1) , \V165(0) , \V165(7) , \V165(6) ,
    \V165(9) , \V165(8) , \V150(0) ;
  wire n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n391,
    n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
    n2382, n2383, n2384, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2708, n2709, n2710, n2711,
    n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523;
  assign n215 = ~\V133(1)  & ~\V133(9) ;
  assign n216 = ~\V133(2)  & n215;
  assign n217 = ~\V133(6)  & n216;
  assign n218 = ~\V133(4)  & n217;
  assign n219 = ~\V133(5)  & n218;
  assign n220 = \V133(7)  & n216;
  assign n221 = ~\V133(1)  & ~\V118(1) ;
  assign n222 = ~\V133(2)  & n221;
  assign n223 = ~\V118(0)  & n222;
  assign n224 = ~\V133(10)  & n223;
  assign n225 = \V133(5)  & n224;
  assign n226 = ~\V133(9)  & n225;
  assign n227 = ~\V133(7)  & n226;
  assign n228 = \V116(3)  & ~n227;
  assign n229 = ~n220 & n228;
  assign n230 = ~n219 & n229;
  assign n231 = ~\V133(10)  & n230;
  assign n232 = \V133(9)  & n231;
  assign n233 = ~\V133(10)  & n232;
  assign n234 = ~n220 & n227;
  assign n235 = ~n219 & n234;
  assign n236 = ~\V133(10)  & n235;
  assign n237 = \V84(20)  & ~n220;
  assign n238 = ~n219 & n237;
  assign n239 = \V133(10)  & n238;
  assign n240 = \V84(20)  & n220;
  assign n241 = ~n219 & n240;
  assign n242 = \V84(20)  & n219;
  assign n243 = ~n241 & ~n242;
  assign n244 = ~n239 & n243;
  assign n245 = ~n236 & n244;
  assign \V212(3)  = n233 | ~n245;
  assign n247 = \V116(2)  & ~n227;
  assign n248 = ~n220 & n247;
  assign n249 = ~n219 & n248;
  assign n250 = ~\V133(10)  & n249;
  assign n251 = \V133(9)  & n250;
  assign n252 = ~\V133(10)  & n251;
  assign n253 = \V84(19)  & ~n220;
  assign n254 = ~n219 & n253;
  assign n255 = \V133(10)  & n254;
  assign n256 = \V84(19)  & n220;
  assign n257 = ~n219 & n256;
  assign n258 = \V84(19)  & n219;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~n255 & n259;
  assign n261 = ~n236 & n260;
  assign \V212(2)  = n252 | ~n261;
  assign n263 = \V116(5)  & ~n227;
  assign n264 = ~n220 & n263;
  assign n265 = ~n219 & n264;
  assign n266 = ~\V133(10)  & n265;
  assign n267 = \V133(9)  & n266;
  assign n268 = ~\V133(10)  & n267;
  assign n269 = \V84(22)  & ~n220;
  assign n270 = ~n219 & n269;
  assign n271 = \V133(10)  & n270;
  assign n272 = \V84(22)  & n220;
  assign n273 = ~n219 & n272;
  assign n274 = \V84(22)  & n219;
  assign n275 = ~n273 & ~n274;
  assign n276 = ~n271 & n275;
  assign n277 = ~n236 & n276;
  assign \V212(5)  = n268 | ~n277;
  assign n279 = \V116(4)  & ~n227;
  assign n280 = ~n220 & n279;
  assign n281 = ~n219 & n280;
  assign n282 = ~\V133(10)  & n281;
  assign n283 = \V133(9)  & n282;
  assign n284 = ~\V133(10)  & n283;
  assign n285 = \V84(21)  & ~n220;
  assign n286 = ~n219 & n285;
  assign n287 = \V133(10)  & n286;
  assign n288 = \V84(21)  & n220;
  assign n289 = ~n219 & n288;
  assign n290 = \V84(21)  & n219;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n287 & n291;
  assign n293 = ~n236 & n292;
  assign \V212(4)  = n284 | ~n293;
  assign n295 = \V116(1)  & ~n227;
  assign n296 = ~n220 & n295;
  assign n297 = ~n219 & n296;
  assign n298 = ~\V133(10)  & n297;
  assign n299 = \V133(9)  & n298;
  assign n300 = ~\V133(10)  & n299;
  assign n301 = \V84(18)  & ~n220;
  assign n302 = ~n219 & n301;
  assign n303 = \V133(10)  & n302;
  assign n304 = \V84(18)  & n220;
  assign n305 = ~n219 & n304;
  assign n306 = \V84(18)  & n219;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~n303 & n307;
  assign n309 = ~n236 & n308;
  assign \V212(1)  = n300 | ~n309;
  assign n311 = \V116(0)  & ~n227;
  assign n312 = ~n220 & n311;
  assign n313 = ~n219 & n312;
  assign n314 = ~\V133(10)  & n313;
  assign n315 = \V133(9)  & n314;
  assign n316 = ~\V133(10)  & n315;
  assign n317 = \V84(17)  & ~n220;
  assign n318 = ~n219 & n317;
  assign n319 = \V133(10)  & n318;
  assign n320 = \V84(17)  & n220;
  assign n321 = ~n219 & n320;
  assign n322 = \V84(17)  & n219;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~n319 & n323;
  assign n325 = ~n236 & n324;
  assign \V212(0)  = n316 | ~n325;
  assign n327 = \V116(7)  & ~n227;
  assign n328 = ~n220 & n327;
  assign n329 = ~n219 & n328;
  assign n330 = ~\V133(10)  & n329;
  assign n331 = \V133(9)  & n330;
  assign n332 = ~\V133(10)  & n331;
  assign n333 = \V84(24)  & ~n220;
  assign n334 = ~n219 & n333;
  assign n335 = \V133(10)  & n334;
  assign n336 = \V84(24)  & n220;
  assign n337 = ~n219 & n336;
  assign n338 = \V84(24)  & n219;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~n335 & n339;
  assign n341 = ~n236 & n340;
  assign \V212(7)  = n332 | ~n341;
  assign n343 = \V116(6)  & ~n227;
  assign n344 = ~n220 & n343;
  assign n345 = ~n219 & n344;
  assign n346 = ~\V133(10)  & n345;
  assign n347 = \V133(9)  & n346;
  assign n348 = ~\V133(10)  & n347;
  assign n349 = \V84(23)  & ~n220;
  assign n350 = ~n219 & n349;
  assign n351 = \V133(10)  & n350;
  assign n352 = \V84(23)  & n220;
  assign n353 = ~n219 & n352;
  assign n354 = \V84(23)  & n219;
  assign n355 = ~n353 & ~n354;
  assign n356 = ~n351 & n355;
  assign n357 = ~n236 & n356;
  assign \V212(6)  = n348 | ~n357;
  assign n359 = \V116(9)  & ~n227;
  assign n360 = ~n220 & n359;
  assign n361 = ~n219 & n360;
  assign n362 = ~\V133(10)  & n361;
  assign n363 = \V133(9)  & n362;
  assign n364 = ~\V133(10)  & n363;
  assign n365 = \V84(26)  & ~n220;
  assign n366 = ~n219 & n365;
  assign n367 = \V133(10)  & n366;
  assign n368 = \V84(26)  & n220;
  assign n369 = ~n219 & n368;
  assign n370 = \V84(26)  & n219;
  assign n371 = ~n369 & ~n370;
  assign n372 = ~n367 & n371;
  assign n373 = ~n236 & n372;
  assign \V212(9)  = n364 | ~n373;
  assign n375 = \V116(8)  & ~n227;
  assign n376 = ~n220 & n375;
  assign n377 = ~n219 & n376;
  assign n378 = ~\V133(10)  & n377;
  assign n379 = \V133(9)  & n378;
  assign n380 = ~\V133(10)  & n379;
  assign n381 = \V84(25)  & ~n220;
  assign n382 = ~n219 & n381;
  assign n383 = \V133(10)  & n382;
  assign n384 = \V84(25)  & n220;
  assign n385 = ~n219 & n384;
  assign n386 = \V84(25)  & n219;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~n383 & n387;
  assign n389 = ~n236 & n388;
  assign \V212(8)  = n380 | ~n389;
  assign n391 = ~\V133(9)  & ~\V133(10) ;
  assign n392 = \V133(7)  & n391;
  assign n393 = \V133(1)  & ~\V133(10) ;
  assign n394 = \V133(2)  & n393;
  assign n395 = ~\V133(9)  & n394;
  assign n396 = \V122(0)  & ~n395;
  assign n397 = ~n392 & n396;
  assign n398 = \V133(10)  & n397;
  assign n399 = ~n392 & n395;
  assign n400 = \V121(17)  & n392;
  assign n401 = ~n399 & ~n400;
  assign \V214(0)  = n398 | ~n401;
  assign n403 = \V133(7)  & ~\V133(9) ;
  assign n404 = ~\V133(4)  & ~\V133(9) ;
  assign n405 = \V116(9)  & ~\V133(10) ;
  assign n406 = ~n404 & n405;
  assign n407 = ~n403 & n406;
  assign n408 = \V133(9)  & n407;
  assign n409 = ~\V133(10)  & n408;
  assign n410 = ~\V133(5)  & ~\V133(10) ;
  assign n411 = ~\V133(1)  & n410;
  assign n412 = \V133(0)  & n411;
  assign n413 = \V133(2)  & n412;
  assign n414 = ~\V133(6)  & n413;
  assign n415 = ~\V133(10)  & \V133(2) ;
  assign n416 = \V133(1)  & n415;
  assign n417 = ~\V133(3)  & n416;
  assign n418 = ~\V133(1)  & n415;
  assign n419 = \V133(8)  & n418;
  assign n420 = ~n417 & ~n419;
  assign n421 = ~n414 & n420;
  assign n422 = \V133(1)  & \V133(3) ;
  assign n423 = \V133(2)  & n422;
  assign n424 = ~\V133(10)  & ~n423;
  assign n425 = ~\V133(0)  & ~\V133(10) ;
  assign n426 = \V133(7)  & n425;
  assign n427 = ~\V133(5)  & n425;
  assign n428 = \V133(1)  & n410;
  assign n429 = ~\V133(2)  & n428;
  assign n430 = ~\V133(6)  & n429;
  assign n431 = \V133(8)  & n393;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~n427 & n432;
  assign n434 = ~n426 & n433;
  assign n435 = ~\V133(2)  & n411;
  assign n436 = ~\V133(6)  & n435;
  assign n437 = ~\V133(10)  & ~\V133(2) ;
  assign n438 = ~\V133(1)  & n437;
  assign n439 = \V133(7)  & n438;
  assign n440 = ~n436 & ~n439;
  assign n441 = n434 & n440;
  assign n442 = n424 & n441;
  assign n443 = n421 & n442;
  assign n444 = \V15(8)  & n421;
  assign n445 = n424 & n444;
  assign n446 = n434 & n445;
  assign n447 = ~n440 & n446;
  assign n448 = \V84(9)  & n434;
  assign n449 = n424 & n448;
  assign n450 = ~n421 & n449;
  assign n451 = \V47(1)  & ~n434;
  assign n452 = n424 & n451;
  assign n453 = \V47(9)  & ~n424;
  assign n454 = ~n452 & ~n453;
  assign n455 = ~n450 & n454;
  assign n456 = ~n447 & n455;
  assign n457 = ~n443 & n456;
  assign n458 = ~n403 & ~n457;
  assign n459 = ~n404 & n458;
  assign n460 = \V133(10)  & n459;
  assign n461 = n403 & ~n457;
  assign n462 = ~n404 & n461;
  assign n463 = n404 & ~n457;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~n460 & n464;
  assign \V143(0)  = n409 | ~n465;
  assign n467 = ~\V133(6)  & ~\V133(9) ;
  assign n468 = ~\V133(4)  & n467;
  assign n469 = ~\V133(10)  & \V116(11) ;
  assign n470 = ~n468 & n469;
  assign n471 = ~n403 & n470;
  assign n472 = \V133(9)  & n471;
  assign n473 = ~\V133(10)  & n472;
  assign n474 = \V15(10)  & n421;
  assign n475 = n424 & n474;
  assign n476 = n434 & n475;
  assign n477 = ~n440 & n476;
  assign n478 = \V84(11)  & n434;
  assign n479 = n424 & n478;
  assign n480 = ~n421 & n479;
  assign n481 = \V47(3)  & ~n434;
  assign n482 = n424 & n481;
  assign n483 = \V47(11)  & ~n424;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n480 & n484;
  assign n486 = ~n477 & n485;
  assign n487 = ~n443 & n486;
  assign n488 = ~n403 & ~n487;
  assign n489 = ~n468 & n488;
  assign n490 = \V133(10)  & n489;
  assign n491 = n403 & ~n487;
  assign n492 = ~n468 & n491;
  assign n493 = n468 & ~n487;
  assign n494 = ~n492 & ~n493;
  assign n495 = ~n490 & n494;
  assign \V145(1)  = n473 | ~n495;
  assign n497 = ~\V133(10)  & \V116(10) ;
  assign n498 = ~n468 & n497;
  assign n499 = ~n403 & n498;
  assign n500 = \V133(9)  & n499;
  assign n501 = ~\V133(10)  & n500;
  assign n502 = \V15(9)  & n421;
  assign n503 = n424 & n502;
  assign n504 = n434 & n503;
  assign n505 = ~n440 & n504;
  assign n506 = \V84(10)  & n434;
  assign n507 = n424 & n506;
  assign n508 = ~n421 & n507;
  assign n509 = \V47(2)  & ~n434;
  assign n510 = n424 & n509;
  assign n511 = \V47(10)  & ~n424;
  assign n512 = ~n510 & ~n511;
  assign n513 = ~n508 & n512;
  assign n514 = ~n505 & n513;
  assign n515 = ~n443 & n514;
  assign n516 = ~n403 & ~n515;
  assign n517 = ~n468 & n516;
  assign n518 = \V133(10)  & n517;
  assign n519 = n403 & ~n515;
  assign n520 = ~n468 & n519;
  assign n521 = n468 & ~n515;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~n518 & n522;
  assign \V145(0)  = n501 | ~n523;
  assign n525 = \V133(3)  & n404;
  assign n526 = ~\V133(6)  & n215;
  assign n527 = ~\V133(4)  & n526;
  assign n528 = ~\V133(2)  & n467;
  assign n529 = ~\V133(4)  & n528;
  assign n530 = \V133(9)  & ~\V133(10) ;
  assign n531 = \V84(15)  & ~n530;
  assign n532 = ~n403 & n531;
  assign n533 = ~n529 & n532;
  assign n534 = ~n527 & n533;
  assign n535 = ~n525 & n534;
  assign n536 = ~\V133(10)  & n535;
  assign n537 = ~\V133(7)  & n536;
  assign n538 = ~\V133(9)  & n537;
  assign n539 = ~\V133(4)  & n538;
  assign n540 = ~\V133(3)  & n539;
  assign n541 = \V133(2)  & n540;
  assign n542 = \V133(1)  & n541;
  assign n543 = ~\V133(10)  & n542;
  assign n544 = \V116(15)  & ~\V133(10) ;
  assign n545 = ~n525 & n544;
  assign n546 = ~n527 & n545;
  assign n547 = ~n529 & n546;
  assign n548 = ~n403 & n547;
  assign n549 = n530 & n548;
  assign n550 = \V15(14)  & n421;
  assign n551 = n424 & n550;
  assign n552 = n434 & n551;
  assign n553 = ~n440 & n552;
  assign n554 = \V47(4)  & n434;
  assign n555 = n424 & n554;
  assign n556 = ~n421 & n555;
  assign n557 = \V47(7)  & ~n434;
  assign n558 = n424 & n557;
  assign n559 = \V47(15)  & ~n424;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n556 & n560;
  assign n562 = ~n553 & n561;
  assign n563 = ~n443 & n562;
  assign n564 = ~n403 & ~n563;
  assign n565 = ~n529 & n564;
  assign n566 = ~n527 & n565;
  assign n567 = ~n525 & n566;
  assign n568 = \V133(10)  & n567;
  assign n569 = ~n525 & ~n563;
  assign n570 = ~n527 & n569;
  assign n571 = ~n529 & n570;
  assign n572 = n403 & n571;
  assign n573 = ~n529 & ~n563;
  assign n574 = ~n527 & n573;
  assign n575 = n525 & n574;
  assign n576 = n529 & ~n563;
  assign n577 = ~n527 & n576;
  assign n578 = n527 & ~n563;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n575 & n579;
  assign n581 = ~n572 & n580;
  assign n582 = ~n568 & n581;
  assign n583 = ~n549 & n582;
  assign \V149(2)  = n543 | ~n583;
  assign n585 = \V84(14)  & ~n530;
  assign n586 = ~n403 & n585;
  assign n587 = ~n529 & n586;
  assign n588 = ~n527 & n587;
  assign n589 = ~n525 & n588;
  assign n590 = ~\V133(10)  & n589;
  assign n591 = ~\V133(7)  & n590;
  assign n592 = ~\V133(9)  & n591;
  assign n593 = ~\V133(4)  & n592;
  assign n594 = ~\V133(3)  & n593;
  assign n595 = \V133(2)  & n594;
  assign n596 = \V133(1)  & n595;
  assign n597 = ~\V133(10)  & n596;
  assign n598 = \V116(14)  & ~\V133(10) ;
  assign n599 = ~n525 & n598;
  assign n600 = ~n527 & n599;
  assign n601 = ~n529 & n600;
  assign n602 = ~n403 & n601;
  assign n603 = n530 & n602;
  assign n604 = \V15(13)  & n421;
  assign n605 = n424 & n604;
  assign n606 = n434 & n605;
  assign n607 = ~n440 & n606;
  assign n608 = \V47(3)  & n434;
  assign n609 = n424 & n608;
  assign n610 = ~n421 & n609;
  assign n611 = \V47(6)  & ~n434;
  assign n612 = n424 & n611;
  assign n613 = \V47(14)  & ~n424;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n610 & n614;
  assign n616 = ~n607 & n615;
  assign n617 = ~n443 & n616;
  assign n618 = ~n403 & ~n617;
  assign n619 = ~n529 & n618;
  assign n620 = ~n527 & n619;
  assign n621 = ~n525 & n620;
  assign n622 = \V133(10)  & n621;
  assign n623 = ~n525 & ~n617;
  assign n624 = ~n527 & n623;
  assign n625 = ~n529 & n624;
  assign n626 = n403 & n625;
  assign n627 = ~n529 & ~n617;
  assign n628 = ~n527 & n627;
  assign n629 = n525 & n628;
  assign n630 = n529 & ~n617;
  assign n631 = ~n527 & n630;
  assign n632 = n527 & ~n617;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~n629 & n633;
  assign n635 = ~n626 & n634;
  assign n636 = ~n622 & n635;
  assign n637 = ~n603 & n636;
  assign \V149(1)  = n597 | ~n637;
  assign n639 = \V84(13)  & ~n530;
  assign n640 = ~n403 & n639;
  assign n641 = ~n529 & n640;
  assign n642 = ~n527 & n641;
  assign n643 = ~n525 & n642;
  assign n644 = ~\V133(10)  & n643;
  assign n645 = ~\V133(7)  & n644;
  assign n646 = ~\V133(9)  & n645;
  assign n647 = ~\V133(4)  & n646;
  assign n648 = ~\V133(3)  & n647;
  assign n649 = \V133(2)  & n648;
  assign n650 = \V133(1)  & n649;
  assign n651 = ~\V133(10)  & n650;
  assign n652 = ~\V133(10)  & \V116(13) ;
  assign n653 = ~n525 & n652;
  assign n654 = ~n527 & n653;
  assign n655 = ~n529 & n654;
  assign n656 = ~n403 & n655;
  assign n657 = n530 & n656;
  assign n658 = \V15(12)  & n421;
  assign n659 = n424 & n658;
  assign n660 = n434 & n659;
  assign n661 = ~n440 & n660;
  assign n662 = \V47(2)  & n434;
  assign n663 = n424 & n662;
  assign n664 = ~n421 & n663;
  assign n665 = \V47(5)  & ~n434;
  assign n666 = n424 & n665;
  assign n667 = \V47(13)  & ~n424;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n664 & n668;
  assign n670 = ~n661 & n669;
  assign n671 = ~n443 & n670;
  assign n672 = ~n403 & ~n671;
  assign n673 = ~n529 & n672;
  assign n674 = ~n527 & n673;
  assign n675 = ~n525 & n674;
  assign n676 = \V133(10)  & n675;
  assign n677 = ~n525 & ~n671;
  assign n678 = ~n527 & n677;
  assign n679 = ~n529 & n678;
  assign n680 = n403 & n679;
  assign n681 = ~n529 & ~n671;
  assign n682 = ~n527 & n681;
  assign n683 = n525 & n682;
  assign n684 = n529 & ~n671;
  assign n685 = ~n527 & n684;
  assign n686 = n527 & ~n671;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n683 & n687;
  assign n689 = ~n680 & n688;
  assign n690 = ~n676 & n689;
  assign n691 = ~n657 & n690;
  assign \V149(0)  = n651 | ~n691;
  assign n693 = ~\V133(2)  & n391;
  assign n694 = \V133(7)  & n693;
  assign n695 = ~\V133(1)  & ~\V133(10) ;
  assign n696 = ~\V133(9)  & n695;
  assign n697 = \V133(7)  & n696;
  assign n698 = ~\V133(7)  & n391;
  assign n699 = ~\V133(10)  & ~n698;
  assign n700 = ~n697 & n699;
  assign n701 = ~n694 & n700;
  assign n702 = ~n530 & n701;
  assign n703 = \V84(0)  & ~n530;
  assign n704 = ~n694 & n703;
  assign n705 = ~n697 & n704;
  assign n706 = ~n698 & n705;
  assign n707 = \V133(10)  & n706;
  assign n708 = \V116(0)  & ~n698;
  assign n709 = ~n697 & n708;
  assign n710 = ~n694 & n709;
  assign n711 = n530 & n710;
  assign n712 = \V49(0)  & ~n694;
  assign n713 = ~n697 & n712;
  assign n714 = n698 & n713;
  assign n715 = \V48(0)  & n694;
  assign n716 = ~n697 & n715;
  assign n717 = \V48(0)  & n697;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n714 & n718;
  assign n720 = ~n711 & n719;
  assign n721 = ~n707 & n720;
  assign \V134(0)  = n702 | ~n721;
  assign n723 = ~\V133(7)  & n693;
  assign n724 = \V133(8)  & n391;
  assign n725 = ~\V133(9)  & ~\V133(8) ;
  assign n726 = \V133(7)  & n725;
  assign n727 = \V133(1)  & ~\V133(9) ;
  assign n728 = \V133(2)  & n727;
  assign n729 = ~\V133(8)  & n728;
  assign n730 = ~\V133(4)  & n729;
  assign n731 = ~\V133(7)  & n696;
  assign n732 = \V52(0)  & ~n731;
  assign n733 = ~\V133(10)  & n732;
  assign n734 = ~n730 & n733;
  assign n735 = ~n726 & n734;
  assign n736 = ~n724 & n735;
  assign n737 = n723 & n736;
  assign n738 = \V52(0)  & ~n724;
  assign n739 = ~n726 & n738;
  assign n740 = ~n730 & n739;
  assign n741 = ~\V133(10)  & n740;
  assign n742 = n731 & n741;
  assign n743 = \V116(2)  & ~n723;
  assign n744 = ~n724 & n743;
  assign n745 = ~n726 & n744;
  assign n746 = ~n730 & n745;
  assign n747 = ~\V133(10)  & n746;
  assign n748 = ~n731 & n747;
  assign n749 = \V133(9)  & n748;
  assign n750 = ~\V133(10)  & n749;
  assign n751 = \V15(1)  & n421;
  assign n752 = n424 & n751;
  assign n753 = n434 & n752;
  assign n754 = ~n440 & n753;
  assign n755 = \V84(2)  & n434;
  assign n756 = n424 & n755;
  assign n757 = ~n421 & n756;
  assign n758 = \V47(2)  & ~n424;
  assign n759 = ~n443 & ~n758;
  assign n760 = ~n757 & n759;
  assign n761 = ~n754 & n760;
  assign n762 = ~n726 & ~n761;
  assign n763 = ~n730 & n762;
  assign n764 = \V133(10)  & n763;
  assign n765 = n726 & ~n761;
  assign n766 = ~n730 & n765;
  assign n767 = n730 & ~n761;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n764 & n768;
  assign n770 = ~n750 & n769;
  assign n771 = ~n742 & n770;
  assign \V136(1)  = n737 | ~n771;
  assign n773 = \V116(1)  & ~n723;
  assign n774 = ~n724 & n773;
  assign n775 = ~n726 & n774;
  assign n776 = ~n730 & n775;
  assign n777 = ~\V133(10)  & n776;
  assign n778 = ~n731 & n777;
  assign n779 = \V133(9)  & n778;
  assign n780 = ~\V133(10)  & n779;
  assign n781 = \V51(0)  & ~n731;
  assign n782 = ~\V133(10)  & n781;
  assign n783 = ~n730 & n782;
  assign n784 = ~n726 & n783;
  assign n785 = ~n724 & n784;
  assign n786 = n723 & n785;
  assign n787 = \V51(0)  & ~n724;
  assign n788 = ~n726 & n787;
  assign n789 = ~n730 & n788;
  assign n790 = ~\V133(10)  & n789;
  assign n791 = n731 & n790;
  assign n792 = \V50(0)  & ~\V133(10) ;
  assign n793 = ~n730 & n792;
  assign n794 = ~n726 & n793;
  assign n795 = n724 & n794;
  assign n796 = \V15(0)  & n421;
  assign n797 = n424 & n796;
  assign n798 = n434 & n797;
  assign n799 = ~n440 & n798;
  assign n800 = \V84(1)  & n434;
  assign n801 = n424 & n800;
  assign n802 = ~n421 & n801;
  assign n803 = \V47(1)  & ~n424;
  assign n804 = ~n443 & ~n803;
  assign n805 = ~n802 & n804;
  assign n806 = ~n799 & n805;
  assign n807 = ~n726 & ~n806;
  assign n808 = ~n730 & n807;
  assign n809 = \V133(10)  & n808;
  assign n810 = n726 & ~n806;
  assign n811 = ~n730 & n810;
  assign n812 = n730 & ~n806;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n809 & n813;
  assign n815 = ~n795 & n814;
  assign n816 = ~n791 & n815;
  assign n817 = ~n786 & n816;
  assign \V136(0)  = n780 | ~n817;
  assign n819 = \V84(28)  & ~n530;
  assign n820 = ~n403 & n819;
  assign n821 = ~n529 & n820;
  assign n822 = ~n527 & n821;
  assign n823 = ~n525 & n822;
  assign n824 = ~\V133(10)  & n823;
  assign n825 = ~\V133(7)  & n824;
  assign n826 = ~\V133(9)  & n825;
  assign n827 = ~\V133(4)  & n826;
  assign n828 = ~\V133(3)  & n827;
  assign n829 = \V133(2)  & n828;
  assign n830 = \V133(1)  & n829;
  assign n831 = ~\V133(10)  & n830;
  assign n832 = ~\V133(10)  & \V116(28) ;
  assign n833 = ~n525 & n832;
  assign n834 = ~n527 & n833;
  assign n835 = ~n529 & n834;
  assign n836 = ~n403 & n835;
  assign n837 = n530 & n836;
  assign n838 = \V47(13)  & n421;
  assign n839 = n424 & n838;
  assign n840 = n434 & n839;
  assign n841 = ~n440 & n840;
  assign n842 = \V47(17)  & n434;
  assign n843 = n424 & n842;
  assign n844 = ~n421 & n843;
  assign n845 = \V47(20)  & ~n434;
  assign n846 = n424 & n845;
  assign n847 = \V47(28)  & ~n424;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n844 & n848;
  assign n850 = ~n841 & n849;
  assign n851 = ~n443 & n850;
  assign n852 = ~n403 & ~n851;
  assign n853 = ~n529 & n852;
  assign n854 = ~n527 & n853;
  assign n855 = ~n525 & n854;
  assign n856 = \V133(10)  & n855;
  assign n857 = ~n525 & ~n851;
  assign n858 = ~n527 & n857;
  assign n859 = ~n529 & n858;
  assign n860 = n403 & n859;
  assign n861 = ~n529 & ~n851;
  assign n862 = ~n527 & n861;
  assign n863 = n525 & n862;
  assign n864 = n529 & ~n851;
  assign n865 = ~n527 & n864;
  assign n866 = n527 & ~n851;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n863 & n867;
  assign n869 = ~n860 & n868;
  assign n870 = ~n856 & n869;
  assign n871 = ~n837 & n870;
  assign \V165(11)  = n831 | ~n871;
  assign n873 = \V133(7)  & n215;
  assign n874 = ~\V133(1)  & ~\V133(0) ;
  assign n875 = ~\V133(9)  & n874;
  assign n876 = \V133(5)  & n875;
  assign n877 = ~\V133(5)  & n526;
  assign n878 = ~\V133(4)  & n877;
  assign n879 = ~\V133(1)  & \V133(0) ;
  assign n880 = ~\V118(0)  & n879;
  assign n881 = ~\V133(9)  & n880;
  assign n882 = \V133(5)  & n881;
  assign n883 = \V133(3)  & n728;
  assign n884 = ~\V133(4)  & n883;
  assign n885 = ~\V133(6)  & n884;
  assign n886 = \V116(3)  & ~\V133(10) ;
  assign n887 = ~n885 & n886;
  assign n888 = ~n882 & n887;
  assign n889 = ~n878 & n888;
  assign n890 = ~n876 & n889;
  assign n891 = ~n873 & n890;
  assign n892 = \V133(9)  & n891;
  assign n893 = ~\V133(10)  & n892;
  assign n894 = \V47(20)  & n421;
  assign n895 = n424 & n894;
  assign n896 = n434 & n895;
  assign n897 = ~n440 & n896;
  assign n898 = \V47(24)  & n434;
  assign n899 = n424 & n898;
  assign n900 = ~n421 & n899;
  assign n901 = \V47(27)  & ~n434;
  assign n902 = n424 & n901;
  assign n903 = \V84(3)  & ~n424;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n900 & n904;
  assign n906 = ~n897 & n905;
  assign n907 = ~n443 & n906;
  assign n908 = ~n873 & ~n907;
  assign n909 = ~n876 & n908;
  assign n910 = ~n878 & n909;
  assign n911 = ~n882 & n910;
  assign n912 = ~n885 & n911;
  assign n913 = \V133(10)  & n912;
  assign n914 = ~n885 & ~n907;
  assign n915 = ~n882 & n914;
  assign n916 = ~n878 & n915;
  assign n917 = ~n876 & n916;
  assign n918 = n873 & n917;
  assign n919 = ~n876 & ~n907;
  assign n920 = ~n878 & n919;
  assign n921 = ~n882 & n920;
  assign n922 = n885 & n921;
  assign n923 = ~n882 & ~n907;
  assign n924 = ~n878 & n923;
  assign n925 = n876 & n924;
  assign n926 = n882 & ~n907;
  assign n927 = ~n878 & n926;
  assign n928 = n878 & ~n907;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n925 & n929;
  assign n931 = ~n922 & n930;
  assign n932 = ~n918 & n931;
  assign n933 = ~n913 & n932;
  assign \V197(3)  = n893 | ~n933;
  assign n935 = \V84(27)  & ~n530;
  assign n936 = ~n403 & n935;
  assign n937 = ~n529 & n936;
  assign n938 = ~n527 & n937;
  assign n939 = ~n525 & n938;
  assign n940 = ~\V133(10)  & n939;
  assign n941 = ~\V133(7)  & n940;
  assign n942 = ~\V133(9)  & n941;
  assign n943 = ~\V133(4)  & n942;
  assign n944 = ~\V133(3)  & n943;
  assign n945 = \V133(2)  & n944;
  assign n946 = \V133(1)  & n945;
  assign n947 = ~\V133(10)  & n946;
  assign n948 = ~\V133(10)  & \V116(27) ;
  assign n949 = ~n525 & n948;
  assign n950 = ~n527 & n949;
  assign n951 = ~n529 & n950;
  assign n952 = ~n403 & n951;
  assign n953 = n530 & n952;
  assign n954 = \V47(12)  & n421;
  assign n955 = n424 & n954;
  assign n956 = n434 & n955;
  assign n957 = ~n440 & n956;
  assign n958 = \V47(16)  & n434;
  assign n959 = n424 & n958;
  assign n960 = ~n421 & n959;
  assign n961 = \V47(19)  & ~n434;
  assign n962 = n424 & n961;
  assign n963 = \V47(27)  & ~n424;
  assign n964 = ~n962 & ~n963;
  assign n965 = ~n960 & n964;
  assign n966 = ~n957 & n965;
  assign n967 = ~n443 & n966;
  assign n968 = ~n403 & ~n967;
  assign n969 = ~n529 & n968;
  assign n970 = ~n527 & n969;
  assign n971 = ~n525 & n970;
  assign n972 = \V133(10)  & n971;
  assign n973 = ~n525 & ~n967;
  assign n974 = ~n527 & n973;
  assign n975 = ~n529 & n974;
  assign n976 = n403 & n975;
  assign n977 = ~n529 & ~n967;
  assign n978 = ~n527 & n977;
  assign n979 = n525 & n978;
  assign n980 = n529 & ~n967;
  assign n981 = ~n527 & n980;
  assign n982 = n527 & ~n967;
  assign n983 = ~n981 & ~n982;
  assign n984 = ~n979 & n983;
  assign n985 = ~n976 & n984;
  assign n986 = ~n972 & n985;
  assign n987 = ~n953 & n986;
  assign \V165(10)  = n947 | ~n987;
  assign n989 = \V116(2)  & ~\V133(10) ;
  assign n990 = ~n885 & n989;
  assign n991 = ~n882 & n990;
  assign n992 = ~n878 & n991;
  assign n993 = ~n876 & n992;
  assign n994 = ~n873 & n993;
  assign n995 = \V133(9)  & n994;
  assign n996 = ~\V133(10)  & n995;
  assign n997 = \V47(19)  & n421;
  assign n998 = n424 & n997;
  assign n999 = n434 & n998;
  assign n1000 = ~n440 & n999;
  assign n1001 = \V47(23)  & n434;
  assign n1002 = n424 & n1001;
  assign n1003 = ~n421 & n1002;
  assign n1004 = \V47(26)  & ~n434;
  assign n1005 = n424 & n1004;
  assign n1006 = \V84(2)  & ~n424;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1003 & n1007;
  assign n1009 = ~n1000 & n1008;
  assign n1010 = ~n443 & n1009;
  assign n1011 = ~n873 & ~n1010;
  assign n1012 = ~n876 & n1011;
  assign n1013 = ~n878 & n1012;
  assign n1014 = ~n882 & n1013;
  assign n1015 = ~n885 & n1014;
  assign n1016 = \V133(10)  & n1015;
  assign n1017 = ~n885 & ~n1010;
  assign n1018 = ~n882 & n1017;
  assign n1019 = ~n878 & n1018;
  assign n1020 = ~n876 & n1019;
  assign n1021 = n873 & n1020;
  assign n1022 = ~n876 & ~n1010;
  assign n1023 = ~n878 & n1022;
  assign n1024 = ~n882 & n1023;
  assign n1025 = n885 & n1024;
  assign n1026 = ~n882 & ~n1010;
  assign n1027 = ~n878 & n1026;
  assign n1028 = n876 & n1027;
  assign n1029 = n882 & ~n1010;
  assign n1030 = ~n878 & n1029;
  assign n1031 = n878 & ~n1010;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = ~n1028 & n1032;
  assign n1034 = ~n1025 & n1033;
  assign n1035 = ~n1021 & n1034;
  assign n1036 = ~n1016 & n1035;
  assign \V197(2)  = n996 | ~n1036;
  assign n1038 = \V84(30)  & ~n530;
  assign n1039 = ~n403 & n1038;
  assign n1040 = ~n529 & n1039;
  assign n1041 = ~n527 & n1040;
  assign n1042 = ~n525 & n1041;
  assign n1043 = ~\V133(10)  & n1042;
  assign n1044 = ~\V133(7)  & n1043;
  assign n1045 = ~\V133(9)  & n1044;
  assign n1046 = ~\V133(4)  & n1045;
  assign n1047 = ~\V133(3)  & n1046;
  assign n1048 = \V133(2)  & n1047;
  assign n1049 = \V133(1)  & n1048;
  assign n1050 = ~\V133(10)  & n1049;
  assign n1051 = \V116(30)  & ~\V133(10) ;
  assign n1052 = ~n525 & n1051;
  assign n1053 = ~n527 & n1052;
  assign n1054 = ~n529 & n1053;
  assign n1055 = ~n403 & n1054;
  assign n1056 = n530 & n1055;
  assign n1057 = \V47(15)  & n421;
  assign n1058 = n424 & n1057;
  assign n1059 = n434 & n1058;
  assign n1060 = ~n440 & n1059;
  assign n1061 = \V47(19)  & n434;
  assign n1062 = n424 & n1061;
  assign n1063 = ~n421 & n1062;
  assign n1064 = \V47(22)  & ~n434;
  assign n1065 = n424 & n1064;
  assign n1066 = \V47(30)  & ~n424;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~n1063 & n1067;
  assign n1069 = ~n1060 & n1068;
  assign n1070 = ~n443 & n1069;
  assign n1071 = ~n403 & ~n1070;
  assign n1072 = ~n529 & n1071;
  assign n1073 = ~n527 & n1072;
  assign n1074 = ~n525 & n1073;
  assign n1075 = \V133(10)  & n1074;
  assign n1076 = ~n525 & ~n1070;
  assign n1077 = ~n527 & n1076;
  assign n1078 = ~n529 & n1077;
  assign n1079 = n403 & n1078;
  assign n1080 = ~n529 & ~n1070;
  assign n1081 = ~n527 & n1080;
  assign n1082 = n525 & n1081;
  assign n1083 = n529 & ~n1070;
  assign n1084 = ~n527 & n1083;
  assign n1085 = n527 & ~n1070;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1082 & n1086;
  assign n1088 = ~n1079 & n1087;
  assign n1089 = ~n1075 & n1088;
  assign n1090 = ~n1056 & n1089;
  assign \V165(13)  = n1050 | ~n1090;
  assign n1092 = \V116(5)  & ~\V133(10) ;
  assign n1093 = ~n885 & n1092;
  assign n1094 = ~n882 & n1093;
  assign n1095 = ~n878 & n1094;
  assign n1096 = ~n876 & n1095;
  assign n1097 = ~n873 & n1096;
  assign n1098 = \V133(9)  & n1097;
  assign n1099 = ~\V133(10)  & n1098;
  assign n1100 = \V47(22)  & n421;
  assign n1101 = n424 & n1100;
  assign n1102 = n434 & n1101;
  assign n1103 = ~n440 & n1102;
  assign n1104 = \V47(26)  & n434;
  assign n1105 = n424 & n1104;
  assign n1106 = ~n421 & n1105;
  assign n1107 = \V47(29)  & ~n434;
  assign n1108 = n424 & n1107;
  assign n1109 = \V84(5)  & ~n424;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1106 & n1110;
  assign n1112 = ~n1103 & n1111;
  assign n1113 = ~n443 & n1112;
  assign n1114 = ~n873 & ~n1113;
  assign n1115 = ~n876 & n1114;
  assign n1116 = ~n878 & n1115;
  assign n1117 = ~n882 & n1116;
  assign n1118 = ~n885 & n1117;
  assign n1119 = \V133(10)  & n1118;
  assign n1120 = ~n885 & ~n1113;
  assign n1121 = ~n882 & n1120;
  assign n1122 = ~n878 & n1121;
  assign n1123 = ~n876 & n1122;
  assign n1124 = n873 & n1123;
  assign n1125 = ~n876 & ~n1113;
  assign n1126 = ~n878 & n1125;
  assign n1127 = ~n882 & n1126;
  assign n1128 = n885 & n1127;
  assign n1129 = ~n882 & ~n1113;
  assign n1130 = ~n878 & n1129;
  assign n1131 = n876 & n1130;
  assign n1132 = n882 & ~n1113;
  assign n1133 = ~n878 & n1132;
  assign n1134 = n878 & ~n1113;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = ~n1131 & n1135;
  assign n1137 = ~n1128 & n1136;
  assign n1138 = ~n1124 & n1137;
  assign n1139 = ~n1119 & n1138;
  assign \V197(5)  = n1099 | ~n1139;
  assign n1141 = \V84(29)  & ~n530;
  assign n1142 = ~n403 & n1141;
  assign n1143 = ~n529 & n1142;
  assign n1144 = ~n527 & n1143;
  assign n1145 = ~n525 & n1144;
  assign n1146 = ~\V133(10)  & n1145;
  assign n1147 = ~\V133(7)  & n1146;
  assign n1148 = ~\V133(9)  & n1147;
  assign n1149 = ~\V133(4)  & n1148;
  assign n1150 = ~\V133(3)  & n1149;
  assign n1151 = \V133(2)  & n1150;
  assign n1152 = \V133(1)  & n1151;
  assign n1153 = ~\V133(10)  & n1152;
  assign n1154 = ~\V133(10)  & \V116(29) ;
  assign n1155 = ~n525 & n1154;
  assign n1156 = ~n527 & n1155;
  assign n1157 = ~n529 & n1156;
  assign n1158 = ~n403 & n1157;
  assign n1159 = n530 & n1158;
  assign n1160 = \V47(14)  & n421;
  assign n1161 = n424 & n1160;
  assign n1162 = n434 & n1161;
  assign n1163 = ~n440 & n1162;
  assign n1164 = \V47(18)  & n434;
  assign n1165 = n424 & n1164;
  assign n1166 = ~n421 & n1165;
  assign n1167 = \V47(21)  & ~n434;
  assign n1168 = n424 & n1167;
  assign n1169 = \V47(29)  & ~n424;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1166 & n1170;
  assign n1172 = ~n1163 & n1171;
  assign n1173 = ~n443 & n1172;
  assign n1174 = ~n403 & ~n1173;
  assign n1175 = ~n529 & n1174;
  assign n1176 = ~n527 & n1175;
  assign n1177 = ~n525 & n1176;
  assign n1178 = \V133(10)  & n1177;
  assign n1179 = ~n525 & ~n1173;
  assign n1180 = ~n527 & n1179;
  assign n1181 = ~n529 & n1180;
  assign n1182 = n403 & n1181;
  assign n1183 = ~n529 & ~n1173;
  assign n1184 = ~n527 & n1183;
  assign n1185 = n525 & n1184;
  assign n1186 = n529 & ~n1173;
  assign n1187 = ~n527 & n1186;
  assign n1188 = n527 & ~n1173;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1185 & n1189;
  assign n1191 = ~n1182 & n1190;
  assign n1192 = ~n1178 & n1191;
  assign n1193 = ~n1159 & n1192;
  assign \V165(12)  = n1153 | ~n1193;
  assign n1195 = \V116(4)  & ~\V133(10) ;
  assign n1196 = ~n885 & n1195;
  assign n1197 = ~n882 & n1196;
  assign n1198 = ~n878 & n1197;
  assign n1199 = ~n876 & n1198;
  assign n1200 = ~n873 & n1199;
  assign n1201 = \V133(9)  & n1200;
  assign n1202 = ~\V133(10)  & n1201;
  assign n1203 = \V47(21)  & n421;
  assign n1204 = n424 & n1203;
  assign n1205 = n434 & n1204;
  assign n1206 = ~n440 & n1205;
  assign n1207 = \V47(25)  & n434;
  assign n1208 = n424 & n1207;
  assign n1209 = ~n421 & n1208;
  assign n1210 = \V47(28)  & ~n434;
  assign n1211 = n424 & n1210;
  assign n1212 = \V84(4)  & ~n424;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = ~n1209 & n1213;
  assign n1215 = ~n1206 & n1214;
  assign n1216 = ~n443 & n1215;
  assign n1217 = ~n873 & ~n1216;
  assign n1218 = ~n876 & n1217;
  assign n1219 = ~n878 & n1218;
  assign n1220 = ~n882 & n1219;
  assign n1221 = ~n885 & n1220;
  assign n1222 = \V133(10)  & n1221;
  assign n1223 = ~n885 & ~n1216;
  assign n1224 = ~n882 & n1223;
  assign n1225 = ~n878 & n1224;
  assign n1226 = ~n876 & n1225;
  assign n1227 = n873 & n1226;
  assign n1228 = ~n876 & ~n1216;
  assign n1229 = ~n878 & n1228;
  assign n1230 = ~n882 & n1229;
  assign n1231 = n885 & n1230;
  assign n1232 = ~n882 & ~n1216;
  assign n1233 = ~n878 & n1232;
  assign n1234 = n876 & n1233;
  assign n1235 = n882 & ~n1216;
  assign n1236 = ~n878 & n1235;
  assign n1237 = n878 & ~n1216;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1234 & n1238;
  assign n1240 = ~n1231 & n1239;
  assign n1241 = ~n1227 & n1240;
  assign n1242 = ~n1222 & n1241;
  assign \V197(4)  = n1202 | ~n1242;
  assign n1244 = ~n885 & n948;
  assign n1245 = ~n882 & n1244;
  assign n1246 = ~n878 & n1245;
  assign n1247 = ~n876 & n1246;
  assign n1248 = ~n873 & n1247;
  assign n1249 = \V133(9)  & n1248;
  assign n1250 = ~\V133(10)  & n1249;
  assign n1251 = \V84(12)  & n421;
  assign n1252 = n424 & n1251;
  assign n1253 = n434 & n1252;
  assign n1254 = ~n440 & n1253;
  assign n1255 = \V84(16)  & n434;
  assign n1256 = n424 & n1255;
  assign n1257 = ~n421 & n1256;
  assign n1258 = \V84(19)  & ~n434;
  assign n1259 = n424 & n1258;
  assign n1260 = \V84(27)  & ~n424;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1257 & n1261;
  assign n1263 = ~n1254 & n1262;
  assign n1264 = ~n443 & n1263;
  assign n1265 = ~n873 & ~n1264;
  assign n1266 = ~n876 & n1265;
  assign n1267 = ~n878 & n1266;
  assign n1268 = ~n882 & n1267;
  assign n1269 = ~n885 & n1268;
  assign n1270 = \V133(10)  & n1269;
  assign n1271 = ~n885 & ~n1264;
  assign n1272 = ~n882 & n1271;
  assign n1273 = ~n878 & n1272;
  assign n1274 = ~n876 & n1273;
  assign n1275 = n873 & n1274;
  assign n1276 = ~n876 & ~n1264;
  assign n1277 = ~n878 & n1276;
  assign n1278 = ~n882 & n1277;
  assign n1279 = n885 & n1278;
  assign n1280 = ~n882 & ~n1264;
  assign n1281 = ~n878 & n1280;
  assign n1282 = n876 & n1281;
  assign n1283 = n882 & ~n1264;
  assign n1284 = ~n878 & n1283;
  assign n1285 = n878 & ~n1264;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1282 & n1286;
  assign n1288 = ~n1279 & n1287;
  assign n1289 = ~n1275 & n1288;
  assign n1290 = ~n1270 & n1289;
  assign \V197(27)  = n1250 | ~n1290;
  assign n1292 = ~\V133(10)  & \V116(26) ;
  assign n1293 = ~n885 & n1292;
  assign n1294 = ~n882 & n1293;
  assign n1295 = ~n878 & n1294;
  assign n1296 = ~n876 & n1295;
  assign n1297 = ~n873 & n1296;
  assign n1298 = \V133(9)  & n1297;
  assign n1299 = ~\V133(10)  & n1298;
  assign n1300 = \V84(11)  & n421;
  assign n1301 = n424 & n1300;
  assign n1302 = n434 & n1301;
  assign n1303 = ~n440 & n1302;
  assign n1304 = \V84(15)  & n434;
  assign n1305 = n424 & n1304;
  assign n1306 = ~n421 & n1305;
  assign n1307 = \V84(18)  & ~n434;
  assign n1308 = n424 & n1307;
  assign n1309 = \V84(26)  & ~n424;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1306 & n1310;
  assign n1312 = ~n1303 & n1311;
  assign n1313 = ~n443 & n1312;
  assign n1314 = ~n873 & ~n1313;
  assign n1315 = ~n876 & n1314;
  assign n1316 = ~n878 & n1315;
  assign n1317 = ~n882 & n1316;
  assign n1318 = ~n885 & n1317;
  assign n1319 = \V133(10)  & n1318;
  assign n1320 = ~n885 & ~n1313;
  assign n1321 = ~n882 & n1320;
  assign n1322 = ~n878 & n1321;
  assign n1323 = ~n876 & n1322;
  assign n1324 = n873 & n1323;
  assign n1325 = ~n876 & ~n1313;
  assign n1326 = ~n878 & n1325;
  assign n1327 = ~n882 & n1326;
  assign n1328 = n885 & n1327;
  assign n1329 = ~n882 & ~n1313;
  assign n1330 = ~n878 & n1329;
  assign n1331 = n876 & n1330;
  assign n1332 = n882 & ~n1313;
  assign n1333 = ~n878 & n1332;
  assign n1334 = n878 & ~n1313;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1331 & n1335;
  assign n1337 = ~n1328 & n1336;
  assign n1338 = ~n1324 & n1337;
  assign n1339 = ~n1319 & n1338;
  assign \V197(26)  = n1299 | ~n1339;
  assign n1341 = \V84(31)  & ~n530;
  assign n1342 = ~n403 & n1341;
  assign n1343 = ~n529 & n1342;
  assign n1344 = ~n527 & n1343;
  assign n1345 = ~n525 & n1344;
  assign n1346 = ~\V133(10)  & n1345;
  assign n1347 = ~\V133(7)  & n1346;
  assign n1348 = ~\V133(9)  & n1347;
  assign n1349 = ~\V133(4)  & n1348;
  assign n1350 = ~\V133(3)  & n1349;
  assign n1351 = \V133(2)  & n1350;
  assign n1352 = \V133(1)  & n1351;
  assign n1353 = ~\V133(10)  & n1352;
  assign n1354 = \V116(31)  & ~\V133(10) ;
  assign n1355 = ~n525 & n1354;
  assign n1356 = ~n527 & n1355;
  assign n1357 = ~n529 & n1356;
  assign n1358 = ~n403 & n1357;
  assign n1359 = n530 & n1358;
  assign n1360 = \V47(16)  & n421;
  assign n1361 = n424 & n1360;
  assign n1362 = n434 & n1361;
  assign n1363 = ~n440 & n1362;
  assign n1364 = \V47(20)  & n434;
  assign n1365 = n424 & n1364;
  assign n1366 = ~n421 & n1365;
  assign n1367 = \V47(23)  & ~n434;
  assign n1368 = n424 & n1367;
  assign n1369 = \V47(31)  & ~n424;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1366 & n1370;
  assign n1372 = ~n1363 & n1371;
  assign n1373 = ~n443 & n1372;
  assign n1374 = ~n403 & ~n1373;
  assign n1375 = ~n529 & n1374;
  assign n1376 = ~n527 & n1375;
  assign n1377 = ~n525 & n1376;
  assign n1378 = \V133(10)  & n1377;
  assign n1379 = ~n525 & ~n1373;
  assign n1380 = ~n527 & n1379;
  assign n1381 = ~n529 & n1380;
  assign n1382 = n403 & n1381;
  assign n1383 = ~n529 & ~n1373;
  assign n1384 = ~n527 & n1383;
  assign n1385 = n525 & n1384;
  assign n1386 = n529 & ~n1373;
  assign n1387 = ~n527 & n1386;
  assign n1388 = n527 & ~n1373;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1385 & n1389;
  assign n1391 = ~n1382 & n1390;
  assign n1392 = ~n1378 & n1391;
  assign n1393 = ~n1359 & n1392;
  assign \V165(14)  = n1353 | ~n1393;
  assign n1395 = ~n885 & n1154;
  assign n1396 = ~n882 & n1395;
  assign n1397 = ~n878 & n1396;
  assign n1398 = ~n876 & n1397;
  assign n1399 = ~n873 & n1398;
  assign n1400 = \V133(9)  & n1399;
  assign n1401 = ~\V133(10)  & n1400;
  assign n1402 = \V84(14)  & n421;
  assign n1403 = n424 & n1402;
  assign n1404 = n434 & n1403;
  assign n1405 = ~n440 & n1404;
  assign n1406 = \V84(18)  & n434;
  assign n1407 = n424 & n1406;
  assign n1408 = ~n421 & n1407;
  assign n1409 = \V84(21)  & ~n434;
  assign n1410 = n424 & n1409;
  assign n1411 = \V84(29)  & ~n424;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~n1408 & n1412;
  assign n1414 = ~n1405 & n1413;
  assign n1415 = ~n443 & n1414;
  assign n1416 = ~n873 & ~n1415;
  assign n1417 = ~n876 & n1416;
  assign n1418 = ~n878 & n1417;
  assign n1419 = ~n882 & n1418;
  assign n1420 = ~n885 & n1419;
  assign n1421 = \V133(10)  & n1420;
  assign n1422 = ~n885 & ~n1415;
  assign n1423 = ~n882 & n1422;
  assign n1424 = ~n878 & n1423;
  assign n1425 = ~n876 & n1424;
  assign n1426 = n873 & n1425;
  assign n1427 = ~n876 & ~n1415;
  assign n1428 = ~n878 & n1427;
  assign n1429 = ~n882 & n1428;
  assign n1430 = n885 & n1429;
  assign n1431 = ~n882 & ~n1415;
  assign n1432 = ~n878 & n1431;
  assign n1433 = n876 & n1432;
  assign n1434 = n882 & ~n1415;
  assign n1435 = ~n878 & n1434;
  assign n1436 = n878 & ~n1415;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1433 & n1437;
  assign n1439 = ~n1430 & n1438;
  assign n1440 = ~n1426 & n1439;
  assign n1441 = ~n1421 & n1440;
  assign \V197(29)  = n1401 | ~n1441;
  assign n1443 = \V116(1)  & ~\V133(10) ;
  assign n1444 = ~n885 & n1443;
  assign n1445 = ~n882 & n1444;
  assign n1446 = ~n878 & n1445;
  assign n1447 = ~n876 & n1446;
  assign n1448 = ~n873 & n1447;
  assign n1449 = \V133(9)  & n1448;
  assign n1450 = ~\V133(10)  & n1449;
  assign n1451 = \V47(18)  & n421;
  assign n1452 = n424 & n1451;
  assign n1453 = n434 & n1452;
  assign n1454 = ~n440 & n1453;
  assign n1455 = \V47(22)  & n434;
  assign n1456 = n424 & n1455;
  assign n1457 = ~n421 & n1456;
  assign n1458 = \V47(25)  & ~n434;
  assign n1459 = n424 & n1458;
  assign n1460 = \V84(1)  & ~n424;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1457 & n1461;
  assign n1463 = ~n1454 & n1462;
  assign n1464 = ~n443 & n1463;
  assign n1465 = ~n873 & ~n1464;
  assign n1466 = ~n876 & n1465;
  assign n1467 = ~n878 & n1466;
  assign n1468 = ~n882 & n1467;
  assign n1469 = ~n885 & n1468;
  assign n1470 = \V133(10)  & n1469;
  assign n1471 = ~n885 & ~n1464;
  assign n1472 = ~n882 & n1471;
  assign n1473 = ~n878 & n1472;
  assign n1474 = ~n876 & n1473;
  assign n1475 = n873 & n1474;
  assign n1476 = ~n876 & ~n1464;
  assign n1477 = ~n878 & n1476;
  assign n1478 = ~n882 & n1477;
  assign n1479 = n885 & n1478;
  assign n1480 = ~n882 & ~n1464;
  assign n1481 = ~n878 & n1480;
  assign n1482 = n876 & n1481;
  assign n1483 = n882 & ~n1464;
  assign n1484 = ~n878 & n1483;
  assign n1485 = n878 & ~n1464;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = ~n1482 & n1486;
  assign n1488 = ~n1479 & n1487;
  assign n1489 = ~n1475 & n1488;
  assign n1490 = ~n1470 & n1489;
  assign \V197(1)  = n1450 | ~n1490;
  assign n1492 = n832 & ~n885;
  assign n1493 = ~n882 & n1492;
  assign n1494 = ~n878 & n1493;
  assign n1495 = ~n876 & n1494;
  assign n1496 = ~n873 & n1495;
  assign n1497 = \V133(9)  & n1496;
  assign n1498 = ~\V133(10)  & n1497;
  assign n1499 = \V84(13)  & n421;
  assign n1500 = n424 & n1499;
  assign n1501 = n434 & n1500;
  assign n1502 = ~n440 & n1501;
  assign n1503 = \V84(17)  & n434;
  assign n1504 = n424 & n1503;
  assign n1505 = ~n421 & n1504;
  assign n1506 = \V84(20)  & ~n434;
  assign n1507 = n424 & n1506;
  assign n1508 = \V84(28)  & ~n424;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n1505 & n1509;
  assign n1511 = ~n1502 & n1510;
  assign n1512 = ~n443 & n1511;
  assign n1513 = ~n873 & ~n1512;
  assign n1514 = ~n876 & n1513;
  assign n1515 = ~n878 & n1514;
  assign n1516 = ~n882 & n1515;
  assign n1517 = ~n885 & n1516;
  assign n1518 = \V133(10)  & n1517;
  assign n1519 = ~n885 & ~n1512;
  assign n1520 = ~n882 & n1519;
  assign n1521 = ~n878 & n1520;
  assign n1522 = ~n876 & n1521;
  assign n1523 = n873 & n1522;
  assign n1524 = ~n876 & ~n1512;
  assign n1525 = ~n878 & n1524;
  assign n1526 = ~n882 & n1525;
  assign n1527 = n885 & n1526;
  assign n1528 = ~n882 & ~n1512;
  assign n1529 = ~n878 & n1528;
  assign n1530 = n876 & n1529;
  assign n1531 = n882 & ~n1512;
  assign n1532 = ~n878 & n1531;
  assign n1533 = n878 & ~n1512;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = ~n1530 & n1534;
  assign n1536 = ~n1527 & n1535;
  assign n1537 = ~n1523 & n1536;
  assign n1538 = ~n1518 & n1537;
  assign \V197(28)  = n1498 | ~n1538;
  assign n1540 = \V116(0)  & ~\V133(10) ;
  assign n1541 = ~n885 & n1540;
  assign n1542 = ~n882 & n1541;
  assign n1543 = ~n878 & n1542;
  assign n1544 = ~n876 & n1543;
  assign n1545 = ~n873 & n1544;
  assign n1546 = \V133(9)  & n1545;
  assign n1547 = ~\V133(10)  & n1546;
  assign n1548 = \V47(17)  & n421;
  assign n1549 = n424 & n1548;
  assign n1550 = n434 & n1549;
  assign n1551 = ~n440 & n1550;
  assign n1552 = \V47(21)  & n434;
  assign n1553 = n424 & n1552;
  assign n1554 = ~n421 & n1553;
  assign n1555 = \V47(24)  & ~n434;
  assign n1556 = n424 & n1555;
  assign n1557 = \V84(0)  & ~n424;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~n1554 & n1558;
  assign n1560 = ~n1551 & n1559;
  assign n1561 = ~n443 & n1560;
  assign n1562 = ~n873 & ~n1561;
  assign n1563 = ~n876 & n1562;
  assign n1564 = ~n878 & n1563;
  assign n1565 = ~n882 & n1564;
  assign n1566 = ~n885 & n1565;
  assign n1567 = \V133(10)  & n1566;
  assign n1568 = ~n885 & ~n1561;
  assign n1569 = ~n882 & n1568;
  assign n1570 = ~n878 & n1569;
  assign n1571 = ~n876 & n1570;
  assign n1572 = n873 & n1571;
  assign n1573 = ~n876 & ~n1561;
  assign n1574 = ~n878 & n1573;
  assign n1575 = ~n882 & n1574;
  assign n1576 = n885 & n1575;
  assign n1577 = ~n882 & ~n1561;
  assign n1578 = ~n878 & n1577;
  assign n1579 = n876 & n1578;
  assign n1580 = n882 & ~n1561;
  assign n1581 = ~n878 & n1580;
  assign n1582 = n878 & ~n1561;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1579 & n1583;
  assign n1585 = ~n1576 & n1584;
  assign n1586 = ~n1572 & n1585;
  assign n1587 = ~n1567 & n1586;
  assign \V197(0)  = n1547 | ~n1587;
  assign n1589 = \V116(7)  & ~\V133(10) ;
  assign n1590 = ~n885 & n1589;
  assign n1591 = ~n882 & n1590;
  assign n1592 = ~n878 & n1591;
  assign n1593 = ~n876 & n1592;
  assign n1594 = ~n873 & n1593;
  assign n1595 = \V133(9)  & n1594;
  assign n1596 = ~\V133(10)  & n1595;
  assign n1597 = \V47(24)  & n421;
  assign n1598 = n424 & n1597;
  assign n1599 = n434 & n1598;
  assign n1600 = ~n440 & n1599;
  assign n1601 = \V47(28)  & n434;
  assign n1602 = n424 & n1601;
  assign n1603 = ~n421 & n1602;
  assign n1604 = \V47(31)  & ~n434;
  assign n1605 = n424 & n1604;
  assign n1606 = \V84(7)  & ~n424;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1603 & n1607;
  assign n1609 = ~n1600 & n1608;
  assign n1610 = ~n443 & n1609;
  assign n1611 = ~n873 & ~n1610;
  assign n1612 = ~n876 & n1611;
  assign n1613 = ~n878 & n1612;
  assign n1614 = ~n882 & n1613;
  assign n1615 = ~n885 & n1614;
  assign n1616 = \V133(10)  & n1615;
  assign n1617 = ~n885 & ~n1610;
  assign n1618 = ~n882 & n1617;
  assign n1619 = ~n878 & n1618;
  assign n1620 = ~n876 & n1619;
  assign n1621 = n873 & n1620;
  assign n1622 = ~n876 & ~n1610;
  assign n1623 = ~n878 & n1622;
  assign n1624 = ~n882 & n1623;
  assign n1625 = n885 & n1624;
  assign n1626 = ~n882 & ~n1610;
  assign n1627 = ~n878 & n1626;
  assign n1628 = n876 & n1627;
  assign n1629 = n882 & ~n1610;
  assign n1630 = ~n878 & n1629;
  assign n1631 = n878 & ~n1610;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~n1628 & n1632;
  assign n1634 = ~n1625 & n1633;
  assign n1635 = ~n1621 & n1634;
  assign n1636 = ~n1616 & n1635;
  assign \V197(7)  = n1596 | ~n1636;
  assign n1638 = \V116(6)  & ~\V133(10) ;
  assign n1639 = ~n885 & n1638;
  assign n1640 = ~n882 & n1639;
  assign n1641 = ~n878 & n1640;
  assign n1642 = ~n876 & n1641;
  assign n1643 = ~n873 & n1642;
  assign n1644 = \V133(9)  & n1643;
  assign n1645 = ~\V133(10)  & n1644;
  assign n1646 = \V47(23)  & n421;
  assign n1647 = n424 & n1646;
  assign n1648 = n434 & n1647;
  assign n1649 = ~n440 & n1648;
  assign n1650 = \V47(27)  & n434;
  assign n1651 = n424 & n1650;
  assign n1652 = ~n421 & n1651;
  assign n1653 = \V47(30)  & ~n434;
  assign n1654 = n424 & n1653;
  assign n1655 = \V84(6)  & ~n424;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1652 & n1656;
  assign n1658 = ~n1649 & n1657;
  assign n1659 = ~n443 & n1658;
  assign n1660 = ~n873 & ~n1659;
  assign n1661 = ~n876 & n1660;
  assign n1662 = ~n878 & n1661;
  assign n1663 = ~n882 & n1662;
  assign n1664 = ~n885 & n1663;
  assign n1665 = \V133(10)  & n1664;
  assign n1666 = ~n885 & ~n1659;
  assign n1667 = ~n882 & n1666;
  assign n1668 = ~n878 & n1667;
  assign n1669 = ~n876 & n1668;
  assign n1670 = n873 & n1669;
  assign n1671 = ~n876 & ~n1659;
  assign n1672 = ~n878 & n1671;
  assign n1673 = ~n882 & n1672;
  assign n1674 = n885 & n1673;
  assign n1675 = ~n882 & ~n1659;
  assign n1676 = ~n878 & n1675;
  assign n1677 = n876 & n1676;
  assign n1678 = n882 & ~n1659;
  assign n1679 = ~n878 & n1678;
  assign n1680 = n878 & ~n1659;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n1677 & n1681;
  assign n1683 = ~n1674 & n1682;
  assign n1684 = ~n1670 & n1683;
  assign n1685 = ~n1665 & n1684;
  assign \V197(6)  = n1645 | ~n1685;
  assign n1687 = ~\V133(10)  & \V116(21) ;
  assign n1688 = ~n885 & n1687;
  assign n1689 = ~n882 & n1688;
  assign n1690 = ~n878 & n1689;
  assign n1691 = ~n876 & n1690;
  assign n1692 = ~n873 & n1691;
  assign n1693 = \V133(9)  & n1692;
  assign n1694 = ~\V133(10)  & n1693;
  assign n1695 = \V84(6)  & n421;
  assign n1696 = n424 & n1695;
  assign n1697 = n434 & n1696;
  assign n1698 = ~n440 & n1697;
  assign n1699 = \V84(13)  & ~n434;
  assign n1700 = n424 & n1699;
  assign n1701 = \V84(21)  & ~n424;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n508 & n1702;
  assign n1704 = ~n1698 & n1703;
  assign n1705 = ~n443 & n1704;
  assign n1706 = ~n873 & ~n1705;
  assign n1707 = ~n876 & n1706;
  assign n1708 = ~n878 & n1707;
  assign n1709 = ~n882 & n1708;
  assign n1710 = ~n885 & n1709;
  assign n1711 = \V133(10)  & n1710;
  assign n1712 = ~n885 & ~n1705;
  assign n1713 = ~n882 & n1712;
  assign n1714 = ~n878 & n1713;
  assign n1715 = ~n876 & n1714;
  assign n1716 = n873 & n1715;
  assign n1717 = ~n876 & ~n1705;
  assign n1718 = ~n878 & n1717;
  assign n1719 = ~n882 & n1718;
  assign n1720 = n885 & n1719;
  assign n1721 = ~n882 & ~n1705;
  assign n1722 = ~n878 & n1721;
  assign n1723 = n876 & n1722;
  assign n1724 = n882 & ~n1705;
  assign n1725 = ~n878 & n1724;
  assign n1726 = n878 & ~n1705;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1723 & n1727;
  assign n1729 = ~n1720 & n1728;
  assign n1730 = ~n1716 & n1729;
  assign n1731 = ~n1711 & n1730;
  assign \V197(21)  = n1694 | ~n1731;
  assign n1733 = n405 & ~n885;
  assign n1734 = ~n882 & n1733;
  assign n1735 = ~n878 & n1734;
  assign n1736 = ~n876 & n1735;
  assign n1737 = ~n873 & n1736;
  assign n1738 = \V133(9)  & n1737;
  assign n1739 = ~\V133(10)  & n1738;
  assign n1740 = \V47(26)  & n421;
  assign n1741 = n424 & n1740;
  assign n1742 = n434 & n1741;
  assign n1743 = ~n440 & n1742;
  assign n1744 = \V47(30)  & n434;
  assign n1745 = n424 & n1744;
  assign n1746 = ~n421 & n1745;
  assign n1747 = \V84(1)  & ~n434;
  assign n1748 = n424 & n1747;
  assign n1749 = \V84(9)  & ~n424;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = ~n1746 & n1750;
  assign n1752 = ~n1743 & n1751;
  assign n1753 = ~n443 & n1752;
  assign n1754 = ~n873 & ~n1753;
  assign n1755 = ~n876 & n1754;
  assign n1756 = ~n878 & n1755;
  assign n1757 = ~n882 & n1756;
  assign n1758 = ~n885 & n1757;
  assign n1759 = \V133(10)  & n1758;
  assign n1760 = ~n885 & ~n1753;
  assign n1761 = ~n882 & n1760;
  assign n1762 = ~n878 & n1761;
  assign n1763 = ~n876 & n1762;
  assign n1764 = n873 & n1763;
  assign n1765 = ~n876 & ~n1753;
  assign n1766 = ~n878 & n1765;
  assign n1767 = ~n882 & n1766;
  assign n1768 = n885 & n1767;
  assign n1769 = ~n882 & ~n1753;
  assign n1770 = ~n878 & n1769;
  assign n1771 = n876 & n1770;
  assign n1772 = n882 & ~n1753;
  assign n1773 = ~n878 & n1772;
  assign n1774 = n878 & ~n1753;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1771 & n1775;
  assign n1777 = ~n1768 & n1776;
  assign n1778 = ~n1764 & n1777;
  assign n1779 = ~n1759 & n1778;
  assign \V197(9)  = n1739 | ~n1779;
  assign n1781 = ~\V133(10)  & \V116(20) ;
  assign n1782 = ~n885 & n1781;
  assign n1783 = ~n882 & n1782;
  assign n1784 = ~n878 & n1783;
  assign n1785 = ~n876 & n1784;
  assign n1786 = ~n873 & n1785;
  assign n1787 = \V133(9)  & n1786;
  assign n1788 = ~\V133(10)  & n1787;
  assign n1789 = \V84(5)  & n421;
  assign n1790 = n424 & n1789;
  assign n1791 = n434 & n1790;
  assign n1792 = ~n440 & n1791;
  assign n1793 = \V84(12)  & ~n434;
  assign n1794 = n424 & n1793;
  assign n1795 = \V84(20)  & ~n424;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~n450 & n1796;
  assign n1798 = ~n1792 & n1797;
  assign n1799 = ~n443 & n1798;
  assign n1800 = ~n873 & ~n1799;
  assign n1801 = ~n876 & n1800;
  assign n1802 = ~n878 & n1801;
  assign n1803 = ~n882 & n1802;
  assign n1804 = ~n885 & n1803;
  assign n1805 = \V133(10)  & n1804;
  assign n1806 = ~n885 & ~n1799;
  assign n1807 = ~n882 & n1806;
  assign n1808 = ~n878 & n1807;
  assign n1809 = ~n876 & n1808;
  assign n1810 = n873 & n1809;
  assign n1811 = ~n876 & ~n1799;
  assign n1812 = ~n878 & n1811;
  assign n1813 = ~n882 & n1812;
  assign n1814 = n885 & n1813;
  assign n1815 = ~n882 & ~n1799;
  assign n1816 = ~n878 & n1815;
  assign n1817 = n876 & n1816;
  assign n1818 = n882 & ~n1799;
  assign n1819 = ~n878 & n1818;
  assign n1820 = n878 & ~n1799;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1817 & n1821;
  assign n1823 = ~n1814 & n1822;
  assign n1824 = ~n1810 & n1823;
  assign n1825 = ~n1805 & n1824;
  assign \V197(20)  = n1788 | ~n1825;
  assign n1827 = \V116(8)  & ~\V133(10) ;
  assign n1828 = ~n885 & n1827;
  assign n1829 = ~n882 & n1828;
  assign n1830 = ~n878 & n1829;
  assign n1831 = ~n876 & n1830;
  assign n1832 = ~n873 & n1831;
  assign n1833 = \V133(9)  & n1832;
  assign n1834 = ~\V133(10)  & n1833;
  assign n1835 = \V47(25)  & n421;
  assign n1836 = n424 & n1835;
  assign n1837 = n434 & n1836;
  assign n1838 = ~n440 & n1837;
  assign n1839 = \V47(29)  & n434;
  assign n1840 = n424 & n1839;
  assign n1841 = ~n421 & n1840;
  assign n1842 = \V84(0)  & ~n434;
  assign n1843 = n424 & n1842;
  assign n1844 = \V84(8)  & ~n424;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1841 & n1845;
  assign n1847 = ~n1838 & n1846;
  assign n1848 = ~n443 & n1847;
  assign n1849 = ~n873 & ~n1848;
  assign n1850 = ~n876 & n1849;
  assign n1851 = ~n878 & n1850;
  assign n1852 = ~n882 & n1851;
  assign n1853 = ~n885 & n1852;
  assign n1854 = \V133(10)  & n1853;
  assign n1855 = ~n885 & ~n1848;
  assign n1856 = ~n882 & n1855;
  assign n1857 = ~n878 & n1856;
  assign n1858 = ~n876 & n1857;
  assign n1859 = n873 & n1858;
  assign n1860 = ~n876 & ~n1848;
  assign n1861 = ~n878 & n1860;
  assign n1862 = ~n882 & n1861;
  assign n1863 = n885 & n1862;
  assign n1864 = ~n882 & ~n1848;
  assign n1865 = ~n878 & n1864;
  assign n1866 = n876 & n1865;
  assign n1867 = n882 & ~n1848;
  assign n1868 = ~n878 & n1867;
  assign n1869 = n878 & ~n1848;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = ~n1866 & n1870;
  assign n1872 = ~n1863 & n1871;
  assign n1873 = ~n1859 & n1872;
  assign n1874 = ~n1854 & n1873;
  assign \V197(8)  = n1834 | ~n1874;
  assign n1876 = ~\V133(10)  & \V116(23) ;
  assign n1877 = ~n885 & n1876;
  assign n1878 = ~n882 & n1877;
  assign n1879 = ~n878 & n1878;
  assign n1880 = ~n876 & n1879;
  assign n1881 = ~n873 & n1880;
  assign n1882 = \V133(9)  & n1881;
  assign n1883 = ~\V133(10)  & n1882;
  assign n1884 = \V84(8)  & n421;
  assign n1885 = n424 & n1884;
  assign n1886 = n434 & n1885;
  assign n1887 = ~n440 & n1886;
  assign n1888 = \V84(12)  & n434;
  assign n1889 = n424 & n1888;
  assign n1890 = ~n421 & n1889;
  assign n1891 = \V84(15)  & ~n434;
  assign n1892 = n424 & n1891;
  assign n1893 = \V84(23)  & ~n424;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~n1890 & n1894;
  assign n1896 = ~n1887 & n1895;
  assign n1897 = ~n443 & n1896;
  assign n1898 = ~n873 & ~n1897;
  assign n1899 = ~n876 & n1898;
  assign n1900 = ~n878 & n1899;
  assign n1901 = ~n882 & n1900;
  assign n1902 = ~n885 & n1901;
  assign n1903 = \V133(10)  & n1902;
  assign n1904 = ~n885 & ~n1897;
  assign n1905 = ~n882 & n1904;
  assign n1906 = ~n878 & n1905;
  assign n1907 = ~n876 & n1906;
  assign n1908 = n873 & n1907;
  assign n1909 = ~n876 & ~n1897;
  assign n1910 = ~n878 & n1909;
  assign n1911 = ~n882 & n1910;
  assign n1912 = n885 & n1911;
  assign n1913 = ~n882 & ~n1897;
  assign n1914 = ~n878 & n1913;
  assign n1915 = n876 & n1914;
  assign n1916 = n882 & ~n1897;
  assign n1917 = ~n878 & n1916;
  assign n1918 = n878 & ~n1897;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = ~n1915 & n1919;
  assign n1921 = ~n1912 & n1920;
  assign n1922 = ~n1908 & n1921;
  assign n1923 = ~n1903 & n1922;
  assign \V197(23)  = n1883 | ~n1923;
  assign n1925 = ~\V133(10)  & \V116(22) ;
  assign n1926 = ~n885 & n1925;
  assign n1927 = ~n882 & n1926;
  assign n1928 = ~n878 & n1927;
  assign n1929 = ~n876 & n1928;
  assign n1930 = ~n873 & n1929;
  assign n1931 = \V133(9)  & n1930;
  assign n1932 = ~\V133(10)  & n1931;
  assign n1933 = \V84(7)  & n421;
  assign n1934 = n424 & n1933;
  assign n1935 = n434 & n1934;
  assign n1936 = ~n440 & n1935;
  assign n1937 = \V84(14)  & ~n434;
  assign n1938 = n424 & n1937;
  assign n1939 = \V84(22)  & ~n424;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n480 & n1940;
  assign n1942 = ~n1936 & n1941;
  assign n1943 = ~n443 & n1942;
  assign n1944 = ~n873 & ~n1943;
  assign n1945 = ~n876 & n1944;
  assign n1946 = ~n878 & n1945;
  assign n1947 = ~n882 & n1946;
  assign n1948 = ~n885 & n1947;
  assign n1949 = \V133(10)  & n1948;
  assign n1950 = ~n885 & ~n1943;
  assign n1951 = ~n882 & n1950;
  assign n1952 = ~n878 & n1951;
  assign n1953 = ~n876 & n1952;
  assign n1954 = n873 & n1953;
  assign n1955 = ~n876 & ~n1943;
  assign n1956 = ~n878 & n1955;
  assign n1957 = ~n882 & n1956;
  assign n1958 = n885 & n1957;
  assign n1959 = ~n882 & ~n1943;
  assign n1960 = ~n878 & n1959;
  assign n1961 = n876 & n1960;
  assign n1962 = n882 & ~n1943;
  assign n1963 = ~n878 & n1962;
  assign n1964 = n878 & ~n1943;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n1961 & n1965;
  assign n1967 = ~n1958 & n1966;
  assign n1968 = ~n1954 & n1967;
  assign n1969 = ~n1949 & n1968;
  assign \V197(22)  = n1932 | ~n1969;
  assign n1971 = ~\V133(10)  & \V116(25) ;
  assign n1972 = ~n885 & n1971;
  assign n1973 = ~n882 & n1972;
  assign n1974 = ~n878 & n1973;
  assign n1975 = ~n876 & n1974;
  assign n1976 = ~n873 & n1975;
  assign n1977 = \V133(9)  & n1976;
  assign n1978 = ~\V133(10)  & n1977;
  assign n1979 = \V84(10)  & n421;
  assign n1980 = n424 & n1979;
  assign n1981 = n434 & n1980;
  assign n1982 = ~n440 & n1981;
  assign n1983 = \V84(14)  & n434;
  assign n1984 = n424 & n1983;
  assign n1985 = ~n421 & n1984;
  assign n1986 = \V84(17)  & ~n434;
  assign n1987 = n424 & n1986;
  assign n1988 = \V84(25)  & ~n424;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1985 & n1989;
  assign n1991 = ~n1982 & n1990;
  assign n1992 = ~n443 & n1991;
  assign n1993 = ~n873 & ~n1992;
  assign n1994 = ~n876 & n1993;
  assign n1995 = ~n878 & n1994;
  assign n1996 = ~n882 & n1995;
  assign n1997 = ~n885 & n1996;
  assign n1998 = \V133(10)  & n1997;
  assign n1999 = ~n885 & ~n1992;
  assign n2000 = ~n882 & n1999;
  assign n2001 = ~n878 & n2000;
  assign n2002 = ~n876 & n2001;
  assign n2003 = n873 & n2002;
  assign n2004 = ~n876 & ~n1992;
  assign n2005 = ~n878 & n2004;
  assign n2006 = ~n882 & n2005;
  assign n2007 = n885 & n2006;
  assign n2008 = ~n882 & ~n1992;
  assign n2009 = ~n878 & n2008;
  assign n2010 = n876 & n2009;
  assign n2011 = n882 & ~n1992;
  assign n2012 = ~n878 & n2011;
  assign n2013 = n878 & ~n1992;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n2010 & n2014;
  assign n2016 = ~n2007 & n2015;
  assign n2017 = ~n2003 & n2016;
  assign n2018 = ~n1998 & n2017;
  assign \V197(25)  = n1978 | ~n2018;
  assign n2020 = ~\V133(10)  & \V116(24) ;
  assign n2021 = ~n885 & n2020;
  assign n2022 = ~n882 & n2021;
  assign n2023 = ~n878 & n2022;
  assign n2024 = ~n876 & n2023;
  assign n2025 = ~n873 & n2024;
  assign n2026 = \V133(9)  & n2025;
  assign n2027 = ~\V133(10)  & n2026;
  assign n2028 = \V84(9)  & n421;
  assign n2029 = n424 & n2028;
  assign n2030 = n434 & n2029;
  assign n2031 = ~n440 & n2030;
  assign n2032 = \V84(13)  & n434;
  assign n2033 = n424 & n2032;
  assign n2034 = ~n421 & n2033;
  assign n2035 = \V84(16)  & ~n434;
  assign n2036 = n424 & n2035;
  assign n2037 = \V84(24)  & ~n424;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~n2034 & n2038;
  assign n2040 = ~n2031 & n2039;
  assign n2041 = ~n443 & n2040;
  assign n2042 = ~n873 & ~n2041;
  assign n2043 = ~n876 & n2042;
  assign n2044 = ~n878 & n2043;
  assign n2045 = ~n882 & n2044;
  assign n2046 = ~n885 & n2045;
  assign n2047 = \V133(10)  & n2046;
  assign n2048 = ~n885 & ~n2041;
  assign n2049 = ~n882 & n2048;
  assign n2050 = ~n878 & n2049;
  assign n2051 = ~n876 & n2050;
  assign n2052 = n873 & n2051;
  assign n2053 = ~n876 & ~n2041;
  assign n2054 = ~n878 & n2053;
  assign n2055 = ~n882 & n2054;
  assign n2056 = n885 & n2055;
  assign n2057 = ~n882 & ~n2041;
  assign n2058 = ~n878 & n2057;
  assign n2059 = n876 & n2058;
  assign n2060 = n882 & ~n2041;
  assign n2061 = ~n878 & n2060;
  assign n2062 = n878 & ~n2041;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2059 & n2063;
  assign n2065 = ~n2056 & n2064;
  assign n2066 = ~n2052 & n2065;
  assign n2067 = ~n2047 & n2066;
  assign \V197(24)  = n2027 | ~n2067;
  assign n2069 = ~\V133(8)  & n391;
  assign n2070 = \V133(7)  & n2069;
  assign n2071 = ~n394 & n724;
  assign n2072 = ~n2070 & n2071;
  assign n2073 = ~n530 & n2072;
  assign n2074 = ~\V133(10)  & n2073;
  assign n2075 = \V119(0)  & ~n394;
  assign n2076 = ~n2070 & n2075;
  assign n2077 = ~n530 & n2076;
  assign n2078 = \V133(10)  & n2077;
  assign n2079 = ~\V133(10)  & n731;
  assign n2080 = ~n530 & n2079;
  assign n2081 = ~n2070 & n2080;
  assign n2082 = ~n394 & n2081;
  assign n2083 = ~n724 & n2082;
  assign n2084 = ~\V133(10)  & ~n731;
  assign n2085 = ~n530 & n2084;
  assign n2086 = ~n2070 & n2085;
  assign n2087 = ~n394 & n2086;
  assign n2088 = ~n724 & n2087;
  assign n2089 = \V121(16)  & n2070;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = ~n2083 & n2090;
  assign n2092 = ~n2078 & n2091;
  assign \V213(0)  = n2074 | ~n2092;
  assign n2094 = ~\V133(10)  & \V116(17) ;
  assign n2095 = ~n885 & n2094;
  assign n2096 = ~n882 & n2095;
  assign n2097 = ~n878 & n2096;
  assign n2098 = ~n876 & n2097;
  assign n2099 = ~n873 & n2098;
  assign n2100 = \V133(9)  & n2099;
  assign n2101 = ~\V133(10)  & n2100;
  assign n2102 = \V84(2)  & n421;
  assign n2103 = n424 & n2102;
  assign n2104 = n434 & n2103;
  assign n2105 = ~n440 & n2104;
  assign n2106 = \V84(6)  & n434;
  assign n2107 = n424 & n2106;
  assign n2108 = ~n421 & n2107;
  assign n2109 = \V84(9)  & ~n434;
  assign n2110 = n424 & n2109;
  assign n2111 = \V84(17)  & ~n424;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~n2108 & n2112;
  assign n2114 = ~n2105 & n2113;
  assign n2115 = ~n443 & n2114;
  assign n2116 = ~n873 & ~n2115;
  assign n2117 = ~n876 & n2116;
  assign n2118 = ~n878 & n2117;
  assign n2119 = ~n882 & n2118;
  assign n2120 = ~n885 & n2119;
  assign n2121 = \V133(10)  & n2120;
  assign n2122 = ~n885 & ~n2115;
  assign n2123 = ~n882 & n2122;
  assign n2124 = ~n878 & n2123;
  assign n2125 = ~n876 & n2124;
  assign n2126 = n873 & n2125;
  assign n2127 = ~n876 & ~n2115;
  assign n2128 = ~n878 & n2127;
  assign n2129 = ~n882 & n2128;
  assign n2130 = n885 & n2129;
  assign n2131 = ~n882 & ~n2115;
  assign n2132 = ~n878 & n2131;
  assign n2133 = n876 & n2132;
  assign n2134 = n882 & ~n2115;
  assign n2135 = ~n878 & n2134;
  assign n2136 = n878 & ~n2115;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2133 & n2137;
  assign n2139 = ~n2130 & n2138;
  assign n2140 = ~n2126 & n2139;
  assign n2141 = ~n2121 & n2140;
  assign \V197(17)  = n2101 | ~n2141;
  assign n2143 = ~\V133(10)  & \V116(16) ;
  assign n2144 = ~n885 & n2143;
  assign n2145 = ~n882 & n2144;
  assign n2146 = ~n878 & n2145;
  assign n2147 = ~n876 & n2146;
  assign n2148 = ~n873 & n2147;
  assign n2149 = \V133(9)  & n2148;
  assign n2150 = ~\V133(10)  & n2149;
  assign n2151 = \V84(1)  & n421;
  assign n2152 = n424 & n2151;
  assign n2153 = n434 & n2152;
  assign n2154 = ~n440 & n2153;
  assign n2155 = \V84(5)  & n434;
  assign n2156 = n424 & n2155;
  assign n2157 = ~n421 & n2156;
  assign n2158 = \V84(8)  & ~n434;
  assign n2159 = n424 & n2158;
  assign n2160 = \V84(16)  & ~n424;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n2157 & n2161;
  assign n2163 = ~n2154 & n2162;
  assign n2164 = ~n443 & n2163;
  assign n2165 = ~n873 & ~n2164;
  assign n2166 = ~n876 & n2165;
  assign n2167 = ~n878 & n2166;
  assign n2168 = ~n882 & n2167;
  assign n2169 = ~n885 & n2168;
  assign n2170 = \V133(10)  & n2169;
  assign n2171 = ~n885 & ~n2164;
  assign n2172 = ~n882 & n2171;
  assign n2173 = ~n878 & n2172;
  assign n2174 = ~n876 & n2173;
  assign n2175 = n873 & n2174;
  assign n2176 = ~n876 & ~n2164;
  assign n2177 = ~n878 & n2176;
  assign n2178 = ~n882 & n2177;
  assign n2179 = n885 & n2178;
  assign n2180 = ~n882 & ~n2164;
  assign n2181 = ~n878 & n2180;
  assign n2182 = n876 & n2181;
  assign n2183 = n882 & ~n2164;
  assign n2184 = ~n878 & n2183;
  assign n2185 = n878 & ~n2164;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2182 & n2186;
  assign n2188 = ~n2179 & n2187;
  assign n2189 = ~n2175 & n2188;
  assign n2190 = ~n2170 & n2189;
  assign \V197(16)  = n2150 | ~n2190;
  assign n2192 = ~\V133(10)  & \V116(19) ;
  assign n2193 = ~n885 & n2192;
  assign n2194 = ~n882 & n2193;
  assign n2195 = ~n878 & n2194;
  assign n2196 = ~n876 & n2195;
  assign n2197 = ~n873 & n2196;
  assign n2198 = \V133(9)  & n2197;
  assign n2199 = ~\V133(10)  & n2198;
  assign n2200 = \V84(4)  & n421;
  assign n2201 = n424 & n2200;
  assign n2202 = n434 & n2201;
  assign n2203 = ~n440 & n2202;
  assign n2204 = \V84(8)  & n434;
  assign n2205 = n424 & n2204;
  assign n2206 = ~n421 & n2205;
  assign n2207 = \V84(11)  & ~n434;
  assign n2208 = n424 & n2207;
  assign n2209 = \V84(19)  & ~n424;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = ~n2206 & n2210;
  assign n2212 = ~n2203 & n2211;
  assign n2213 = ~n443 & n2212;
  assign n2214 = ~n873 & ~n2213;
  assign n2215 = ~n876 & n2214;
  assign n2216 = ~n878 & n2215;
  assign n2217 = ~n882 & n2216;
  assign n2218 = ~n885 & n2217;
  assign n2219 = \V133(10)  & n2218;
  assign n2220 = ~n885 & ~n2213;
  assign n2221 = ~n882 & n2220;
  assign n2222 = ~n878 & n2221;
  assign n2223 = ~n876 & n2222;
  assign n2224 = n873 & n2223;
  assign n2225 = ~n876 & ~n2213;
  assign n2226 = ~n878 & n2225;
  assign n2227 = ~n882 & n2226;
  assign n2228 = n885 & n2227;
  assign n2229 = ~n882 & ~n2213;
  assign n2230 = ~n878 & n2229;
  assign n2231 = n876 & n2230;
  assign n2232 = n882 & ~n2213;
  assign n2233 = ~n878 & n2232;
  assign n2234 = n878 & ~n2213;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = ~n2231 & n2235;
  assign n2237 = ~n2228 & n2236;
  assign n2238 = ~n2224 & n2237;
  assign n2239 = ~n2219 & n2238;
  assign \V197(19)  = n2199 | ~n2239;
  assign n2241 = ~\V133(10)  & \V116(18) ;
  assign n2242 = ~n885 & n2241;
  assign n2243 = ~n882 & n2242;
  assign n2244 = ~n878 & n2243;
  assign n2245 = ~n876 & n2244;
  assign n2246 = ~n873 & n2245;
  assign n2247 = \V133(9)  & n2246;
  assign n2248 = ~\V133(10)  & n2247;
  assign n2249 = \V84(3)  & n421;
  assign n2250 = n424 & n2249;
  assign n2251 = n434 & n2250;
  assign n2252 = ~n440 & n2251;
  assign n2253 = \V84(7)  & n434;
  assign n2254 = n424 & n2253;
  assign n2255 = ~n421 & n2254;
  assign n2256 = \V84(10)  & ~n434;
  assign n2257 = n424 & n2256;
  assign n2258 = \V84(18)  & ~n424;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2255 & n2259;
  assign n2261 = ~n2252 & n2260;
  assign n2262 = ~n443 & n2261;
  assign n2263 = ~n873 & ~n2262;
  assign n2264 = ~n876 & n2263;
  assign n2265 = ~n878 & n2264;
  assign n2266 = ~n882 & n2265;
  assign n2267 = ~n885 & n2266;
  assign n2268 = \V133(10)  & n2267;
  assign n2269 = ~n885 & ~n2262;
  assign n2270 = ~n882 & n2269;
  assign n2271 = ~n878 & n2270;
  assign n2272 = ~n876 & n2271;
  assign n2273 = n873 & n2272;
  assign n2274 = ~n876 & ~n2262;
  assign n2275 = ~n878 & n2274;
  assign n2276 = ~n882 & n2275;
  assign n2277 = n885 & n2276;
  assign n2278 = ~n882 & ~n2262;
  assign n2279 = ~n878 & n2278;
  assign n2280 = n876 & n2279;
  assign n2281 = n882 & ~n2262;
  assign n2282 = ~n878 & n2281;
  assign n2283 = n878 & ~n2262;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2280 & n2284;
  assign n2286 = ~n2277 & n2285;
  assign n2287 = ~n2273 & n2286;
  assign n2288 = ~n2268 & n2287;
  assign \V197(18)  = n2248 | ~n2288;
  assign n2290 = n469 & ~n885;
  assign n2291 = ~n882 & n2290;
  assign n2292 = ~n878 & n2291;
  assign n2293 = ~n876 & n2292;
  assign n2294 = ~n873 & n2293;
  assign n2295 = \V133(9)  & n2294;
  assign n2296 = ~\V133(10)  & n2295;
  assign n2297 = \V47(28)  & n421;
  assign n2298 = n424 & n2297;
  assign n2299 = n434 & n2298;
  assign n2300 = ~n440 & n2299;
  assign n2301 = \V84(0)  & n434;
  assign n2302 = n424 & n2301;
  assign n2303 = ~n421 & n2302;
  assign n2304 = \V84(3)  & ~n434;
  assign n2305 = n424 & n2304;
  assign n2306 = \V84(11)  & ~n424;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2303 & n2307;
  assign n2309 = ~n2300 & n2308;
  assign n2310 = ~n443 & n2309;
  assign n2311 = ~n873 & ~n2310;
  assign n2312 = ~n876 & n2311;
  assign n2313 = ~n878 & n2312;
  assign n2314 = ~n882 & n2313;
  assign n2315 = ~n885 & n2314;
  assign n2316 = \V133(10)  & n2315;
  assign n2317 = ~n885 & ~n2310;
  assign n2318 = ~n882 & n2317;
  assign n2319 = ~n878 & n2318;
  assign n2320 = ~n876 & n2319;
  assign n2321 = n873 & n2320;
  assign n2322 = ~n876 & ~n2310;
  assign n2323 = ~n878 & n2322;
  assign n2324 = ~n882 & n2323;
  assign n2325 = n885 & n2324;
  assign n2326 = ~n882 & ~n2310;
  assign n2327 = ~n878 & n2326;
  assign n2328 = n876 & n2327;
  assign n2329 = n882 & ~n2310;
  assign n2330 = ~n878 & n2329;
  assign n2331 = n878 & ~n2310;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = ~n2328 & n2332;
  assign n2334 = ~n2325 & n2333;
  assign n2335 = ~n2321 & n2334;
  assign n2336 = ~n2316 & n2335;
  assign \V197(11)  = n2296 | ~n2336;
  assign n2338 = n497 & ~n885;
  assign n2339 = ~n882 & n2338;
  assign n2340 = ~n878 & n2339;
  assign n2341 = ~n876 & n2340;
  assign n2342 = ~n873 & n2341;
  assign n2343 = \V133(9)  & n2342;
  assign n2344 = ~\V133(10)  & n2343;
  assign n2345 = \V47(27)  & n421;
  assign n2346 = n424 & n2345;
  assign n2347 = n434 & n2346;
  assign n2348 = ~n440 & n2347;
  assign n2349 = \V47(31)  & n434;
  assign n2350 = n424 & n2349;
  assign n2351 = ~n421 & n2350;
  assign n2352 = \V84(2)  & ~n434;
  assign n2353 = n424 & n2352;
  assign n2354 = \V84(10)  & ~n424;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2351 & n2355;
  assign n2357 = ~n2348 & n2356;
  assign n2358 = ~n443 & n2357;
  assign n2359 = ~n873 & ~n2358;
  assign n2360 = ~n876 & n2359;
  assign n2361 = ~n878 & n2360;
  assign n2362 = ~n882 & n2361;
  assign n2363 = ~n885 & n2362;
  assign n2364 = \V133(10)  & n2363;
  assign n2365 = ~n885 & ~n2358;
  assign n2366 = ~n882 & n2365;
  assign n2367 = ~n878 & n2366;
  assign n2368 = ~n876 & n2367;
  assign n2369 = n873 & n2368;
  assign n2370 = ~n876 & ~n2358;
  assign n2371 = ~n878 & n2370;
  assign n2372 = ~n882 & n2371;
  assign n2373 = n885 & n2372;
  assign n2374 = ~n882 & ~n2358;
  assign n2375 = ~n878 & n2374;
  assign n2376 = n876 & n2375;
  assign n2377 = n882 & ~n2358;
  assign n2378 = ~n878 & n2377;
  assign n2379 = n878 & ~n2358;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = ~n2376 & n2380;
  assign n2382 = ~n2373 & n2381;
  assign n2383 = ~n2369 & n2382;
  assign n2384 = ~n2364 & n2383;
  assign \V197(10)  = n2344 | ~n2384;
  assign n2386 = n652 & ~n885;
  assign n2387 = ~n882 & n2386;
  assign n2388 = ~n878 & n2387;
  assign n2389 = ~n876 & n2388;
  assign n2390 = ~n873 & n2389;
  assign n2391 = \V133(9)  & n2390;
  assign n2392 = ~\V133(10)  & n2391;
  assign n2393 = \V47(30)  & n421;
  assign n2394 = n424 & n2393;
  assign n2395 = n434 & n2394;
  assign n2396 = ~n440 & n2395;
  assign n2397 = \V84(5)  & ~n434;
  assign n2398 = n424 & n2397;
  assign n2399 = \V84(13)  & ~n424;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n757 & n2400;
  assign n2402 = ~n2396 & n2401;
  assign n2403 = ~n443 & n2402;
  assign n2404 = ~n873 & ~n2403;
  assign n2405 = ~n876 & n2404;
  assign n2406 = ~n878 & n2405;
  assign n2407 = ~n882 & n2406;
  assign n2408 = ~n885 & n2407;
  assign n2409 = \V133(10)  & n2408;
  assign n2410 = ~n885 & ~n2403;
  assign n2411 = ~n882 & n2410;
  assign n2412 = ~n878 & n2411;
  assign n2413 = ~n876 & n2412;
  assign n2414 = n873 & n2413;
  assign n2415 = ~n876 & ~n2403;
  assign n2416 = ~n878 & n2415;
  assign n2417 = ~n882 & n2416;
  assign n2418 = n885 & n2417;
  assign n2419 = ~n882 & ~n2403;
  assign n2420 = ~n878 & n2419;
  assign n2421 = n876 & n2420;
  assign n2422 = n882 & ~n2403;
  assign n2423 = ~n878 & n2422;
  assign n2424 = n878 & ~n2403;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~n2421 & n2425;
  assign n2427 = ~n2418 & n2426;
  assign n2428 = ~n2414 & n2427;
  assign n2429 = ~n2409 & n2428;
  assign \V197(13)  = n2392 | ~n2429;
  assign n2431 = \V116(12)  & ~\V133(10) ;
  assign n2432 = ~n885 & n2431;
  assign n2433 = ~n882 & n2432;
  assign n2434 = ~n878 & n2433;
  assign n2435 = ~n876 & n2434;
  assign n2436 = ~n873 & n2435;
  assign n2437 = \V133(9)  & n2436;
  assign n2438 = ~\V133(10)  & n2437;
  assign n2439 = \V47(29)  & n421;
  assign n2440 = n424 & n2439;
  assign n2441 = n434 & n2440;
  assign n2442 = ~n440 & n2441;
  assign n2443 = \V84(4)  & ~n434;
  assign n2444 = n424 & n2443;
  assign n2445 = \V84(12)  & ~n424;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n802 & n2446;
  assign n2448 = ~n2442 & n2447;
  assign n2449 = ~n443 & n2448;
  assign n2450 = ~n873 & ~n2449;
  assign n2451 = ~n876 & n2450;
  assign n2452 = ~n878 & n2451;
  assign n2453 = ~n882 & n2452;
  assign n2454 = ~n885 & n2453;
  assign n2455 = \V133(10)  & n2454;
  assign n2456 = ~n885 & ~n2449;
  assign n2457 = ~n882 & n2456;
  assign n2458 = ~n878 & n2457;
  assign n2459 = ~n876 & n2458;
  assign n2460 = n873 & n2459;
  assign n2461 = ~n876 & ~n2449;
  assign n2462 = ~n878 & n2461;
  assign n2463 = ~n882 & n2462;
  assign n2464 = n885 & n2463;
  assign n2465 = ~n882 & ~n2449;
  assign n2466 = ~n878 & n2465;
  assign n2467 = n876 & n2466;
  assign n2468 = n882 & ~n2449;
  assign n2469 = ~n878 & n2468;
  assign n2470 = n878 & ~n2449;
  assign n2471 = ~n2469 & ~n2470;
  assign n2472 = ~n2467 & n2471;
  assign n2473 = ~n2464 & n2472;
  assign n2474 = ~n2460 & n2473;
  assign n2475 = ~n2455 & n2474;
  assign \V197(12)  = n2438 | ~n2475;
  assign n2477 = n544 & ~n885;
  assign n2478 = ~n882 & n2477;
  assign n2479 = ~n878 & n2478;
  assign n2480 = ~n876 & n2479;
  assign n2481 = ~n873 & n2480;
  assign n2482 = \V133(9)  & n2481;
  assign n2483 = ~\V133(10)  & n2482;
  assign n2484 = \V84(0)  & n421;
  assign n2485 = n424 & n2484;
  assign n2486 = n434 & n2485;
  assign n2487 = ~n440 & n2486;
  assign n2488 = \V84(4)  & n434;
  assign n2489 = n424 & n2488;
  assign n2490 = ~n421 & n2489;
  assign n2491 = \V84(7)  & ~n434;
  assign n2492 = n424 & n2491;
  assign n2493 = \V84(15)  & ~n424;
  assign n2494 = ~n2492 & ~n2493;
  assign n2495 = ~n2490 & n2494;
  assign n2496 = ~n2487 & n2495;
  assign n2497 = ~n443 & n2496;
  assign n2498 = ~n873 & ~n2497;
  assign n2499 = ~n876 & n2498;
  assign n2500 = ~n878 & n2499;
  assign n2501 = ~n882 & n2500;
  assign n2502 = ~n885 & n2501;
  assign n2503 = \V133(10)  & n2502;
  assign n2504 = ~n885 & ~n2497;
  assign n2505 = ~n882 & n2504;
  assign n2506 = ~n878 & n2505;
  assign n2507 = ~n876 & n2506;
  assign n2508 = n873 & n2507;
  assign n2509 = ~n876 & ~n2497;
  assign n2510 = ~n878 & n2509;
  assign n2511 = ~n882 & n2510;
  assign n2512 = n885 & n2511;
  assign n2513 = ~n882 & ~n2497;
  assign n2514 = ~n878 & n2513;
  assign n2515 = n876 & n2514;
  assign n2516 = n882 & ~n2497;
  assign n2517 = ~n878 & n2516;
  assign n2518 = n878 & ~n2497;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = ~n2515 & n2519;
  assign n2521 = ~n2512 & n2520;
  assign n2522 = ~n2508 & n2521;
  assign n2523 = ~n2503 & n2522;
  assign \V197(15)  = n2483 | ~n2523;
  assign n2525 = n598 & ~n885;
  assign n2526 = ~n882 & n2525;
  assign n2527 = ~n878 & n2526;
  assign n2528 = ~n876 & n2527;
  assign n2529 = ~n873 & n2528;
  assign n2530 = \V133(9)  & n2529;
  assign n2531 = ~\V133(10)  & n2530;
  assign n2532 = \V47(31)  & n421;
  assign n2533 = n424 & n2532;
  assign n2534 = n434 & n2533;
  assign n2535 = ~n440 & n2534;
  assign n2536 = \V84(3)  & n434;
  assign n2537 = n424 & n2536;
  assign n2538 = ~n421 & n2537;
  assign n2539 = \V84(6)  & ~n434;
  assign n2540 = n424 & n2539;
  assign n2541 = \V84(14)  & ~n424;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = ~n2538 & n2542;
  assign n2544 = ~n2535 & n2543;
  assign n2545 = ~n443 & n2544;
  assign n2546 = ~n873 & ~n2545;
  assign n2547 = ~n876 & n2546;
  assign n2548 = ~n878 & n2547;
  assign n2549 = ~n882 & n2548;
  assign n2550 = ~n885 & n2549;
  assign n2551 = \V133(10)  & n2550;
  assign n2552 = ~n885 & ~n2545;
  assign n2553 = ~n882 & n2552;
  assign n2554 = ~n878 & n2553;
  assign n2555 = ~n876 & n2554;
  assign n2556 = n873 & n2555;
  assign n2557 = ~n876 & ~n2545;
  assign n2558 = ~n878 & n2557;
  assign n2559 = ~n882 & n2558;
  assign n2560 = n885 & n2559;
  assign n2561 = ~n882 & ~n2545;
  assign n2562 = ~n878 & n2561;
  assign n2563 = n876 & n2562;
  assign n2564 = n882 & ~n2545;
  assign n2565 = ~n878 & n2564;
  assign n2566 = n878 & ~n2545;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = ~n2563 & n2567;
  assign n2569 = ~n2560 & n2568;
  assign n2570 = ~n2556 & n2569;
  assign n2571 = ~n2551 & n2570;
  assign \V197(14)  = n2531 | ~n2571;
  assign n2573 = ~n468 & n1638;
  assign n2574 = ~n403 & n2573;
  assign n2575 = \V133(9)  & n2574;
  assign n2576 = ~\V133(10)  & n2575;
  assign n2577 = \V15(5)  & n421;
  assign n2578 = n424 & n2577;
  assign n2579 = n434 & n2578;
  assign n2580 = ~n440 & n2579;
  assign n2581 = \V47(6)  & ~n424;
  assign n2582 = ~n443 & ~n2581;
  assign n2583 = ~n2108 & n2582;
  assign n2584 = ~n2580 & n2583;
  assign n2585 = ~n403 & ~n2584;
  assign n2586 = ~n468 & n2585;
  assign n2587 = \V133(10)  & n2586;
  assign n2588 = n403 & ~n2584;
  assign n2589 = ~n468 & n2588;
  assign n2590 = n468 & ~n2584;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = ~n2587 & n2591;
  assign \V142(3)  = n2576 | ~n2592;
  assign n2594 = ~n468 & n1092;
  assign n2595 = ~n403 & n2594;
  assign n2596 = \V133(9)  & n2595;
  assign n2597 = ~\V133(10)  & n2596;
  assign n2598 = \V15(4)  & n421;
  assign n2599 = n424 & n2598;
  assign n2600 = n434 & n2599;
  assign n2601 = ~n440 & n2600;
  assign n2602 = \V47(5)  & ~n424;
  assign n2603 = ~n443 & ~n2602;
  assign n2604 = ~n2157 & n2603;
  assign n2605 = ~n2601 & n2604;
  assign n2606 = ~n403 & ~n2605;
  assign n2607 = ~n468 & n2606;
  assign n2608 = \V133(10)  & n2607;
  assign n2609 = n403 & ~n2605;
  assign n2610 = ~n468 & n2609;
  assign n2611 = n468 & ~n2605;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2608 & n2612;
  assign \V142(2)  = n2597 | ~n2613;
  assign n2615 = ~n468 & n1827;
  assign n2616 = ~n403 & n2615;
  assign n2617 = \V133(9)  & n2616;
  assign n2618 = ~\V133(10)  & n2617;
  assign n2619 = \V15(7)  & n421;
  assign n2620 = n424 & n2619;
  assign n2621 = n434 & n2620;
  assign n2622 = ~n440 & n2621;
  assign n2623 = \V47(0)  & ~n434;
  assign n2624 = n424 & n2623;
  assign n2625 = \V47(8)  & ~n424;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2206 & n2626;
  assign n2628 = ~n2622 & n2627;
  assign n2629 = ~n443 & n2628;
  assign n2630 = ~n403 & ~n2629;
  assign n2631 = ~n468 & n2630;
  assign n2632 = \V133(10)  & n2631;
  assign n2633 = n403 & ~n2629;
  assign n2634 = ~n468 & n2633;
  assign n2635 = n468 & ~n2629;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = ~n2632 & n2636;
  assign \V142(5)  = n2618 | ~n2637;
  assign n2639 = ~n468 & n1589;
  assign n2640 = ~n403 & n2639;
  assign n2641 = \V133(9)  & n2640;
  assign n2642 = ~\V133(10)  & n2641;
  assign n2643 = \V15(6)  & n421;
  assign n2644 = n424 & n2643;
  assign n2645 = n434 & n2644;
  assign n2646 = ~n440 & n2645;
  assign n2647 = \V47(7)  & ~n424;
  assign n2648 = ~n443 & ~n2647;
  assign n2649 = ~n2255 & n2648;
  assign n2650 = ~n2646 & n2649;
  assign n2651 = ~n403 & ~n2650;
  assign n2652 = ~n468 & n2651;
  assign n2653 = \V133(10)  & n2652;
  assign n2654 = n403 & ~n2650;
  assign n2655 = ~n468 & n2654;
  assign n2656 = n468 & ~n2650;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = ~n2653 & n2657;
  assign \V142(4)  = n2642 | ~n2658;
  assign n2660 = ~n885 & n1354;
  assign n2661 = ~n882 & n2660;
  assign n2662 = ~n878 & n2661;
  assign n2663 = ~n876 & n2662;
  assign n2664 = ~n873 & n2663;
  assign n2665 = \V133(9)  & n2664;
  assign n2666 = ~\V133(10)  & n2665;
  assign n2667 = \V84(16)  & n421;
  assign n2668 = n424 & n2667;
  assign n2669 = n434 & n2668;
  assign n2670 = ~n440 & n2669;
  assign n2671 = \V84(20)  & n434;
  assign n2672 = n424 & n2671;
  assign n2673 = ~n421 & n2672;
  assign n2674 = \V84(23)  & ~n434;
  assign n2675 = n424 & n2674;
  assign n2676 = \V84(31)  & ~n424;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = ~n2673 & n2677;
  assign n2679 = ~n2670 & n2678;
  assign n2680 = ~n443 & n2679;
  assign n2681 = ~n873 & ~n2680;
  assign n2682 = ~n876 & n2681;
  assign n2683 = ~n878 & n2682;
  assign n2684 = ~n882 & n2683;
  assign n2685 = ~n885 & n2684;
  assign n2686 = \V133(10)  & n2685;
  assign n2687 = ~n885 & ~n2680;
  assign n2688 = ~n882 & n2687;
  assign n2689 = ~n878 & n2688;
  assign n2690 = ~n876 & n2689;
  assign n2691 = n873 & n2690;
  assign n2692 = ~n876 & ~n2680;
  assign n2693 = ~n878 & n2692;
  assign n2694 = ~n882 & n2693;
  assign n2695 = n885 & n2694;
  assign n2696 = ~n882 & ~n2680;
  assign n2697 = ~n878 & n2696;
  assign n2698 = n876 & n2697;
  assign n2699 = n882 & ~n2680;
  assign n2700 = ~n878 & n2699;
  assign n2701 = n878 & ~n2680;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = ~n2698 & n2702;
  assign n2704 = ~n2695 & n2703;
  assign n2705 = ~n2691 & n2704;
  assign n2706 = ~n2686 & n2705;
  assign \V197(31)  = n2666 | ~n2706;
  assign n2708 = ~n468 & n1195;
  assign n2709 = ~n403 & n2708;
  assign n2710 = \V133(9)  & n2709;
  assign n2711 = ~\V133(10)  & n2710;
  assign n2712 = \V15(3)  & n421;
  assign n2713 = n424 & n2712;
  assign n2714 = n434 & n2713;
  assign n2715 = ~n440 & n2714;
  assign n2716 = \V47(4)  & ~n424;
  assign n2717 = ~n443 & ~n2716;
  assign n2718 = ~n2490 & n2717;
  assign n2719 = ~n2715 & n2718;
  assign n2720 = ~n403 & ~n2719;
  assign n2721 = ~n468 & n2720;
  assign n2722 = \V133(10)  & n2721;
  assign n2723 = n403 & ~n2719;
  assign n2724 = ~n468 & n2723;
  assign n2725 = n468 & ~n2719;
  assign n2726 = ~n2724 & ~n2725;
  assign n2727 = ~n2722 & n2726;
  assign \V142(1)  = n2711 | ~n2727;
  assign n2729 = ~n885 & n1051;
  assign n2730 = ~n882 & n2729;
  assign n2731 = ~n878 & n2730;
  assign n2732 = ~n876 & n2731;
  assign n2733 = ~n873 & n2732;
  assign n2734 = \V133(9)  & n2733;
  assign n2735 = ~\V133(10)  & n2734;
  assign n2736 = \V84(15)  & n421;
  assign n2737 = n424 & n2736;
  assign n2738 = n434 & n2737;
  assign n2739 = ~n440 & n2738;
  assign n2740 = \V84(19)  & n434;
  assign n2741 = n424 & n2740;
  assign n2742 = ~n421 & n2741;
  assign n2743 = \V84(22)  & ~n434;
  assign n2744 = n424 & n2743;
  assign n2745 = \V84(30)  & ~n424;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = ~n2742 & n2746;
  assign n2748 = ~n2739 & n2747;
  assign n2749 = ~n443 & n2748;
  assign n2750 = ~n873 & ~n2749;
  assign n2751 = ~n876 & n2750;
  assign n2752 = ~n878 & n2751;
  assign n2753 = ~n882 & n2752;
  assign n2754 = ~n885 & n2753;
  assign n2755 = \V133(10)  & n2754;
  assign n2756 = ~n885 & ~n2749;
  assign n2757 = ~n882 & n2756;
  assign n2758 = ~n878 & n2757;
  assign n2759 = ~n876 & n2758;
  assign n2760 = n873 & n2759;
  assign n2761 = ~n876 & ~n2749;
  assign n2762 = ~n878 & n2761;
  assign n2763 = ~n882 & n2762;
  assign n2764 = n885 & n2763;
  assign n2765 = ~n882 & ~n2749;
  assign n2766 = ~n878 & n2765;
  assign n2767 = n876 & n2766;
  assign n2768 = n882 & ~n2749;
  assign n2769 = ~n878 & n2768;
  assign n2770 = n878 & ~n2749;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = ~n2767 & n2771;
  assign n2773 = ~n2764 & n2772;
  assign n2774 = ~n2760 & n2773;
  assign n2775 = ~n2755 & n2774;
  assign \V197(30)  = n2735 | ~n2775;
  assign n2777 = ~n468 & n886;
  assign n2778 = ~n403 & n2777;
  assign n2779 = \V133(9)  & n2778;
  assign n2780 = ~\V133(10)  & n2779;
  assign n2781 = \V15(2)  & n421;
  assign n2782 = n424 & n2781;
  assign n2783 = n434 & n2782;
  assign n2784 = ~n440 & n2783;
  assign n2785 = \V47(3)  & ~n424;
  assign n2786 = ~n443 & ~n2785;
  assign n2787 = ~n2538 & n2786;
  assign n2788 = ~n2784 & n2787;
  assign n2789 = ~n403 & ~n2788;
  assign n2790 = ~n468 & n2789;
  assign n2791 = \V133(10)  & n2790;
  assign n2792 = n403 & ~n2788;
  assign n2793 = ~n468 & n2792;
  assign n2794 = n468 & ~n2788;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2791 & n2795;
  assign \V142(0)  = n2780 | ~n2796;
  assign n2798 = \V84(20)  & ~n530;
  assign n2799 = ~n403 & n2798;
  assign n2800 = ~n529 & n2799;
  assign n2801 = ~n527 & n2800;
  assign n2802 = ~n525 & n2801;
  assign n2803 = ~\V133(10)  & n2802;
  assign n2804 = ~\V133(7)  & n2803;
  assign n2805 = ~\V133(9)  & n2804;
  assign n2806 = ~\V133(4)  & n2805;
  assign n2807 = ~\V133(3)  & n2806;
  assign n2808 = \V133(2)  & n2807;
  assign n2809 = \V133(1)  & n2808;
  assign n2810 = ~\V133(10)  & n2809;
  assign n2811 = ~n525 & n1781;
  assign n2812 = ~n527 & n2811;
  assign n2813 = ~n529 & n2812;
  assign n2814 = ~n403 & n2813;
  assign n2815 = n530 & n2814;
  assign n2816 = \V47(5)  & n421;
  assign n2817 = n424 & n2816;
  assign n2818 = n434 & n2817;
  assign n2819 = ~n440 & n2818;
  assign n2820 = \V47(9)  & n434;
  assign n2821 = n424 & n2820;
  assign n2822 = ~n421 & n2821;
  assign n2823 = \V47(12)  & ~n434;
  assign n2824 = n424 & n2823;
  assign n2825 = \V47(20)  & ~n424;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = ~n2822 & n2826;
  assign n2828 = ~n2819 & n2827;
  assign n2829 = ~n443 & n2828;
  assign n2830 = ~n403 & ~n2829;
  assign n2831 = ~n529 & n2830;
  assign n2832 = ~n527 & n2831;
  assign n2833 = ~n525 & n2832;
  assign n2834 = \V133(10)  & n2833;
  assign n2835 = ~n525 & ~n2829;
  assign n2836 = ~n527 & n2835;
  assign n2837 = ~n529 & n2836;
  assign n2838 = n403 & n2837;
  assign n2839 = ~n529 & ~n2829;
  assign n2840 = ~n527 & n2839;
  assign n2841 = n525 & n2840;
  assign n2842 = n529 & ~n2829;
  assign n2843 = ~n527 & n2842;
  assign n2844 = n527 & ~n2829;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = ~n2841 & n2845;
  assign n2847 = ~n2838 & n2846;
  assign n2848 = ~n2834 & n2847;
  assign n2849 = ~n2815 & n2848;
  assign \V165(3)  = n2810 | ~n2849;
  assign n2851 = \V116(11)  & ~n227;
  assign n2852 = ~n220 & n2851;
  assign n2853 = ~n219 & n2852;
  assign n2854 = ~\V133(10)  & n2853;
  assign n2855 = \V133(9)  & n2854;
  assign n2856 = ~\V133(10)  & n2855;
  assign n2857 = \V84(28)  & ~n220;
  assign n2858 = ~n219 & n2857;
  assign n2859 = \V133(10)  & n2858;
  assign n2860 = \V84(28)  & n220;
  assign n2861 = ~n219 & n2860;
  assign n2862 = \V84(28)  & n219;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = ~n2859 & n2863;
  assign n2865 = ~n236 & n2864;
  assign \V212(11)  = n2856 | ~n2865;
  assign n2867 = \V84(19)  & ~n530;
  assign n2868 = ~n403 & n2867;
  assign n2869 = ~n529 & n2868;
  assign n2870 = ~n527 & n2869;
  assign n2871 = ~n525 & n2870;
  assign n2872 = ~\V133(10)  & n2871;
  assign n2873 = ~\V133(7)  & n2872;
  assign n2874 = ~\V133(9)  & n2873;
  assign n2875 = ~\V133(4)  & n2874;
  assign n2876 = ~\V133(3)  & n2875;
  assign n2877 = \V133(2)  & n2876;
  assign n2878 = \V133(1)  & n2877;
  assign n2879 = ~\V133(10)  & n2878;
  assign n2880 = ~n525 & n2192;
  assign n2881 = ~n527 & n2880;
  assign n2882 = ~n529 & n2881;
  assign n2883 = ~n403 & n2882;
  assign n2884 = n530 & n2883;
  assign n2885 = \V47(4)  & n421;
  assign n2886 = n424 & n2885;
  assign n2887 = n434 & n2886;
  assign n2888 = ~n440 & n2887;
  assign n2889 = \V47(8)  & n434;
  assign n2890 = n424 & n2889;
  assign n2891 = ~n421 & n2890;
  assign n2892 = \V47(11)  & ~n434;
  assign n2893 = n424 & n2892;
  assign n2894 = \V47(19)  & ~n424;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = ~n2891 & n2895;
  assign n2897 = ~n2888 & n2896;
  assign n2898 = ~n443 & n2897;
  assign n2899 = ~n403 & ~n2898;
  assign n2900 = ~n529 & n2899;
  assign n2901 = ~n527 & n2900;
  assign n2902 = ~n525 & n2901;
  assign n2903 = \V133(10)  & n2902;
  assign n2904 = ~n525 & ~n2898;
  assign n2905 = ~n527 & n2904;
  assign n2906 = ~n529 & n2905;
  assign n2907 = n403 & n2906;
  assign n2908 = ~n529 & ~n2898;
  assign n2909 = ~n527 & n2908;
  assign n2910 = n525 & n2909;
  assign n2911 = n529 & ~n2898;
  assign n2912 = ~n527 & n2911;
  assign n2913 = n527 & ~n2898;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = ~n2910 & n2914;
  assign n2916 = ~n2907 & n2915;
  assign n2917 = ~n2903 & n2916;
  assign n2918 = ~n2884 & n2917;
  assign \V165(2)  = n2879 | ~n2918;
  assign n2920 = \V116(10)  & ~n227;
  assign n2921 = ~n220 & n2920;
  assign n2922 = ~n219 & n2921;
  assign n2923 = ~\V133(10)  & n2922;
  assign n2924 = \V133(9)  & n2923;
  assign n2925 = ~\V133(10)  & n2924;
  assign n2926 = \V84(27)  & ~n220;
  assign n2927 = ~n219 & n2926;
  assign n2928 = \V133(10)  & n2927;
  assign n2929 = \V84(27)  & n220;
  assign n2930 = ~n219 & n2929;
  assign n2931 = \V84(27)  & n219;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = ~n2928 & n2932;
  assign n2934 = ~n236 & n2933;
  assign \V212(10)  = n2925 | ~n2934;
  assign n2936 = \V84(22)  & ~n530;
  assign n2937 = ~n403 & n2936;
  assign n2938 = ~n529 & n2937;
  assign n2939 = ~n527 & n2938;
  assign n2940 = ~n525 & n2939;
  assign n2941 = ~\V133(10)  & n2940;
  assign n2942 = ~\V133(7)  & n2941;
  assign n2943 = ~\V133(9)  & n2942;
  assign n2944 = ~\V133(4)  & n2943;
  assign n2945 = ~\V133(3)  & n2944;
  assign n2946 = \V133(2)  & n2945;
  assign n2947 = \V133(1)  & n2946;
  assign n2948 = ~\V133(10)  & n2947;
  assign n2949 = ~n525 & n1925;
  assign n2950 = ~n527 & n2949;
  assign n2951 = ~n529 & n2950;
  assign n2952 = ~n403 & n2951;
  assign n2953 = n530 & n2952;
  assign n2954 = \V47(7)  & n421;
  assign n2955 = n424 & n2954;
  assign n2956 = n434 & n2955;
  assign n2957 = ~n440 & n2956;
  assign n2958 = \V47(11)  & n434;
  assign n2959 = n424 & n2958;
  assign n2960 = ~n421 & n2959;
  assign n2961 = \V47(14)  & ~n434;
  assign n2962 = n424 & n2961;
  assign n2963 = \V47(22)  & ~n424;
  assign n2964 = ~n2962 & ~n2963;
  assign n2965 = ~n2960 & n2964;
  assign n2966 = ~n2957 & n2965;
  assign n2967 = ~n443 & n2966;
  assign n2968 = ~n403 & ~n2967;
  assign n2969 = ~n529 & n2968;
  assign n2970 = ~n527 & n2969;
  assign n2971 = ~n525 & n2970;
  assign n2972 = \V133(10)  & n2971;
  assign n2973 = ~n525 & ~n2967;
  assign n2974 = ~n527 & n2973;
  assign n2975 = ~n529 & n2974;
  assign n2976 = n403 & n2975;
  assign n2977 = ~n529 & ~n2967;
  assign n2978 = ~n527 & n2977;
  assign n2979 = n525 & n2978;
  assign n2980 = n529 & ~n2967;
  assign n2981 = ~n527 & n2980;
  assign n2982 = n527 & ~n2967;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2979 & n2983;
  assign n2985 = ~n2976 & n2984;
  assign n2986 = ~n2972 & n2985;
  assign n2987 = ~n2953 & n2986;
  assign \V165(5)  = n2948 | ~n2987;
  assign n2989 = \V116(13)  & ~n227;
  assign n2990 = ~n220 & n2989;
  assign n2991 = ~n219 & n2990;
  assign n2992 = ~\V133(10)  & n2991;
  assign n2993 = \V133(9)  & n2992;
  assign n2994 = ~\V133(10)  & n2993;
  assign n2995 = \V84(30)  & ~n220;
  assign n2996 = ~n219 & n2995;
  assign n2997 = \V133(10)  & n2996;
  assign n2998 = \V84(30)  & n220;
  assign n2999 = ~n219 & n2998;
  assign n3000 = \V84(30)  & n219;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = ~n2997 & n3001;
  assign n3003 = ~n236 & n3002;
  assign \V212(13)  = n2994 | ~n3003;
  assign n3005 = \V84(21)  & ~n530;
  assign n3006 = ~n403 & n3005;
  assign n3007 = ~n529 & n3006;
  assign n3008 = ~n527 & n3007;
  assign n3009 = ~n525 & n3008;
  assign n3010 = ~\V133(10)  & n3009;
  assign n3011 = ~\V133(7)  & n3010;
  assign n3012 = ~\V133(9)  & n3011;
  assign n3013 = ~\V133(4)  & n3012;
  assign n3014 = ~\V133(3)  & n3013;
  assign n3015 = \V133(2)  & n3014;
  assign n3016 = \V133(1)  & n3015;
  assign n3017 = ~\V133(10)  & n3016;
  assign n3018 = ~n525 & n1687;
  assign n3019 = ~n527 & n3018;
  assign n3020 = ~n529 & n3019;
  assign n3021 = ~n403 & n3020;
  assign n3022 = n530 & n3021;
  assign n3023 = \V47(6)  & n421;
  assign n3024 = n424 & n3023;
  assign n3025 = n434 & n3024;
  assign n3026 = ~n440 & n3025;
  assign n3027 = \V47(10)  & n434;
  assign n3028 = n424 & n3027;
  assign n3029 = ~n421 & n3028;
  assign n3030 = \V47(13)  & ~n434;
  assign n3031 = n424 & n3030;
  assign n3032 = \V47(21)  & ~n424;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = ~n3029 & n3033;
  assign n3035 = ~n3026 & n3034;
  assign n3036 = ~n443 & n3035;
  assign n3037 = ~n403 & ~n3036;
  assign n3038 = ~n529 & n3037;
  assign n3039 = ~n527 & n3038;
  assign n3040 = ~n525 & n3039;
  assign n3041 = \V133(10)  & n3040;
  assign n3042 = ~n525 & ~n3036;
  assign n3043 = ~n527 & n3042;
  assign n3044 = ~n529 & n3043;
  assign n3045 = n403 & n3044;
  assign n3046 = ~n529 & ~n3036;
  assign n3047 = ~n527 & n3046;
  assign n3048 = n525 & n3047;
  assign n3049 = n529 & ~n3036;
  assign n3050 = ~n527 & n3049;
  assign n3051 = n527 & ~n3036;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = ~n3048 & n3052;
  assign n3054 = ~n3045 & n3053;
  assign n3055 = ~n3041 & n3054;
  assign n3056 = ~n3022 & n3055;
  assign \V165(4)  = n3017 | ~n3056;
  assign n3058 = \V116(12)  & ~n227;
  assign n3059 = ~n220 & n3058;
  assign n3060 = ~n219 & n3059;
  assign n3061 = ~\V133(10)  & n3060;
  assign n3062 = \V133(9)  & n3061;
  assign n3063 = ~\V133(10)  & n3062;
  assign n3064 = \V84(29)  & ~n220;
  assign n3065 = ~n219 & n3064;
  assign n3066 = \V133(10)  & n3065;
  assign n3067 = \V84(29)  & n220;
  assign n3068 = ~n219 & n3067;
  assign n3069 = \V84(29)  & n219;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3066 & n3070;
  assign n3072 = ~n236 & n3071;
  assign \V212(12)  = n3063 | ~n3072;
  assign n3074 = ~\V133(4)  & n215;
  assign n3075 = \V84(12)  & ~n530;
  assign n3076 = ~n403 & n3075;
  assign n3077 = ~n529 & n3076;
  assign n3078 = ~n3074 & n3077;
  assign n3079 = ~n525 & n3078;
  assign n3080 = ~\V133(10)  & n3079;
  assign n3081 = ~\V133(7)  & n3080;
  assign n3082 = ~\V133(9)  & n3081;
  assign n3083 = ~\V133(4)  & n3082;
  assign n3084 = ~\V133(3)  & n3083;
  assign n3085 = \V133(2)  & n3084;
  assign n3086 = \V133(1)  & n3085;
  assign n3087 = ~\V133(10)  & n3086;
  assign n3088 = ~n525 & n2431;
  assign n3089 = ~n3074 & n3088;
  assign n3090 = ~n529 & n3089;
  assign n3091 = ~n403 & n3090;
  assign n3092 = n530 & n3091;
  assign n3093 = \V15(11)  & n421;
  assign n3094 = n424 & n3093;
  assign n3095 = n434 & n3094;
  assign n3096 = ~n440 & n3095;
  assign n3097 = \V47(1)  & n434;
  assign n3098 = n424 & n3097;
  assign n3099 = ~n421 & n3098;
  assign n3100 = \V47(4)  & ~n434;
  assign n3101 = n424 & n3100;
  assign n3102 = \V47(12)  & ~n424;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n3099 & n3103;
  assign n3105 = ~n3096 & n3104;
  assign n3106 = ~n443 & n3105;
  assign n3107 = ~n403 & ~n3106;
  assign n3108 = ~n529 & n3107;
  assign n3109 = ~n3074 & n3108;
  assign n3110 = ~n525 & n3109;
  assign n3111 = \V133(10)  & n3110;
  assign n3112 = ~n525 & ~n3106;
  assign n3113 = ~n3074 & n3112;
  assign n3114 = ~n529 & n3113;
  assign n3115 = n403 & n3114;
  assign n3116 = ~n529 & ~n3106;
  assign n3117 = ~n3074 & n3116;
  assign n3118 = n525 & n3117;
  assign n3119 = n529 & ~n3106;
  assign n3120 = ~n3074 & n3119;
  assign n3121 = n3074 & ~n3106;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = ~n3118 & n3122;
  assign n3124 = ~n3115 & n3123;
  assign n3125 = ~n3111 & n3124;
  assign n3126 = ~n3092 & n3125;
  assign \V146(0)  = n3087 | ~n3126;
  assign n3128 = \V116(14)  & ~n227;
  assign n3129 = ~n220 & n3128;
  assign n3130 = ~n219 & n3129;
  assign n3131 = ~\V133(10)  & n3130;
  assign n3132 = \V133(9)  & n3131;
  assign n3133 = ~\V133(10)  & n3132;
  assign n3134 = \V84(31)  & ~n220;
  assign n3135 = ~n219 & n3134;
  assign n3136 = \V133(10)  & n3135;
  assign n3137 = \V84(31)  & n220;
  assign n3138 = ~n219 & n3137;
  assign n3139 = \V84(31)  & n219;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~n3136 & n3140;
  assign n3142 = ~n236 & n3141;
  assign \V212(14)  = n3133 | ~n3142;
  assign n3144 = \V84(18)  & ~n530;
  assign n3145 = ~n403 & n3144;
  assign n3146 = ~n529 & n3145;
  assign n3147 = ~n527 & n3146;
  assign n3148 = ~n525 & n3147;
  assign n3149 = ~\V133(10)  & n3148;
  assign n3150 = ~\V133(7)  & n3149;
  assign n3151 = ~\V133(9)  & n3150;
  assign n3152 = ~\V133(4)  & n3151;
  assign n3153 = ~\V133(3)  & n3152;
  assign n3154 = \V133(2)  & n3153;
  assign n3155 = \V133(1)  & n3154;
  assign n3156 = ~\V133(10)  & n3155;
  assign n3157 = ~n525 & n2241;
  assign n3158 = ~n527 & n3157;
  assign n3159 = ~n529 & n3158;
  assign n3160 = ~n403 & n3159;
  assign n3161 = n530 & n3160;
  assign n3162 = \V47(3)  & n421;
  assign n3163 = n424 & n3162;
  assign n3164 = n434 & n3163;
  assign n3165 = ~n440 & n3164;
  assign n3166 = \V47(7)  & n434;
  assign n3167 = n424 & n3166;
  assign n3168 = ~n421 & n3167;
  assign n3169 = \V47(10)  & ~n434;
  assign n3170 = n424 & n3169;
  assign n3171 = \V47(18)  & ~n424;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = ~n3168 & n3172;
  assign n3174 = ~n3165 & n3173;
  assign n3175 = ~n443 & n3174;
  assign n3176 = ~n403 & ~n3175;
  assign n3177 = ~n529 & n3176;
  assign n3178 = ~n527 & n3177;
  assign n3179 = ~n525 & n3178;
  assign n3180 = \V133(10)  & n3179;
  assign n3181 = ~n525 & ~n3175;
  assign n3182 = ~n527 & n3181;
  assign n3183 = ~n529 & n3182;
  assign n3184 = n403 & n3183;
  assign n3185 = ~n529 & ~n3175;
  assign n3186 = ~n527 & n3185;
  assign n3187 = n525 & n3186;
  assign n3188 = n529 & ~n3175;
  assign n3189 = ~n527 & n3188;
  assign n3190 = n527 & ~n3175;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = ~n3187 & n3191;
  assign n3193 = ~n3184 & n3192;
  assign n3194 = ~n3180 & n3193;
  assign n3195 = ~n3161 & n3194;
  assign \V165(1)  = n3156 | ~n3195;
  assign n3197 = \V84(17)  & ~n530;
  assign n3198 = ~n403 & n3197;
  assign n3199 = ~n529 & n3198;
  assign n3200 = ~n527 & n3199;
  assign n3201 = ~n525 & n3200;
  assign n3202 = ~\V133(10)  & n3201;
  assign n3203 = ~\V133(7)  & n3202;
  assign n3204 = ~\V133(9)  & n3203;
  assign n3205 = ~\V133(4)  & n3204;
  assign n3206 = ~\V133(3)  & n3205;
  assign n3207 = \V133(2)  & n3206;
  assign n3208 = \V133(1)  & n3207;
  assign n3209 = ~\V133(10)  & n3208;
  assign n3210 = ~n525 & n2094;
  assign n3211 = ~n527 & n3210;
  assign n3212 = ~n529 & n3211;
  assign n3213 = ~n403 & n3212;
  assign n3214 = n530 & n3213;
  assign n3215 = \V47(2)  & n421;
  assign n3216 = n424 & n3215;
  assign n3217 = n434 & n3216;
  assign n3218 = ~n440 & n3217;
  assign n3219 = \V47(6)  & n434;
  assign n3220 = n424 & n3219;
  assign n3221 = ~n421 & n3220;
  assign n3222 = \V47(9)  & ~n434;
  assign n3223 = n424 & n3222;
  assign n3224 = \V47(17)  & ~n424;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = ~n3221 & n3225;
  assign n3227 = ~n3218 & n3226;
  assign n3228 = ~n443 & n3227;
  assign n3229 = ~n403 & ~n3228;
  assign n3230 = ~n529 & n3229;
  assign n3231 = ~n527 & n3230;
  assign n3232 = ~n525 & n3231;
  assign n3233 = \V133(10)  & n3232;
  assign n3234 = ~n525 & ~n3228;
  assign n3235 = ~n527 & n3234;
  assign n3236 = ~n529 & n3235;
  assign n3237 = n403 & n3236;
  assign n3238 = ~n529 & ~n3228;
  assign n3239 = ~n527 & n3238;
  assign n3240 = n525 & n3239;
  assign n3241 = n529 & ~n3228;
  assign n3242 = ~n527 & n3241;
  assign n3243 = n527 & ~n3228;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = ~n3240 & n3244;
  assign n3246 = ~n3237 & n3245;
  assign n3247 = ~n3233 & n3246;
  assign n3248 = ~n3214 & n3247;
  assign \V165(0)  = n3209 | ~n3248;
  assign n3250 = \V84(24)  & ~n530;
  assign n3251 = ~n403 & n3250;
  assign n3252 = ~n529 & n3251;
  assign n3253 = ~n527 & n3252;
  assign n3254 = ~n525 & n3253;
  assign n3255 = ~\V133(10)  & n3254;
  assign n3256 = ~\V133(7)  & n3255;
  assign n3257 = ~\V133(9)  & n3256;
  assign n3258 = ~\V133(4)  & n3257;
  assign n3259 = ~\V133(3)  & n3258;
  assign n3260 = \V133(2)  & n3259;
  assign n3261 = \V133(1)  & n3260;
  assign n3262 = ~\V133(10)  & n3261;
  assign n3263 = ~n525 & n2020;
  assign n3264 = ~n527 & n3263;
  assign n3265 = ~n529 & n3264;
  assign n3266 = ~n403 & n3265;
  assign n3267 = n530 & n3266;
  assign n3268 = \V47(9)  & n421;
  assign n3269 = n424 & n3268;
  assign n3270 = n434 & n3269;
  assign n3271 = ~n440 & n3270;
  assign n3272 = \V47(13)  & n434;
  assign n3273 = n424 & n3272;
  assign n3274 = ~n421 & n3273;
  assign n3275 = \V47(16)  & ~n434;
  assign n3276 = n424 & n3275;
  assign n3277 = \V47(24)  & ~n424;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n3274 & n3278;
  assign n3280 = ~n3271 & n3279;
  assign n3281 = ~n443 & n3280;
  assign n3282 = ~n403 & ~n3281;
  assign n3283 = ~n529 & n3282;
  assign n3284 = ~n527 & n3283;
  assign n3285 = ~n525 & n3284;
  assign n3286 = \V133(10)  & n3285;
  assign n3287 = ~n525 & ~n3281;
  assign n3288 = ~n527 & n3287;
  assign n3289 = ~n529 & n3288;
  assign n3290 = n403 & n3289;
  assign n3291 = ~n529 & ~n3281;
  assign n3292 = ~n527 & n3291;
  assign n3293 = n525 & n3292;
  assign n3294 = n529 & ~n3281;
  assign n3295 = ~n527 & n3294;
  assign n3296 = n527 & ~n3281;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n3293 & n3297;
  assign n3299 = ~n3290 & n3298;
  assign n3300 = ~n3286 & n3299;
  assign n3301 = ~n3267 & n3300;
  assign \V165(7)  = n3262 | ~n3301;
  assign n3303 = \V84(23)  & ~n530;
  assign n3304 = ~n403 & n3303;
  assign n3305 = ~n529 & n3304;
  assign n3306 = ~n527 & n3305;
  assign n3307 = ~n525 & n3306;
  assign n3308 = ~\V133(10)  & n3307;
  assign n3309 = ~\V133(7)  & n3308;
  assign n3310 = ~\V133(9)  & n3309;
  assign n3311 = ~\V133(4)  & n3310;
  assign n3312 = ~\V133(3)  & n3311;
  assign n3313 = \V133(2)  & n3312;
  assign n3314 = \V133(1)  & n3313;
  assign n3315 = ~\V133(10)  & n3314;
  assign n3316 = ~n525 & n1876;
  assign n3317 = ~n527 & n3316;
  assign n3318 = ~n529 & n3317;
  assign n3319 = ~n403 & n3318;
  assign n3320 = n530 & n3319;
  assign n3321 = \V47(8)  & n421;
  assign n3322 = n424 & n3321;
  assign n3323 = n434 & n3322;
  assign n3324 = ~n440 & n3323;
  assign n3325 = \V47(12)  & n434;
  assign n3326 = n424 & n3325;
  assign n3327 = ~n421 & n3326;
  assign n3328 = \V47(15)  & ~n434;
  assign n3329 = n424 & n3328;
  assign n3330 = \V47(23)  & ~n424;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = ~n3327 & n3331;
  assign n3333 = ~n3324 & n3332;
  assign n3334 = ~n443 & n3333;
  assign n3335 = ~n403 & ~n3334;
  assign n3336 = ~n529 & n3335;
  assign n3337 = ~n527 & n3336;
  assign n3338 = ~n525 & n3337;
  assign n3339 = \V133(10)  & n3338;
  assign n3340 = ~n525 & ~n3334;
  assign n3341 = ~n527 & n3340;
  assign n3342 = ~n529 & n3341;
  assign n3343 = n403 & n3342;
  assign n3344 = ~n529 & ~n3334;
  assign n3345 = ~n527 & n3344;
  assign n3346 = n525 & n3345;
  assign n3347 = n529 & ~n3334;
  assign n3348 = ~n527 & n3347;
  assign n3349 = n527 & ~n3334;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = ~n3346 & n3350;
  assign n3352 = ~n3343 & n3351;
  assign n3353 = ~n3339 & n3352;
  assign n3354 = ~n3320 & n3353;
  assign \V165(6)  = n3315 | ~n3354;
  assign n3356 = \V84(26)  & ~n530;
  assign n3357 = ~n403 & n3356;
  assign n3358 = ~n529 & n3357;
  assign n3359 = ~n527 & n3358;
  assign n3360 = ~n525 & n3359;
  assign n3361 = ~\V133(10)  & n3360;
  assign n3362 = ~\V133(7)  & n3361;
  assign n3363 = ~\V133(9)  & n3362;
  assign n3364 = ~\V133(4)  & n3363;
  assign n3365 = ~\V133(3)  & n3364;
  assign n3366 = \V133(2)  & n3365;
  assign n3367 = \V133(1)  & n3366;
  assign n3368 = ~\V133(10)  & n3367;
  assign n3369 = ~n525 & n1292;
  assign n3370 = ~n527 & n3369;
  assign n3371 = ~n529 & n3370;
  assign n3372 = ~n403 & n3371;
  assign n3373 = n530 & n3372;
  assign n3374 = \V47(11)  & n421;
  assign n3375 = n424 & n3374;
  assign n3376 = n434 & n3375;
  assign n3377 = ~n440 & n3376;
  assign n3378 = \V47(15)  & n434;
  assign n3379 = n424 & n3378;
  assign n3380 = ~n421 & n3379;
  assign n3381 = \V47(18)  & ~n434;
  assign n3382 = n424 & n3381;
  assign n3383 = \V47(26)  & ~n424;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = ~n3380 & n3384;
  assign n3386 = ~n3377 & n3385;
  assign n3387 = ~n443 & n3386;
  assign n3388 = ~n403 & ~n3387;
  assign n3389 = ~n529 & n3388;
  assign n3390 = ~n527 & n3389;
  assign n3391 = ~n525 & n3390;
  assign n3392 = \V133(10)  & n3391;
  assign n3393 = ~n525 & ~n3387;
  assign n3394 = ~n527 & n3393;
  assign n3395 = ~n529 & n3394;
  assign n3396 = n403 & n3395;
  assign n3397 = ~n529 & ~n3387;
  assign n3398 = ~n527 & n3397;
  assign n3399 = n525 & n3398;
  assign n3400 = n529 & ~n3387;
  assign n3401 = ~n527 & n3400;
  assign n3402 = n527 & ~n3387;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = ~n3399 & n3403;
  assign n3405 = ~n3396 & n3404;
  assign n3406 = ~n3392 & n3405;
  assign n3407 = ~n3373 & n3406;
  assign \V165(9)  = n3368 | ~n3407;
  assign n3409 = \V84(25)  & ~n530;
  assign n3410 = ~n403 & n3409;
  assign n3411 = ~n529 & n3410;
  assign n3412 = ~n527 & n3411;
  assign n3413 = ~n525 & n3412;
  assign n3414 = ~\V133(10)  & n3413;
  assign n3415 = ~\V133(7)  & n3414;
  assign n3416 = ~\V133(9)  & n3415;
  assign n3417 = ~\V133(4)  & n3416;
  assign n3418 = ~\V133(3)  & n3417;
  assign n3419 = \V133(2)  & n3418;
  assign n3420 = \V133(1)  & n3419;
  assign n3421 = ~\V133(10)  & n3420;
  assign n3422 = ~n525 & n1971;
  assign n3423 = ~n527 & n3422;
  assign n3424 = ~n529 & n3423;
  assign n3425 = ~n403 & n3424;
  assign n3426 = n530 & n3425;
  assign n3427 = \V47(10)  & n421;
  assign n3428 = n424 & n3427;
  assign n3429 = n434 & n3428;
  assign n3430 = ~n440 & n3429;
  assign n3431 = \V47(14)  & n434;
  assign n3432 = n424 & n3431;
  assign n3433 = ~n421 & n3432;
  assign n3434 = \V47(17)  & ~n434;
  assign n3435 = n424 & n3434;
  assign n3436 = \V47(25)  & ~n424;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = ~n3433 & n3437;
  assign n3439 = ~n3430 & n3438;
  assign n3440 = ~n443 & n3439;
  assign n3441 = ~n403 & ~n3440;
  assign n3442 = ~n529 & n3441;
  assign n3443 = ~n527 & n3442;
  assign n3444 = ~n525 & n3443;
  assign n3445 = \V133(10)  & n3444;
  assign n3446 = ~n525 & ~n3440;
  assign n3447 = ~n527 & n3446;
  assign n3448 = ~n529 & n3447;
  assign n3449 = n403 & n3448;
  assign n3450 = ~n529 & ~n3440;
  assign n3451 = ~n527 & n3450;
  assign n3452 = n525 & n3451;
  assign n3453 = n529 & ~n3440;
  assign n3454 = ~n527 & n3453;
  assign n3455 = n527 & ~n3440;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = ~n3452 & n3456;
  assign n3458 = ~n3449 & n3457;
  assign n3459 = ~n3445 & n3458;
  assign n3460 = ~n3426 & n3459;
  assign \V165(8)  = n3421 | ~n3460;
  assign n3462 = ~\V133(4)  & n216;
  assign n3463 = \V84(16)  & ~n530;
  assign n3464 = ~n403 & n3463;
  assign n3465 = ~n529 & n3464;
  assign n3466 = ~n3462 & n3465;
  assign n3467 = ~n527 & n3466;
  assign n3468 = ~n525 & n3467;
  assign n3469 = ~\V133(10)  & n3468;
  assign n3470 = ~\V133(7)  & n3469;
  assign n3471 = ~\V133(9)  & n3470;
  assign n3472 = ~\V133(4)  & n3471;
  assign n3473 = ~\V133(3)  & n3472;
  assign n3474 = \V133(2)  & n3473;
  assign n3475 = \V133(1)  & n3474;
  assign n3476 = ~\V133(10)  & n3475;
  assign n3477 = ~n525 & n2143;
  assign n3478 = ~n527 & n3477;
  assign n3479 = ~n3462 & n3478;
  assign n3480 = ~n529 & n3479;
  assign n3481 = ~n403 & n3480;
  assign n3482 = n530 & n3481;
  assign n3483 = \V47(1)  & n421;
  assign n3484 = n424 & n3483;
  assign n3485 = n434 & n3484;
  assign n3486 = ~n440 & n3485;
  assign n3487 = \V47(5)  & n434;
  assign n3488 = n424 & n3487;
  assign n3489 = ~n421 & n3488;
  assign n3490 = \V47(8)  & ~n434;
  assign n3491 = n424 & n3490;
  assign n3492 = \V47(16)  & ~n424;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = ~n3489 & n3493;
  assign n3495 = ~n3486 & n3494;
  assign n3496 = ~n443 & n3495;
  assign n3497 = ~n403 & ~n3496;
  assign n3498 = ~n529 & n3497;
  assign n3499 = ~n3462 & n3498;
  assign n3500 = ~n527 & n3499;
  assign n3501 = ~n525 & n3500;
  assign n3502 = \V133(10)  & n3501;
  assign n3503 = ~n525 & ~n3496;
  assign n3504 = ~n527 & n3503;
  assign n3505 = ~n3462 & n3504;
  assign n3506 = ~n529 & n3505;
  assign n3507 = n403 & n3506;
  assign n3508 = ~n529 & ~n3496;
  assign n3509 = ~n3462 & n3508;
  assign n3510 = ~n527 & n3509;
  assign n3511 = n525 & n3510;
  assign n3512 = ~n527 & ~n3496;
  assign n3513 = ~n3462 & n3512;
  assign n3514 = n529 & n3513;
  assign n3515 = n527 & ~n3496;
  assign n3516 = ~n3462 & n3515;
  assign n3517 = n3462 & ~n3496;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~n3514 & n3518;
  assign n3520 = ~n3511 & n3519;
  assign n3521 = ~n3507 & n3520;
  assign n3522 = ~n3502 & n3521;
  assign n3523 = ~n3482 & n3522;
  assign \V150(0)  = n3476 | ~n3523;
endmodule


