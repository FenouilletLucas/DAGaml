// Benchmark "i3" written by ABC on Tue May 16 16:07:50 2017

module i3 ( 
    \V132(5) , \V28(13) , \V126(1) , \V88(21) , \V132(4) , \V28(12) ,
    \V126(0) , \V88(20) , \V28(15) , \V28(14) , \V132(1) , \V132(0) ,
    \V28(11) , \V88(27) , \V28(10) , \V88(0) , \V88(26) , \V88(1) ,
    \V88(29) , \V88(2) , \V88(28) , \V88(3) , \V88(4) , \V28(17) ,
    \V88(5) , \V120(31) , \V28(16) , \V88(6) , \V120(30) , \V56(13) ,
    \V28(19) , \V88(7) , \V56(12) , \V28(18) , \V88(8) , \V56(15) ,
    \V28(23) , \V88(9) , \V88(31) , \V56(14) , \V28(22) , \V88(30) ,
    \V28(25) , \V28(24) , \V56(11) , \V56(10) , \V28(21) , \V28(20) ,
    \V120(27) , \V120(26) , \V120(29) , \V56(17) , \V120(28) , \V120(3) ,
    \V56(0) , \V56(16) , \V120(2) , \V56(1) , \V56(19) , \V28(27) ,
    \V120(5) , \V56(2) , \V56(18) , \V28(26) , \V120(4) , \V56(3) ,
    \V56(23) , \V56(4) , \V56(22) , \V56(5) , \V56(25) , \V120(1) ,
    \V56(6) , \V56(24) , \V120(21) , \V120(0) , \V56(7) , \V120(20) ,
    \V56(8) , \V120(23) , \V56(9) , \V56(21) , \V120(22) , \V56(20) ,
    \V120(25) , \V120(24) , \V120(7) , \V120(17) , \V120(6) , \V120(16) ,
    \V120(9) , \V120(19) , \V120(8) , \V56(27) , \V120(18) , \V56(26) ,
    \V88(13) , \V28(0) , \V88(12) , \V28(1) , \V88(15) , \V120(11) ,
    \V28(2) , \V88(14) , \V120(10) , \V28(3) , \V120(13) , \V28(4) ,
    \V120(12) , \V28(5) , \V88(11) , \V120(15) , \V28(6) , \V88(10) ,
    \V120(14) , \V28(7) , \V28(8) , \V28(9) , \V88(17) , \V88(16) ,
    \V88(19) , \V88(18) , \V126(3) , \V88(23) , \V126(2) , \V88(22) ,
    \V126(5) , \V88(25) , \V126(4) , \V88(24) , \V132(3) , \V132(2) ,
    \V138(3) , \V138(2) , \V134(1) , \V134(0) , \V138(1) , \V138(0)   );
  input  \V132(5) , \V28(13) , \V126(1) , \V88(21) , \V132(4) ,
    \V28(12) , \V126(0) , \V88(20) , \V28(15) , \V28(14) , \V132(1) ,
    \V132(0) , \V28(11) , \V88(27) , \V28(10) , \V88(0) , \V88(26) ,
    \V88(1) , \V88(29) , \V88(2) , \V88(28) , \V88(3) , \V88(4) ,
    \V28(17) , \V88(5) , \V120(31) , \V28(16) , \V88(6) , \V120(30) ,
    \V56(13) , \V28(19) , \V88(7) , \V56(12) , \V28(18) , \V88(8) ,
    \V56(15) , \V28(23) , \V88(9) , \V88(31) , \V56(14) , \V28(22) ,
    \V88(30) , \V28(25) , \V28(24) , \V56(11) , \V56(10) , \V28(21) ,
    \V28(20) , \V120(27) , \V120(26) , \V120(29) , \V56(17) , \V120(28) ,
    \V120(3) , \V56(0) , \V56(16) , \V120(2) , \V56(1) , \V56(19) ,
    \V28(27) , \V120(5) , \V56(2) , \V56(18) , \V28(26) , \V120(4) ,
    \V56(3) , \V56(23) , \V56(4) , \V56(22) , \V56(5) , \V56(25) ,
    \V120(1) , \V56(6) , \V56(24) , \V120(21) , \V120(0) , \V56(7) ,
    \V120(20) , \V56(8) , \V120(23) , \V56(9) , \V56(21) , \V120(22) ,
    \V56(20) , \V120(25) , \V120(24) , \V120(7) , \V120(17) , \V120(6) ,
    \V120(16) , \V120(9) , \V120(19) , \V120(8) , \V56(27) , \V120(18) ,
    \V56(26) , \V88(13) , \V28(0) , \V88(12) , \V28(1) , \V88(15) ,
    \V120(11) , \V28(2) , \V88(14) , \V120(10) , \V28(3) , \V120(13) ,
    \V28(4) , \V120(12) , \V28(5) , \V88(11) , \V120(15) , \V28(6) ,
    \V88(10) , \V120(14) , \V28(7) , \V28(8) , \V28(9) , \V88(17) ,
    \V88(16) , \V88(19) , \V88(18) , \V126(3) , \V88(23) , \V126(2) ,
    \V88(22) , \V126(5) , \V88(25) , \V126(4) , \V88(24) , \V132(3) ,
    \V132(2) ;
  output \V138(3) , \V138(2) , \V134(1) , \V134(0) , \V138(1) , \V138(0) ;
  wire n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447;
  assign n139 = ~\V126(3)  & ~\V132(3) ;
  assign n140 = ~\V126(2)  & ~\V132(2) ;
  assign n141 = ~\V126(1)  & ~\V132(1) ;
  assign n142 = ~\V126(0)  & ~\V132(0) ;
  assign n143 = ~\V120(31)  & ~\V88(31) ;
  assign n144 = ~\V120(30)  & ~\V88(30) ;
  assign n145 = ~\V88(29)  & ~\V120(29) ;
  assign n146 = ~\V88(28)  & ~\V120(28) ;
  assign n147 = ~\V88(27)  & ~\V120(27) ;
  assign n148 = ~\V88(26)  & ~\V120(26) ;
  assign n149 = ~\V120(25)  & ~\V88(25) ;
  assign n150 = ~\V120(24)  & ~\V88(24) ;
  assign n151 = ~\V120(23)  & ~\V88(23) ;
  assign n152 = ~\V120(22)  & ~\V88(22) ;
  assign n153 = \V126(5)  & \V126(4) ;
  assign n154 = ~n152 & n153;
  assign n155 = ~n151 & n154;
  assign n156 = ~n150 & n155;
  assign n157 = ~n149 & n156;
  assign n158 = ~n148 & n157;
  assign n159 = ~n147 & n158;
  assign n160 = ~n146 & n159;
  assign n161 = ~n145 & n160;
  assign n162 = ~n144 & n161;
  assign n163 = ~n143 & n162;
  assign n164 = ~n142 & n163;
  assign n165 = ~n141 & n164;
  assign n166 = ~n140 & n165;
  assign n167 = ~n139 & n166;
  assign n168 = \V132(4)  & \V126(5) ;
  assign n169 = ~n152 & n168;
  assign n170 = ~n151 & n169;
  assign n171 = ~n150 & n170;
  assign n172 = ~n149 & n171;
  assign n173 = ~n148 & n172;
  assign n174 = ~n147 & n173;
  assign n175 = ~n146 & n174;
  assign n176 = ~n145 & n175;
  assign n177 = ~n144 & n176;
  assign n178 = ~n143 & n177;
  assign n179 = ~n142 & n178;
  assign n180 = ~n141 & n179;
  assign n181 = ~n140 & n180;
  assign n182 = ~n139 & n181;
  assign n183 = \V132(5)  & \V126(4) ;
  assign n184 = ~n152 & n183;
  assign n185 = ~n151 & n184;
  assign n186 = ~n150 & n185;
  assign n187 = ~n149 & n186;
  assign n188 = ~n148 & n187;
  assign n189 = ~n147 & n188;
  assign n190 = ~n146 & n189;
  assign n191 = ~n145 & n190;
  assign n192 = ~n144 & n191;
  assign n193 = ~n143 & n192;
  assign n194 = ~n142 & n193;
  assign n195 = ~n141 & n194;
  assign n196 = ~n140 & n195;
  assign n197 = ~n139 & n196;
  assign n198 = \V132(5)  & \V132(4) ;
  assign n199 = ~n152 & n198;
  assign n200 = ~n151 & n199;
  assign n201 = ~n150 & n200;
  assign n202 = ~n149 & n201;
  assign n203 = ~n148 & n202;
  assign n204 = ~n147 & n203;
  assign n205 = ~n146 & n204;
  assign n206 = ~n145 & n205;
  assign n207 = ~n144 & n206;
  assign n208 = ~n143 & n207;
  assign n209 = ~n142 & n208;
  assign n210 = ~n141 & n209;
  assign n211 = ~n140 & n210;
  assign n212 = ~n139 & n211;
  assign n213 = ~n197 & ~n212;
  assign n214 = ~n182 & n213;
  assign \V138(3)  = n167 | ~n214;
  assign n216 = ~\V120(19)  & ~\V88(19) ;
  assign n217 = ~\V120(18)  & ~\V88(18) ;
  assign n218 = ~\V120(17)  & ~\V88(17) ;
  assign n219 = ~\V120(16)  & ~\V88(16) ;
  assign n220 = ~\V88(15)  & ~\V120(15) ;
  assign n221 = ~\V88(14)  & ~\V120(14) ;
  assign n222 = ~\V88(13)  & ~\V120(13) ;
  assign n223 = ~\V88(12)  & ~\V120(12) ;
  assign n224 = ~\V120(11)  & ~\V88(11) ;
  assign n225 = ~\V120(10)  & ~\V88(10) ;
  assign n226 = ~\V88(9)  & ~\V120(9) ;
  assign n227 = ~\V88(8)  & ~\V120(8) ;
  assign n228 = ~\V88(7)  & ~\V120(7) ;
  assign n229 = ~\V88(6)  & ~\V120(6) ;
  assign n230 = \V88(21)  & \V88(20) ;
  assign n231 = ~n229 & n230;
  assign n232 = ~n228 & n231;
  assign n233 = ~n227 & n232;
  assign n234 = ~n226 & n233;
  assign n235 = ~n225 & n234;
  assign n236 = ~n224 & n235;
  assign n237 = ~n223 & n236;
  assign n238 = ~n222 & n237;
  assign n239 = ~n221 & n238;
  assign n240 = ~n220 & n239;
  assign n241 = ~n219 & n240;
  assign n242 = ~n218 & n241;
  assign n243 = ~n217 & n242;
  assign n244 = ~n216 & n243;
  assign n245 = \V88(21)  & \V120(20) ;
  assign n246 = ~n229 & n245;
  assign n247 = ~n228 & n246;
  assign n248 = ~n227 & n247;
  assign n249 = ~n226 & n248;
  assign n250 = ~n225 & n249;
  assign n251 = ~n224 & n250;
  assign n252 = ~n223 & n251;
  assign n253 = ~n222 & n252;
  assign n254 = ~n221 & n253;
  assign n255 = ~n220 & n254;
  assign n256 = ~n219 & n255;
  assign n257 = ~n218 & n256;
  assign n258 = ~n217 & n257;
  assign n259 = ~n216 & n258;
  assign n260 = \V88(20)  & \V120(21) ;
  assign n261 = ~n229 & n260;
  assign n262 = ~n228 & n261;
  assign n263 = ~n227 & n262;
  assign n264 = ~n226 & n263;
  assign n265 = ~n225 & n264;
  assign n266 = ~n224 & n265;
  assign n267 = ~n223 & n266;
  assign n268 = ~n222 & n267;
  assign n269 = ~n221 & n268;
  assign n270 = ~n220 & n269;
  assign n271 = ~n219 & n270;
  assign n272 = ~n218 & n271;
  assign n273 = ~n217 & n272;
  assign n274 = ~n216 & n273;
  assign n275 = \V120(21)  & \V120(20) ;
  assign n276 = ~n229 & n275;
  assign n277 = ~n228 & n276;
  assign n278 = ~n227 & n277;
  assign n279 = ~n226 & n278;
  assign n280 = ~n225 & n279;
  assign n281 = ~n224 & n280;
  assign n282 = ~n223 & n281;
  assign n283 = ~n222 & n282;
  assign n284 = ~n221 & n283;
  assign n285 = ~n220 & n284;
  assign n286 = ~n219 & n285;
  assign n287 = ~n218 & n286;
  assign n288 = ~n217 & n287;
  assign n289 = ~n216 & n288;
  assign n290 = ~n274 & ~n289;
  assign n291 = ~n259 & n290;
  assign \V138(2)  = n244 | ~n291;
  assign \V134(1)  = \V56(1)  | \V28(1) ;
  assign \V134(0)  = \V56(0)  | \V28(0) ;
  assign n295 = ~\V88(3)  & ~\V120(3) ;
  assign n296 = ~\V88(2)  & ~\V120(2) ;
  assign n297 = ~\V88(1)  & ~\V120(1) ;
  assign n298 = ~\V88(0)  & ~\V120(0) ;
  assign n299 = ~\V28(27)  & ~\V56(27) ;
  assign n300 = ~\V28(26)  & ~\V56(26) ;
  assign n301 = ~\V28(25)  & ~\V56(25) ;
  assign n302 = ~\V28(24)  & ~\V56(24) ;
  assign n303 = ~\V28(23)  & ~\V56(23) ;
  assign n304 = ~\V28(22)  & ~\V56(22) ;
  assign n305 = ~\V28(21)  & ~\V56(21) ;
  assign n306 = ~\V28(20)  & ~\V56(20) ;
  assign n307 = ~\V28(19)  & ~\V56(19) ;
  assign n308 = ~\V28(18)  & ~\V56(18) ;
  assign n309 = \V88(4)  & \V88(5) ;
  assign n310 = ~n308 & n309;
  assign n311 = ~n307 & n310;
  assign n312 = ~n306 & n311;
  assign n313 = ~n305 & n312;
  assign n314 = ~n304 & n313;
  assign n315 = ~n303 & n314;
  assign n316 = ~n302 & n315;
  assign n317 = ~n301 & n316;
  assign n318 = ~n300 & n317;
  assign n319 = ~n299 & n318;
  assign n320 = ~n298 & n319;
  assign n321 = ~n297 & n320;
  assign n322 = ~n296 & n321;
  assign n323 = ~n295 & n322;
  assign n324 = \V88(5)  & \V120(4) ;
  assign n325 = ~n308 & n324;
  assign n326 = ~n307 & n325;
  assign n327 = ~n306 & n326;
  assign n328 = ~n305 & n327;
  assign n329 = ~n304 & n328;
  assign n330 = ~n303 & n329;
  assign n331 = ~n302 & n330;
  assign n332 = ~n301 & n331;
  assign n333 = ~n300 & n332;
  assign n334 = ~n299 & n333;
  assign n335 = ~n298 & n334;
  assign n336 = ~n297 & n335;
  assign n337 = ~n296 & n336;
  assign n338 = ~n295 & n337;
  assign n339 = \V88(4)  & \V120(5) ;
  assign n340 = ~n308 & n339;
  assign n341 = ~n307 & n340;
  assign n342 = ~n306 & n341;
  assign n343 = ~n305 & n342;
  assign n344 = ~n304 & n343;
  assign n345 = ~n303 & n344;
  assign n346 = ~n302 & n345;
  assign n347 = ~n301 & n346;
  assign n348 = ~n300 & n347;
  assign n349 = ~n299 & n348;
  assign n350 = ~n298 & n349;
  assign n351 = ~n297 & n350;
  assign n352 = ~n296 & n351;
  assign n353 = ~n295 & n352;
  assign n354 = \V120(5)  & \V120(4) ;
  assign n355 = ~n308 & n354;
  assign n356 = ~n307 & n355;
  assign n357 = ~n306 & n356;
  assign n358 = ~n305 & n357;
  assign n359 = ~n304 & n358;
  assign n360 = ~n303 & n359;
  assign n361 = ~n302 & n360;
  assign n362 = ~n301 & n361;
  assign n363 = ~n300 & n362;
  assign n364 = ~n299 & n363;
  assign n365 = ~n298 & n364;
  assign n366 = ~n297 & n365;
  assign n367 = ~n296 & n366;
  assign n368 = ~n295 & n367;
  assign n369 = ~n353 & ~n368;
  assign n370 = ~n338 & n369;
  assign \V138(1)  = n323 | ~n370;
  assign n372 = ~\V28(15)  & ~\V56(15) ;
  assign n373 = ~\V28(14)  & ~\V56(14) ;
  assign n374 = ~\V28(13)  & ~\V56(13) ;
  assign n375 = ~\V28(12)  & ~\V56(12) ;
  assign n376 = ~\V28(11)  & ~\V56(11) ;
  assign n377 = ~\V28(10)  & ~\V56(10) ;
  assign n378 = ~\V56(9)  & ~\V28(9) ;
  assign n379 = ~\V56(8)  & ~\V28(8) ;
  assign n380 = ~\V56(7)  & ~\V28(7) ;
  assign n381 = ~\V56(6)  & ~\V28(6) ;
  assign n382 = ~\V56(5)  & ~\V28(5) ;
  assign n383 = ~\V56(4)  & ~\V28(4) ;
  assign n384 = ~\V56(3)  & ~\V28(3) ;
  assign n385 = ~\V56(2)  & ~\V28(2) ;
  assign n386 = \V28(17)  & \V28(16) ;
  assign n387 = ~n385 & n386;
  assign n388 = ~n384 & n387;
  assign n389 = ~n383 & n388;
  assign n390 = ~n382 & n389;
  assign n391 = ~n381 & n390;
  assign n392 = ~n380 & n391;
  assign n393 = ~n379 & n392;
  assign n394 = ~n378 & n393;
  assign n395 = ~n377 & n394;
  assign n396 = ~n376 & n395;
  assign n397 = ~n375 & n396;
  assign n398 = ~n374 & n397;
  assign n399 = ~n373 & n398;
  assign n400 = ~n372 & n399;
  assign n401 = \V28(17)  & \V56(16) ;
  assign n402 = ~n385 & n401;
  assign n403 = ~n384 & n402;
  assign n404 = ~n383 & n403;
  assign n405 = ~n382 & n404;
  assign n406 = ~n381 & n405;
  assign n407 = ~n380 & n406;
  assign n408 = ~n379 & n407;
  assign n409 = ~n378 & n408;
  assign n410 = ~n377 & n409;
  assign n411 = ~n376 & n410;
  assign n412 = ~n375 & n411;
  assign n413 = ~n374 & n412;
  assign n414 = ~n373 & n413;
  assign n415 = ~n372 & n414;
  assign n416 = \V28(16)  & \V56(17) ;
  assign n417 = ~n385 & n416;
  assign n418 = ~n384 & n417;
  assign n419 = ~n383 & n418;
  assign n420 = ~n382 & n419;
  assign n421 = ~n381 & n420;
  assign n422 = ~n380 & n421;
  assign n423 = ~n379 & n422;
  assign n424 = ~n378 & n423;
  assign n425 = ~n377 & n424;
  assign n426 = ~n376 & n425;
  assign n427 = ~n375 & n426;
  assign n428 = ~n374 & n427;
  assign n429 = ~n373 & n428;
  assign n430 = ~n372 & n429;
  assign n431 = \V56(17)  & \V56(16) ;
  assign n432 = ~n385 & n431;
  assign n433 = ~n384 & n432;
  assign n434 = ~n383 & n433;
  assign n435 = ~n382 & n434;
  assign n436 = ~n381 & n435;
  assign n437 = ~n380 & n436;
  assign n438 = ~n379 & n437;
  assign n439 = ~n378 & n438;
  assign n440 = ~n377 & n439;
  assign n441 = ~n376 & n440;
  assign n442 = ~n375 & n441;
  assign n443 = ~n374 & n442;
  assign n444 = ~n373 & n443;
  assign n445 = ~n372 & n444;
  assign n446 = ~n430 & ~n445;
  assign n447 = ~n415 & n446;
  assign \V138(0)  = n400 | ~n447;
endmodule


