// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:20 2016

module TOP ( clock, 
    Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_, Pkey_251_,
    Pkey_250_, Pkey_249_, Pkey_248_, Pkey_247_, Pkey_246_, Pkey_245_,
    Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_, Pkey_239_,
    Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_, Pkey_233_,
    Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, Pkey_228_, Pkey_227_,
    Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_, Pkey_221_,
    Pkey_220_, Pkey_219_, Pkey_218_, Pkey_217_, Pkey_216_, Pkey_215_,
    Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_, Pkey_209_,
    Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_, Pkey_203_,
    Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, Pkey_198_, Pkey_197_,
    Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_, Pkey_191_,
    Pkey_190_, Pkey_189_, Pkey_188_, Pkey_187_, Pkey_186_, Pkey_185_,
    Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_, Pkey_179_,
    Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_, Pkey_173_,
    Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, Pkey_168_, Pkey_167_,
    Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_, Pkey_161_,
    Pkey_160_, Pkey_159_, Pkey_158_, Pkey_157_, Pkey_156_, Pkey_155_,
    Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_, Pkey_149_,
    Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_, Pkey_143_,
    Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, Pkey_138_, Pkey_137_,
    Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_, Pkey_131_,
    Pkey_130_, Pkey_129_, Pkey_128_, Pkey_127_, Pkey_126_, Pkey_125_,
    Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_, Pkey_119_,
    Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_, Pkey_113_,
    Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, Pkey_108_, Pkey_107_,
    Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_, Pkey_101_,
    Pkey_100_, Pkey_99_, Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_, Pkey_94_,
    Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, Pkey_88_, Pkey_87_,
    Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_, Pkey_80_,
    Pkey_79_, Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_, Pkey_73_,
    Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, Pkey_68_, Pkey_67_, Pkey_66_,
    Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_, Pkey_59_,
    Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_, Pkey_52_,
    Pkey_51_, Pkey_50_, Pkey_49_, Pkey_48_, Pkey_47_, Pkey_46_, Pkey_45_,
    Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_, Pkey_38_,
    Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_, Pkey_31_,
    Pkey_30_, Pkey_29_, Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_, Pkey_24_,
    Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, Pkey_18_, Pkey_17_,
    Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_, Pkey_10_,
    Pkey_9_, Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_, Pkey_3_, Pkey_2_,
    Pkey_1_, Pkey_0_, Pencrypt_0_, Pcount_3_, Pcount_2_, Pcount_1_,
    Pcount_0_, PCLK,
    Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_,
    Pdata_ready_0_, PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_,
    PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, PKSi_181_,
    PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_,
    PKSi_174_, PKSi_173_, PKSi_172_, PKSi_171_, PKSi_170_, PKSi_169_,
    PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_,
    PKSi_162_, PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_,
    PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, PKSi_151_,
    PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_,
    PKSi_144_, PKSi_143_, PKSi_142_, PKSi_141_, PKSi_140_, PKSi_139_,
    PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_,
    PKSi_132_, PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_,
    PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, PKSi_121_,
    PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_,
    PKSi_114_, PKSi_113_, PKSi_112_, PKSi_111_, PKSi_110_, PKSi_109_,
    PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_,
    PKSi_102_, PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_,
    PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, PKSi_91_, PKSi_90_,
    PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_,
    PKSi_82_, PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_,
    PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, PKSi_71_, PKSi_70_, PKSi_69_,
    PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_,
    PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_,
    PKSi_54_, PKSi_53_, PKSi_52_, PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_,
    PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, PKSi_41_,
    PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_,
    PKSi_33_, PKSi_32_, PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_,
    PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, PKSi_21_, PKSi_20_,
    PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_,
    PKSi_12_, PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_,
    PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, PKSi_1_, PKSi_0_  );
  input  clock;
  input  Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_,
    Pkey_251_, Pkey_250_, Pkey_249_, Pkey_248_, Pkey_247_, Pkey_246_,
    Pkey_245_, Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_,
    Pkey_239_, Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_,
    Pkey_233_, Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, Pkey_228_,
    Pkey_227_, Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_,
    Pkey_221_, Pkey_220_, Pkey_219_, Pkey_218_, Pkey_217_, Pkey_216_,
    Pkey_215_, Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_,
    Pkey_209_, Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_,
    Pkey_203_, Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, Pkey_198_,
    Pkey_197_, Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_,
    Pkey_191_, Pkey_190_, Pkey_189_, Pkey_188_, Pkey_187_, Pkey_186_,
    Pkey_185_, Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_,
    Pkey_179_, Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_,
    Pkey_173_, Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, Pkey_168_,
    Pkey_167_, Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_,
    Pkey_161_, Pkey_160_, Pkey_159_, Pkey_158_, Pkey_157_, Pkey_156_,
    Pkey_155_, Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_,
    Pkey_149_, Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_,
    Pkey_143_, Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, Pkey_138_,
    Pkey_137_, Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_,
    Pkey_131_, Pkey_130_, Pkey_129_, Pkey_128_, Pkey_127_, Pkey_126_,
    Pkey_125_, Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_,
    Pkey_119_, Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_,
    Pkey_113_, Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, Pkey_108_,
    Pkey_107_, Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_,
    Pkey_101_, Pkey_100_, Pkey_99_, Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_,
    Pkey_94_, Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, Pkey_88_,
    Pkey_87_, Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_,
    Pkey_80_, Pkey_79_, Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_,
    Pkey_73_, Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, Pkey_68_, Pkey_67_,
    Pkey_66_, Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_,
    Pkey_59_, Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_,
    Pkey_52_, Pkey_51_, Pkey_50_, Pkey_49_, Pkey_48_, Pkey_47_, Pkey_46_,
    Pkey_45_, Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_,
    Pkey_38_, Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_,
    Pkey_31_, Pkey_30_, Pkey_29_, Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_,
    Pkey_24_, Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, Pkey_18_,
    Pkey_17_, Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_,
    Pkey_10_, Pkey_9_, Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_,
    Pkey_3_, Pkey_2_, Pkey_1_, Pkey_0_, Pencrypt_0_, Pcount_3_, Pcount_2_,
    Pcount_1_, Pcount_0_, PCLK;
  output Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_,
    Pdata_ready_0_, PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_,
    PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, PKSi_181_,
    PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_,
    PKSi_174_, PKSi_173_, PKSi_172_, PKSi_171_, PKSi_170_, PKSi_169_,
    PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_,
    PKSi_162_, PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_,
    PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, PKSi_151_,
    PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_,
    PKSi_144_, PKSi_143_, PKSi_142_, PKSi_141_, PKSi_140_, PKSi_139_,
    PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_,
    PKSi_132_, PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_,
    PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, PKSi_121_,
    PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_,
    PKSi_114_, PKSi_113_, PKSi_112_, PKSi_111_, PKSi_110_, PKSi_109_,
    PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_,
    PKSi_102_, PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_,
    PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, PKSi_91_, PKSi_90_,
    PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_,
    PKSi_82_, PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_,
    PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, PKSi_71_, PKSi_70_, PKSi_69_,
    PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_,
    PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_,
    PKSi_54_, PKSi_53_, PKSi_52_, PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_,
    PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, PKSi_41_,
    PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_,
    PKSi_33_, PKSi_32_, PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_,
    PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, PKSi_21_, PKSi_20_,
    PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_,
    PKSi_12_, PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_,
    PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, PKSi_1_, PKSi_0_;
  reg PKSi_79_, PKSi_92_, \[333] , N_N2737, PKSi_75_, PKSi_84_, N_N2741,
    PKSi_82_, PKSi_93_, PKSi_85_, N_N2746, PKSi_73_, N_N2749, PKSi_80_,
    PKSi_72_, PKSi_94_, PKSi_86_, PKSi_74_, PKSi_83_, N_N2757, PKSi_89_,
    PKSi_91_, PKSi_81_, PKSi_77_, PKSi_87_, PKSi_78_, PKSi_95_, PKSi_76_,
    PKSi_55_, PKSi_68_, PKSi_64_, N_N2770, PKSi_51_, PKSi_60_, N_N2774,
    PKSi_58_, PKSi_69_, PKSi_61_, N_N2779, PKSi_49_, PKSi_66_, PKSi_56_,
    PKSi_48_, PKSi_70_, PKSi_62_, PKSi_50_, PKSi_59_, N_N2789, PKSi_65_,
    PKSi_67_, PKSi_57_, PKSi_53_, PKSi_63_, PKSi_54_, PKSi_71_, PKSi_52_,
    PKSi_31_, PKSi_44_, PKSi_40_, N_N2802, PKSi_27_, PKSi_36_, N_N2806,
    PKSi_34_, PKSi_45_, PKSi_37_, N_N2811, PKSi_25_, PKSi_42_, PKSi_32_,
    PKSi_24_, PKSi_46_, PKSi_38_, PKSi_26_, PKSi_35_, N_N2821, PKSi_41_,
    PKSi_43_, PKSi_33_, PKSi_29_, PKSi_39_, PKSi_30_, PKSi_47_, PKSi_28_,
    PKSi_7_, PKSi_20_, PKSi_16_, N_N2834, PKSi_3_, PKSi_12_, N_N2838,
    PKSi_10_, PKSi_21_, PKSi_13_, N_N2843, PKSi_1_, PKSi_18_, PKSi_8_,
    PKSi_0_, PKSi_22_, PKSi_14_, PKSi_2_, PKSi_11_, N_N2853, PKSi_17_,
    PKSi_19_, PKSi_9_, PKSi_5_, PKSi_15_, PKSi_6_, PKSi_23_, PKSi_4_,
    PKSi_183_, PKSi_173_, N_N2865, PKSi_185_, PKSi_169_, PKSi_176_,
    PKSi_188_, \[253] , PKSi_179_, PKSi_172_, PKSi_186_, PKSi_177_,
    PKSi_180_, N_N2877, N_N2879, N_N2881, PKSi_175_, PKSi_182_, N_N2885,
    PKSi_171_, PKSi_189_, N_N2889, PKSi_184_, PKSi_178_, \[234] ,
    PKSi_170_, PKSi_174_, PKSi_190_, PKSi_159_, PKSi_149_, N_N2899,
    PKSi_161_, PKSi_145_, PKSi_152_, PKSi_164_, PKSi_157_, PKSi_155_,
    PKSi_148_, PKSi_162_, N_N2909, PKSi_156_, PKSi_153_, PKSi_163_,
    PKSi_144_, PKSi_151_, PKSi_158_, N_N2917, PKSi_147_, PKSi_165_,
    N_N2921, PKSi_160_, PKSi_154_, PKSi_167_, PKSi_146_, PKSi_150_,
    PKSi_166_, PKSi_135_, PKSi_125_, N_N2931, PKSi_137_, PKSi_121_,
    PKSi_128_, PKSi_140_, PKSi_133_, PKSi_131_, PKSi_124_, PKSi_138_,
    PKSi_129_, PKSi_132_, N_N2943, N_N2945, PKSi_120_, PKSi_127_,
    PKSi_134_, N_N2950, PKSi_123_, PKSi_141_, N_N2954, PKSi_136_,
    PKSi_130_, \[282] , PKSi_122_, PKSi_126_, PKSi_142_, PKSi_111_,
    PKSi_101_, N_N2964, PKSi_113_, PKSi_97_, PKSi_104_, PKSi_116_,
    PKSi_109_, PKSi_107_, PKSi_100_, PKSi_114_, PKSi_105_, PKSi_108_,
    N_N2976, PKSi_115_, PKSi_96_, PKSi_103_, PKSi_110_, N_N2982, PKSi_99_,
    PKSi_117_, N_N2986, PKSi_112_, PKSi_106_, PKSi_119_, PKSi_98_,
    PKSi_102_, PKSi_118_;
  wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1165, n1166, n1167, n1168_1, n1170, n1172, n1174, n1175, n1176,
    n1177_1, n1178, n1179, n1180, n1181_1, n1182, n1183, n1184, n1185,
    n1186_1, n1187, n1188, n1189, n1190_1, n1191, n1192, n1193, n1194_1,
    n1195, n1196, n1197, n1198_1, n1199, n1200, n1202, n1203_1, n1204,
    n1205, n1206, n1207_1, n1208, n1209, n1210, n1211_1, n1212, n1213,
    n1214, n1216, n1217, n1218, n1219_1, n1220, n1221, n1222, n1223_1,
    n1224, n1225, n1226, n1227_1, n1228, n1230, n1231_1, n1232, n1233,
    n1234, n1235_1, n1236, n1237, n1238, n1239, n1240_1, n1241, n1242,
    n1244_1, n1245, n1246, n1247, n1248_1, n1249, n1250, n1251, n1252_1,
    n1253, n1254, n1255, n1256_1, n1258, n1259, n1260_1, n1261, n1262,
    n1263, n1264_1, n1265, n1266, n1267, n1268_1, n1269, n1270, n1272_1,
    n1273, n1274, n1275, n1276_1, n1277, n1278, n1279, n1280_1, n1281,
    n1282, n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742_1, n1743, n1744,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755_1,
    n1756, n1757, n1758, n1760, n1761, n1762, n1763_1, n1764, n1765, n1766,
    n1767_1, n1768, n1769, n1770, n1771_1, n1772, n1774, n1775_1, n1776,
    n1777, n1778, n1779_1, n1780, n1781, n1782, n1783_1, n1784, n1785,
    n1786, n1788, n1789, n1790, n1791_1, n1792, n1793, n1794, n1795_1,
    n1796, n1797, n1798, n1799, n1800, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1816, n1817,
    n1818, n1819, n1820, n1821_1, n1822, n1823, n1824, n1825_1, n1826,
    n1827, n1828, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
    n2387, n2388, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2736, n2737, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
    n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3556,
    n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3611,
    n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3622,
    n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3677,
    n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3732,
    n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n922_1, n926, n930_1,
    n935_1, n940_1, n944_1, n948_1, n953, n957, n961, n965, n970_1, n974_1,
    n979, n983, n987, n991, n995, n999, n1003, n1008_1, n1012_1, n1016_1,
    n1020_1, n1024_1, n1028_1, n1032_1, n1036_1, n1040_1, n1044_1, n1048_1,
    n1052_1, n1057, n1061, n1065, n1070_1, n1074_1, n1078_1, n1082_1,
    n1087, n1091, n1095, n1099, n1103, n1107, n1111, n1115, n1119, n1124_1,
    n1128_1, n1132_1, n1136_1, n1140_1, n1144_1, n1148_1, n1152_1, n1156_1,
    n1160_1, n1164, n1168, n1173, n1177, n1181, n1186, n1190, n1194, n1198,
    n1203, n1207, n1211, n1215, n1219, n1223, n1227, n1231, n1235, n1240,
    n1244, n1248, n1252, n1256, n1260, n1264, n1268, n1272, n1276, n1280,
    n1284_1, n1289_1, n1293_1, n1297_1, n1302_1, n1306_1, n1310_1, n1314_1,
    n1319_1, n1323_1, n1327_1, n1331_1, n1335_1, n1339_1, n1343_1, n1347_1,
    n1351_1, n1356_1, n1360_1, n1364_1, n1368_1, n1372_1, n1376_1, n1380_1,
    n1384_1, n1388_1, n1392_1, n1396_1, n1401_1, n1405_1, n1409_1, n1413_1,
    n1417_1, n1422_1, n1426_1, n1430_1, n1434_1, n1438_1, n1442_1, n1447_1,
    n1452_1, n1457_1, n1461_1, n1465_1, n1470_1, n1474_1, n1478_1, n1483_1,
    n1487_1, n1491_1, n1496_1, n1500_1, n1504_1, n1508_1, n1512_1, n1516_1,
    n1521_1, n1525_1, n1529_1, n1533_1, n1537_1, n1541_1, n1545_1, n1549_1,
    n1553_1, n1558_1, n1562_1, n1566_1, n1570_1, n1574_1, n1578_1, n1582_1,
    n1587_1, n1591_1, n1595_1, n1600_1, n1604_1, n1608_1, n1612_1, n1616_1,
    n1620_1, n1624_1, n1628_1, n1632_1, n1637_1, n1641_1, n1645_1, n1649_1,
    n1653_1, n1657_1, n1661_1, n1665_1, n1669_1, n1673_1, n1677_1, n1682_1,
    n1687_1, n1691_1, n1695_1, n1699_1, n1704_1, n1708_1, n1712_1, n1717_1,
    n1721_1, n1725_1, n1730_1, n1734_1, n1738_1, n1742, n1746_1, n1750_1,
    n1755, n1759, n1763, n1767, n1771, n1775, n1779, n1783, n1787, n1791,
    n1795, n1800_1, n1804_1, n1808_1, n1812_1, n1816_1, n1821, n1825,
    n1829, n1834_1, n1838_1, n1842_1, n1846_1, n1850_1, n1854_1;
  assign n1133 = ~Pcount_1_ & ~Pcount_0_;
  assign n1134 = ~Pcount_2_ & n1133;
  assign n1135 = ~Pencrypt_0_ & n1134;
  assign n1136 = ~Pstart_0_ & Pcount_3_;
  assign n1137 = Pcount_1_ & Pcount_0_;
  assign n1138 = Pcount_2_ & n1137;
  assign n1139 = Pencrypt_0_ & n1138;
  assign n1140 = n1136 & ~n1139;
  assign n1141 = ~n1135 & n1140;
  assign n1142 = ~Pcount_3_ & n1138;
  assign n1143 = ~Pstart_0_ & Pencrypt_0_;
  assign n1144 = n1142 & n1143;
  assign n1145 = Pstart_0_ & ~Pencrypt_0_;
  assign n1146 = ~Pstart_0_ & ~Pencrypt_0_;
  assign n1147 = ~Pcount_3_ & n1146;
  assign n1148 = n1134 & n1147;
  assign n1149 = ~n1145 & ~n1148;
  assign n1150 = ~n1144 & n1149;
  assign Pnew_count_3_ = n1141 | ~n1150;
  assign n1152 = ~Pencrypt_0_ & Pcount_1_;
  assign n1153 = ~Pcount_0_ & n1143;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = Pcount_2_ & ~n1154;
  assign n1156 = ~n1135 & ~n1155;
  assign n1157 = Pcount_2_ & Pcount_1_;
  assign n1158 = ~Pcount_2_ & ~Pcount_1_;
  assign n1159 = ~Pstart_0_ & Pcount_0_;
  assign n1160 = ~n1152 & n1159;
  assign n1161 = ~n1158 & n1160;
  assign n1162 = ~n1157 & n1161;
  assign n1163 = ~n1145 & ~n1162;
  assign Pnew_count_2_ = ~n1156 | ~n1163;
  assign n1165 = ~n1133 & ~n1137;
  assign n1166 = ~n1143 & ~n1145;
  assign n1167 = n1165 & ~n1166;
  assign n1168_1 = ~Pencrypt_0_ & ~n1165;
  assign Pnew_count_1_ = n1167 | n1168_1;
  assign n1170 = Pstart_0_ & Pencrypt_0_;
  assign Pnew_count_0_ = ~n1159 & ~n1170;
  assign n1172 = n1136 & n1139;
  assign Pdata_ready_0_ = n1148 | n1172;
  assign n1174 = Pkey_56_ & n1170;
  assign n1175 = Pkey_227_ & n1145;
  assign n1176 = ~PKSi_79_ & ~PKSi_183_;
  assign n1177_1 = Pcount_3_ & n1157;
  assign n1178 = Pcount_0_ & n1177_1;
  assign n1179 = ~Pcount_3_ & n1158;
  assign n1180 = ~n1134 & ~n1179;
  assign n1181_1 = ~n1178 & n1180;
  assign n1182 = n1146 & ~n1181_1;
  assign n1183 = n1176 & n1182;
  assign n1184 = n1146 & n1181_1;
  assign n1185 = ~n1176 & n1184;
  assign n1186_1 = ~n1183 & ~n1185;
  assign n1187 = ~n1175 & n1186_1;
  assign n1188 = ~n1174 & n1187;
  assign n1189 = PKSi_79_ & PKSi_183_;
  assign n1190_1 = ~n1177_1 & ~n1179;
  assign n1191 = ~Pcount_0_ & ~n1190_1;
  assign n1192 = ~n1142 & ~n1191;
  assign n1193 = ~Pstart_0_ & ~n1192;
  assign n1194_1 = ~n1146 & ~n1193;
  assign n1195 = n1189 & ~n1194_1;
  assign n1196 = ~n1176 & ~n1189;
  assign n1197 = ~Pstart_0_ & n1192;
  assign n1198_1 = Pencrypt_0_ & n1197;
  assign n1199 = n1196 & n1198_1;
  assign n1200 = ~n1195 & ~n1199;
  assign n922_1 = ~n1188 | ~n1200;
  assign n1202 = Pkey_227_ & n1170;
  assign n1203_1 = Pkey_235_ & n1145;
  assign n1204 = ~PKSi_92_ & ~PKSi_173_;
  assign n1205 = n1182 & n1204;
  assign n1206 = n1184 & ~n1204;
  assign n1207_1 = ~n1205 & ~n1206;
  assign n1208 = ~n1203_1 & n1207_1;
  assign n1209 = ~n1202 & n1208;
  assign n1210 = PKSi_92_ & PKSi_173_;
  assign n1211_1 = ~n1194_1 & n1210;
  assign n1212 = ~n1204 & ~n1210;
  assign n1213 = n1198_1 & n1212;
  assign n1214 = ~n1211_1 & ~n1213;
  assign n926 = ~n1209 | ~n1214;
  assign n1216 = Pkey_235_ & n1170;
  assign n1217 = Pkey_243_ & n1145;
  assign n1218 = ~\[333]  & ~N_N2865;
  assign n1219_1 = n1182 & n1218;
  assign n1220 = n1184 & ~n1218;
  assign n1221 = ~n1219_1 & ~n1220;
  assign n1222 = ~n1217 & n1221;
  assign n1223_1 = ~n1216 & n1222;
  assign n1224 = \[333]  & N_N2865;
  assign n1225 = ~n1194_1 & n1224;
  assign n1226 = ~n1218 & ~n1224;
  assign n1227_1 = n1198_1 & n1226;
  assign n1228 = ~n1225 & ~n1227_1;
  assign n930_1 = ~n1223_1 | ~n1228;
  assign n1230 = Pkey_243_ & n1170;
  assign n1231_1 = Pkey_251_ & n1145;
  assign n1232 = ~N_N2737 & ~PKSi_185_;
  assign n1233 = n1182 & n1232;
  assign n1234 = n1184 & ~n1232;
  assign n1235_1 = ~n1233 & ~n1234;
  assign n1236 = ~n1231_1 & n1235_1;
  assign n1237 = ~n1230 & n1236;
  assign n1238 = N_N2737 & PKSi_185_;
  assign n1239 = ~n1194_1 & n1238;
  assign n1240_1 = ~n1232 & ~n1238;
  assign n1241 = n1198_1 & n1240_1;
  assign n1242 = ~n1239 & ~n1241;
  assign n935_1 = ~n1237 | ~n1242;
  assign n1244_1 = Pkey_251_ & n1170;
  assign n1245 = Pkey_194_ & n1145;
  assign n1246 = ~PKSi_75_ & ~PKSi_169_;
  assign n1247 = n1182 & n1246;
  assign n1248_1 = n1184 & ~n1246;
  assign n1249 = ~n1247 & ~n1248_1;
  assign n1250 = ~n1245 & n1249;
  assign n1251 = ~n1244_1 & n1250;
  assign n1252_1 = PKSi_75_ & PKSi_169_;
  assign n1253 = ~n1194_1 & n1252_1;
  assign n1254 = ~n1246 & ~n1252_1;
  assign n1255 = n1198_1 & n1254;
  assign n1256_1 = ~n1253 & ~n1255;
  assign n940_1 = ~n1251 | ~n1256_1;
  assign n1258 = Pkey_194_ & n1170;
  assign n1259 = Pkey_202_ & n1145;
  assign n1260_1 = ~PKSi_84_ & ~PKSi_176_;
  assign n1261 = n1182 & n1260_1;
  assign n1262 = n1184 & ~n1260_1;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264_1 = ~n1259 & n1263;
  assign n1265 = ~n1258 & n1264_1;
  assign n1266 = PKSi_84_ & PKSi_176_;
  assign n1267 = ~n1194_1 & n1266;
  assign n1268_1 = ~n1260_1 & ~n1266;
  assign n1269 = n1198_1 & n1268_1;
  assign n1270 = ~n1267 & ~n1269;
  assign n944_1 = ~n1265 | ~n1270;
  assign n1272_1 = Pkey_202_ & n1170;
  assign n1273 = Pkey_210_ & n1145;
  assign n1274 = ~N_N2741 & ~PKSi_188_;
  assign n1275 = n1182 & n1274;
  assign n1276_1 = n1184 & ~n1274;
  assign n1277 = ~n1275 & ~n1276_1;
  assign n1278 = ~n1273 & n1277;
  assign n1279 = ~n1272_1 & n1278;
  assign n1280_1 = N_N2741 & PKSi_188_;
  assign n1281 = ~n1194_1 & n1280_1;
  assign n1282 = ~n1274 & ~n1280_1;
  assign n1283 = n1198_1 & n1282;
  assign n1284 = ~n1281 & ~n1283;
  assign n948_1 = ~n1279 | ~n1284;
  assign n1286 = Pkey_210_ & n1170;
  assign n1287 = Pkey_218_ & n1145;
  assign n1288 = ~PKSi_82_ & ~\[253] ;
  assign n1289 = n1182 & n1288;
  assign n1290 = n1184 & ~n1288;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1287 & n1291;
  assign n1293 = ~n1286 & n1292;
  assign n1294 = PKSi_82_ & \[253] ;
  assign n1295 = ~n1194_1 & n1294;
  assign n1296 = ~n1288 & ~n1294;
  assign n1297 = n1198_1 & n1296;
  assign n1298 = ~n1295 & ~n1297;
  assign n953 = ~n1293 | ~n1298;
  assign n1300 = Pkey_218_ & n1170;
  assign n1301 = Pkey_226_ & n1145;
  assign n1302 = ~PKSi_93_ & ~PKSi_179_;
  assign n1303 = n1182 & n1302;
  assign n1304 = n1184 & ~n1302;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = ~n1301 & n1305;
  assign n1307 = ~n1300 & n1306;
  assign n1308 = PKSi_93_ & PKSi_179_;
  assign n1309 = ~n1194_1 & n1308;
  assign n1310 = ~n1302 & ~n1308;
  assign n1311 = n1198_1 & n1310;
  assign n1312 = ~n1309 & ~n1311;
  assign n957 = ~n1307 | ~n1312;
  assign n1314 = Pkey_226_ & n1170;
  assign n1315 = Pkey_234_ & n1145;
  assign n1316 = ~PKSi_85_ & ~PKSi_172_;
  assign n1317 = n1182 & n1316;
  assign n1318 = n1184 & ~n1316;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~n1315 & n1319;
  assign n1321 = ~n1314 & n1320;
  assign n1322 = PKSi_85_ & PKSi_172_;
  assign n1323 = ~n1194_1 & n1322;
  assign n1324 = ~n1316 & ~n1322;
  assign n1325 = n1198_1 & n1324;
  assign n1326 = ~n1323 & ~n1325;
  assign n961 = ~n1321 | ~n1326;
  assign n1328 = N_N2746 & PKSi_186_;
  assign n1329 = ~n1194_1 & n1328;
  assign n1330 = ~N_N2746 & ~PKSi_186_;
  assign n1331 = n1198_1 & ~n1328;
  assign n1332 = ~n1184 & ~n1331;
  assign n1333 = ~n1330 & ~n1332;
  assign n1334 = Pkey_242_ & n1145;
  assign n1335 = Pkey_234_ & n1170;
  assign n1336 = n1182 & n1330;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = ~n1334 & n1337;
  assign n1339 = ~n1333 & n1338;
  assign n965 = n1329 | ~n1339;
  assign n1341 = Pkey_242_ & n1170;
  assign n1342 = Pkey_250_ & n1145;
  assign n1343 = ~PKSi_73_ & ~PKSi_177_;
  assign n1344 = n1182 & n1343;
  assign n1345 = n1184 & ~n1343;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n1342 & n1346;
  assign n1348 = ~n1341 & n1347;
  assign n1349 = PKSi_73_ & PKSi_177_;
  assign n1350 = ~n1194_1 & n1349;
  assign n1351 = ~n1343 & ~n1349;
  assign n1352 = n1198_1 & n1351;
  assign n1353 = ~n1350 & ~n1352;
  assign n970_1 = ~n1348 | ~n1353;
  assign n1355 = Pkey_193_ & n1145;
  assign n1356 = Pkey_250_ & n1170;
  assign n1357 = ~N_N2749 & ~PKSi_180_;
  assign n1358 = n1182 & n1357;
  assign n1359 = n1184 & ~n1357;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1356 & n1360;
  assign n1362 = ~n1355 & n1361;
  assign n1363 = N_N2749 & PKSi_180_;
  assign n1364 = ~n1194_1 & n1363;
  assign n1365 = ~n1357 & ~n1363;
  assign n1366 = n1198_1 & n1365;
  assign n1367 = ~n1364 & ~n1366;
  assign n974_1 = ~n1362 | ~n1367;
  assign n1369 = Pkey_201_ & n1145;
  assign n1370 = Pkey_193_ & n1170;
  assign n1371 = ~PKSi_80_ & ~N_N2877;
  assign n1372 = n1182 & n1371;
  assign n1373 = n1184 & ~n1371;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1370 & n1374;
  assign n1376 = ~n1369 & n1375;
  assign n1377 = PKSi_80_ & N_N2877;
  assign n1378 = ~n1194_1 & n1377;
  assign n1379 = ~n1371 & ~n1377;
  assign n1380 = n1198_1 & n1379;
  assign n1381 = ~n1378 & ~n1380;
  assign n979 = ~n1376 | ~n1381;
  assign n1383 = Pkey_209_ & n1145;
  assign n1384 = Pkey_201_ & n1170;
  assign n1385 = ~PKSi_72_ & ~N_N2879;
  assign n1386 = n1182 & n1385;
  assign n1387 = n1184 & ~n1385;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~n1384 & n1388;
  assign n1390 = ~n1383 & n1389;
  assign n1391 = PKSi_72_ & N_N2879;
  assign n1392 = ~n1194_1 & n1391;
  assign n1393 = ~n1385 & ~n1391;
  assign n1394 = n1198_1 & n1393;
  assign n1395 = ~n1392 & ~n1394;
  assign n983 = ~n1390 | ~n1395;
  assign n1397 = Pkey_209_ & n1170;
  assign n1398 = Pkey_217_ & n1145;
  assign n1399 = ~PKSi_94_ & ~N_N2881;
  assign n1400 = n1182 & n1399;
  assign n1401 = n1184 & ~n1399;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n1398 & n1402;
  assign n1404 = ~n1397 & n1403;
  assign n1405 = PKSi_94_ & N_N2881;
  assign n1406 = ~n1194_1 & n1405;
  assign n1407 = ~n1399 & ~n1405;
  assign n1408 = n1198_1 & n1407;
  assign n1409 = ~n1406 & ~n1408;
  assign n987 = ~n1404 | ~n1409;
  assign n1411 = Pkey_217_ & n1170;
  assign n1412 = Pkey_225_ & n1145;
  assign n1413 = ~PKSi_86_ & ~PKSi_175_;
  assign n1414 = n1182 & n1413;
  assign n1415 = n1184 & ~n1413;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1412 & n1416;
  assign n1418 = ~n1411 & n1417;
  assign n1419 = PKSi_86_ & PKSi_175_;
  assign n1420 = ~n1194_1 & n1419;
  assign n1421 = ~n1413 & ~n1419;
  assign n1422 = n1198_1 & n1421;
  assign n1423 = ~n1420 & ~n1422;
  assign n991 = ~n1418 | ~n1423;
  assign n1425 = Pkey_225_ & n1170;
  assign n1426 = Pkey_233_ & n1145;
  assign n1427 = ~PKSi_74_ & ~PKSi_182_;
  assign n1428 = n1182 & n1427;
  assign n1429 = n1184 & ~n1427;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = ~n1426 & n1430;
  assign n1432 = ~n1425 & n1431;
  assign n1433 = PKSi_74_ & PKSi_182_;
  assign n1434 = ~n1194_1 & n1433;
  assign n1435 = ~n1427 & ~n1433;
  assign n1436 = n1198_1 & n1435;
  assign n1437 = ~n1434 & ~n1436;
  assign n995 = ~n1432 | ~n1437;
  assign n1439 = Pkey_233_ & n1170;
  assign n1440 = Pkey_241_ & n1145;
  assign n1441 = ~PKSi_83_ & ~N_N2885;
  assign n1442 = n1182 & n1441;
  assign n1443 = n1184 & ~n1441;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1440 & n1444;
  assign n1446 = ~n1439 & n1445;
  assign n1447 = PKSi_83_ & N_N2885;
  assign n1448 = ~n1194_1 & n1447;
  assign n1449 = ~n1441 & ~n1447;
  assign n1450 = n1198_1 & n1449;
  assign n1451 = ~n1448 & ~n1450;
  assign n999 = ~n1446 | ~n1451;
  assign n1453 = Pkey_241_ & n1170;
  assign n1454 = Pkey_249_ & n1145;
  assign n1455 = ~N_N2757 & ~PKSi_171_;
  assign n1456 = n1182 & n1455;
  assign n1457 = n1184 & ~n1455;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1454 & n1458;
  assign n1460 = ~n1453 & n1459;
  assign n1461 = N_N2757 & PKSi_171_;
  assign n1462 = ~n1194_1 & n1461;
  assign n1463 = ~n1455 & ~n1461;
  assign n1464 = n1198_1 & n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1003 = ~n1460 | ~n1465;
  assign n1467 = Pkey_249_ & n1170;
  assign n1468 = Pkey_192_ & n1145;
  assign n1469 = ~PKSi_89_ & ~PKSi_189_;
  assign n1470 = n1182 & n1469;
  assign n1471 = n1184 & ~n1469;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n1468 & n1472;
  assign n1474 = ~n1467 & n1473;
  assign n1475 = PKSi_89_ & PKSi_189_;
  assign n1476 = ~n1194_1 & n1475;
  assign n1477 = ~n1469 & ~n1475;
  assign n1478 = n1198_1 & n1477;
  assign n1479 = ~n1476 & ~n1478;
  assign n1008_1 = ~n1474 | ~n1479;
  assign n1481 = Pkey_192_ & n1170;
  assign n1482 = Pkey_200_ & n1145;
  assign n1483 = ~PKSi_91_ & ~N_N2889;
  assign n1484 = n1182 & n1483;
  assign n1485 = n1184 & ~n1483;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = ~n1482 & n1486;
  assign n1488 = ~n1481 & n1487;
  assign n1489 = PKSi_91_ & N_N2889;
  assign n1490 = ~n1194_1 & n1489;
  assign n1491 = ~n1483 & ~n1489;
  assign n1492 = n1198_1 & n1491;
  assign n1493 = ~n1490 & ~n1492;
  assign n1012_1 = ~n1488 | ~n1493;
  assign n1495 = Pkey_200_ & n1170;
  assign n1496 = Pkey_208_ & n1145;
  assign n1497 = ~PKSi_81_ & ~PKSi_184_;
  assign n1498 = n1182 & n1497;
  assign n1499 = n1184 & ~n1497;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1496 & n1500;
  assign n1502 = ~n1495 & n1501;
  assign n1503 = PKSi_81_ & PKSi_184_;
  assign n1504 = ~n1194_1 & n1503;
  assign n1505 = ~n1497 & ~n1503;
  assign n1506 = n1198_1 & n1505;
  assign n1507 = ~n1504 & ~n1506;
  assign n1016_1 = ~n1502 | ~n1507;
  assign n1509 = Pkey_208_ & n1170;
  assign n1510 = Pkey_216_ & n1145;
  assign n1511 = ~PKSi_77_ & ~PKSi_178_;
  assign n1512 = n1182 & n1511;
  assign n1513 = n1184 & ~n1511;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1510 & n1514;
  assign n1516 = ~n1509 & n1515;
  assign n1517 = PKSi_77_ & PKSi_178_;
  assign n1518 = ~n1194_1 & n1517;
  assign n1519 = ~n1511 & ~n1517;
  assign n1520 = n1198_1 & n1519;
  assign n1521 = ~n1518 & ~n1520;
  assign n1020_1 = ~n1516 | ~n1521;
  assign n1523 = Pkey_216_ & n1170;
  assign n1524 = Pkey_224_ & n1145;
  assign n1525 = ~PKSi_87_ & ~\[234] ;
  assign n1526 = n1182 & n1525;
  assign n1527 = n1184 & ~n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1524 & n1528;
  assign n1530 = ~n1523 & n1529;
  assign n1531 = PKSi_87_ & \[234] ;
  assign n1532 = ~n1194_1 & n1531;
  assign n1533 = ~n1525 & ~n1531;
  assign n1534 = n1198_1 & n1533;
  assign n1535 = ~n1532 & ~n1534;
  assign n1024_1 = ~n1530 | ~n1535;
  assign n1537 = Pkey_224_ & n1170;
  assign n1538 = Pkey_232_ & n1145;
  assign n1539 = ~PKSi_78_ & ~PKSi_170_;
  assign n1540 = n1182 & n1539;
  assign n1541 = n1184 & ~n1539;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = ~n1538 & n1542;
  assign n1544 = ~n1537 & n1543;
  assign n1545 = PKSi_78_ & PKSi_170_;
  assign n1546 = ~n1194_1 & n1545;
  assign n1547 = ~n1539 & ~n1545;
  assign n1548 = n1198_1 & n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign n1028_1 = ~n1544 | ~n1549;
  assign n1551 = Pkey_232_ & n1170;
  assign n1552 = Pkey_240_ & n1145;
  assign n1553 = ~PKSi_95_ & ~PKSi_174_;
  assign n1554 = n1182 & n1553;
  assign n1555 = n1184 & ~n1553;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~n1552 & n1556;
  assign n1558 = ~n1551 & n1557;
  assign n1559 = PKSi_95_ & PKSi_174_;
  assign n1560 = ~n1194_1 & n1559;
  assign n1561 = ~n1553 & ~n1559;
  assign n1562 = n1198_1 & n1561;
  assign n1563 = ~n1560 & ~n1562;
  assign n1032_1 = ~n1558 | ~n1563;
  assign n1565 = Pkey_240_ & n1170;
  assign n1566 = Pkey_248_ & n1145;
  assign n1567 = ~PKSi_76_ & ~PKSi_190_;
  assign n1568 = n1182 & n1567;
  assign n1569 = n1184 & ~n1567;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1566 & n1570;
  assign n1572 = ~n1565 & n1571;
  assign n1573 = PKSi_76_ & PKSi_190_;
  assign n1574 = ~n1194_1 & n1573;
  assign n1575 = ~n1567 & ~n1573;
  assign n1576 = n1198_1 & n1575;
  assign n1577 = ~n1574 & ~n1576;
  assign n1036_1 = ~n1572 | ~n1577;
  assign n1579 = Pkey_248_ & n1170;
  assign n1580 = Pkey_163_ & n1145;
  assign n1581 = ~PKSi_55_ & ~PKSi_159_;
  assign n1582 = n1182 & n1581;
  assign n1583 = n1184 & ~n1581;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = ~n1580 & n1584;
  assign n1586 = ~n1579 & n1585;
  assign n1587 = PKSi_55_ & PKSi_159_;
  assign n1588 = ~n1194_1 & n1587;
  assign n1589 = ~n1581 & ~n1587;
  assign n1590 = n1198_1 & n1589;
  assign n1591 = ~n1588 & ~n1590;
  assign n1040_1 = ~n1586 | ~n1591;
  assign n1593 = Pkey_163_ & n1170;
  assign n1594 = Pkey_171_ & n1145;
  assign n1595 = ~PKSi_68_ & ~PKSi_149_;
  assign n1596 = n1182 & n1595;
  assign n1597 = n1184 & ~n1595;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1594 & n1598;
  assign n1600 = ~n1593 & n1599;
  assign n1601 = PKSi_68_ & PKSi_149_;
  assign n1602 = ~n1194_1 & n1601;
  assign n1603 = ~n1595 & ~n1601;
  assign n1604 = n1198_1 & n1603;
  assign n1605 = ~n1602 & ~n1604;
  assign n1044_1 = ~n1600 | ~n1605;
  assign n1607 = Pkey_179_ & n1145;
  assign n1608 = Pkey_171_ & n1170;
  assign n1609 = ~PKSi_64_ & ~N_N2899;
  assign n1610 = n1182 & n1609;
  assign n1611 = n1184 & ~n1609;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~n1608 & n1612;
  assign n1614 = ~n1607 & n1613;
  assign n1615 = PKSi_64_ & N_N2899;
  assign n1616 = ~n1194_1 & n1615;
  assign n1617 = ~n1609 & ~n1615;
  assign n1618 = n1198_1 & n1617;
  assign n1619 = ~n1616 & ~n1618;
  assign n1048_1 = ~n1614 | ~n1619;
  assign n1621 = Pkey_187_ & n1145;
  assign n1622 = Pkey_179_ & n1170;
  assign n1623 = ~N_N2770 & ~PKSi_161_;
  assign n1624 = n1182 & n1623;
  assign n1625 = n1184 & ~n1623;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~n1622 & n1626;
  assign n1628 = ~n1621 & n1627;
  assign n1629 = N_N2770 & PKSi_161_;
  assign n1630 = ~n1194_1 & n1629;
  assign n1631 = ~n1623 & ~n1629;
  assign n1632 = n1198_1 & n1631;
  assign n1633 = ~n1630 & ~n1632;
  assign n1052_1 = ~n1628 | ~n1633;
  assign n1635 = Pkey_187_ & n1170;
  assign n1636 = Pkey_130_ & n1145;
  assign n1637 = ~PKSi_51_ & ~PKSi_145_;
  assign n1638 = n1182 & n1637;
  assign n1639 = n1184 & ~n1637;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = ~n1636 & n1640;
  assign n1642 = ~n1635 & n1641;
  assign n1643 = PKSi_51_ & PKSi_145_;
  assign n1644 = ~n1194_1 & n1643;
  assign n1645 = ~n1637 & ~n1643;
  assign n1646 = n1198_1 & n1645;
  assign n1647 = ~n1644 & ~n1646;
  assign n1057 = ~n1642 | ~n1647;
  assign n1649 = Pkey_130_ & n1170;
  assign n1650 = Pkey_138_ & n1145;
  assign n1651 = ~PKSi_60_ & ~PKSi_152_;
  assign n1652 = n1182 & n1651;
  assign n1653 = n1184 & ~n1651;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1650 & n1654;
  assign n1656 = ~n1649 & n1655;
  assign n1657 = PKSi_60_ & PKSi_152_;
  assign n1658 = ~n1194_1 & n1657;
  assign n1659 = ~n1651 & ~n1657;
  assign n1660 = n1198_1 & n1659;
  assign n1661 = ~n1658 & ~n1660;
  assign n1061 = ~n1656 | ~n1661;
  assign n1663 = Pkey_146_ & n1145;
  assign n1664 = Pkey_138_ & n1170;
  assign n1665 = ~N_N2774 & ~PKSi_164_;
  assign n1666 = n1182 & n1665;
  assign n1667 = n1184 & ~n1665;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~n1664 & n1668;
  assign n1670 = ~n1663 & n1669;
  assign n1671 = N_N2774 & PKSi_164_;
  assign n1672 = ~n1194_1 & n1671;
  assign n1673 = ~n1665 & ~n1671;
  assign n1674 = n1198_1 & n1673;
  assign n1675 = ~n1672 & ~n1674;
  assign n1065 = ~n1670 | ~n1675;
  assign n1677 = Pkey_146_ & n1170;
  assign n1678 = ~PKSi_58_ & ~PKSi_157_;
  assign n1679 = n1182 & n1678;
  assign n1680 = ~n1677 & ~n1679;
  assign n1681 = PKSi_58_ & PKSi_157_;
  assign n1682 = ~n1194_1 & n1681;
  assign n1683 = Pkey_154_ & n1145;
  assign n1684 = n1184 & ~n1678;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1682 & n1685;
  assign n1687 = ~n1678 & ~n1681;
  assign n1688 = n1198_1 & n1687;
  assign n1689 = n1686 & ~n1688;
  assign n1070_1 = ~n1680 | ~n1689;
  assign n1691 = PKSi_69_ & PKSi_155_;
  assign n1692 = ~PKSi_69_ & ~PKSi_155_;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = n1198_1 & n1693;
  assign n1695 = ~n1194_1 & n1691;
  assign n1696 = n1182 & n1692;
  assign n1697 = n1184 & ~n1692;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = Pkey_154_ & n1170;
  assign n1700 = Pkey_162_ & n1145;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = n1698 & n1701;
  assign n1703 = ~n1695 & n1702;
  assign n1074_1 = n1694 | ~n1703;
  assign n1705 = Pkey_162_ & n1170;
  assign n1706 = Pkey_170_ & n1145;
  assign n1707 = ~PKSi_61_ & ~PKSi_148_;
  assign n1708 = n1182 & n1707;
  assign n1709 = n1184 & ~n1707;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~n1706 & n1710;
  assign n1712 = ~n1705 & n1711;
  assign n1713 = PKSi_61_ & PKSi_148_;
  assign n1714 = ~n1194_1 & n1713;
  assign n1715 = ~n1707 & ~n1713;
  assign n1716 = n1198_1 & n1715;
  assign n1717 = ~n1714 & ~n1716;
  assign n1078_1 = ~n1712 | ~n1717;
  assign n1719 = N_N2779 & PKSi_162_;
  assign n1720 = ~n1194_1 & n1719;
  assign n1721 = ~N_N2779 & ~PKSi_162_;
  assign n1722 = n1198_1 & ~n1719;
  assign n1723 = ~n1184 & ~n1722;
  assign n1724 = ~n1721 & ~n1723;
  assign n1725 = Pkey_170_ & n1170;
  assign n1726 = Pkey_178_ & n1145;
  assign n1727 = n1182 & n1721;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n1725 & n1728;
  assign n1730 = ~n1724 & n1729;
  assign n1082_1 = n1720 | ~n1730;
  assign n1732 = Pkey_178_ & n1170;
  assign n1733 = Pkey_186_ & n1145;
  assign n1734 = ~PKSi_49_ & ~N_N2909;
  assign n1735 = n1182 & n1734;
  assign n1736 = n1184 & ~n1734;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1733 & n1737;
  assign n1739 = ~n1732 & n1738;
  assign n1740 = PKSi_49_ & N_N2909;
  assign n1741 = ~n1194_1 & n1740;
  assign n1742_1 = ~n1734 & ~n1740;
  assign n1743 = n1198_1 & n1742_1;
  assign n1744 = ~n1741 & ~n1743;
  assign n1087 = ~n1739 | ~n1744;
  assign n1746 = Pkey_186_ & n1170;
  assign n1747 = Pkey_129_ & n1145;
  assign n1748 = ~PKSi_66_ & ~PKSi_156_;
  assign n1749 = n1182 & n1748;
  assign n1750 = n1184 & ~n1748;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = ~n1747 & n1751;
  assign n1753 = ~n1746 & n1752;
  assign n1754 = PKSi_66_ & PKSi_156_;
  assign n1755_1 = ~n1194_1 & n1754;
  assign n1756 = ~n1748 & ~n1754;
  assign n1757 = n1198_1 & n1756;
  assign n1758 = ~n1755_1 & ~n1757;
  assign n1091 = ~n1753 | ~n1758;
  assign n1760 = Pkey_129_ & n1170;
  assign n1761 = Pkey_137_ & n1145;
  assign n1762 = ~PKSi_56_ & ~PKSi_153_;
  assign n1763_1 = n1182 & n1762;
  assign n1764 = n1184 & ~n1762;
  assign n1765 = ~n1763_1 & ~n1764;
  assign n1766 = ~n1761 & n1765;
  assign n1767_1 = ~n1760 & n1766;
  assign n1768 = PKSi_56_ & PKSi_153_;
  assign n1769 = ~n1194_1 & n1768;
  assign n1770 = ~n1762 & ~n1768;
  assign n1771_1 = n1198_1 & n1770;
  assign n1772 = ~n1769 & ~n1771_1;
  assign n1095 = ~n1767_1 | ~n1772;
  assign n1774 = Pkey_137_ & n1170;
  assign n1775_1 = Pkey_145_ & n1145;
  assign n1776 = ~PKSi_48_ & ~PKSi_163_;
  assign n1777 = n1182 & n1776;
  assign n1778 = n1184 & ~n1776;
  assign n1779_1 = ~n1777 & ~n1778;
  assign n1780 = ~n1775_1 & n1779_1;
  assign n1781 = ~n1774 & n1780;
  assign n1782 = PKSi_48_ & PKSi_163_;
  assign n1783_1 = ~n1194_1 & n1782;
  assign n1784 = ~n1776 & ~n1782;
  assign n1785 = n1198_1 & n1784;
  assign n1786 = ~n1783_1 & ~n1785;
  assign n1099 = ~n1781 | ~n1786;
  assign n1788 = Pkey_145_ & n1170;
  assign n1789 = Pkey_153_ & n1145;
  assign n1790 = ~PKSi_70_ & ~PKSi_144_;
  assign n1791_1 = n1182 & n1790;
  assign n1792 = n1184 & ~n1790;
  assign n1793 = ~n1791_1 & ~n1792;
  assign n1794 = ~n1789 & n1793;
  assign n1795_1 = ~n1788 & n1794;
  assign n1796 = PKSi_70_ & PKSi_144_;
  assign n1797 = ~n1194_1 & n1796;
  assign n1798 = ~n1790 & ~n1796;
  assign n1799 = n1198_1 & n1798;
  assign n1800 = ~n1797 & ~n1799;
  assign n1103 = ~n1795_1 | ~n1800;
  assign n1802 = Pkey_153_ & n1170;
  assign n1803 = Pkey_161_ & n1145;
  assign n1804 = ~PKSi_62_ & ~PKSi_151_;
  assign n1805 = n1182 & n1804;
  assign n1806 = n1184 & ~n1804;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = ~n1803 & n1807;
  assign n1809 = ~n1802 & n1808;
  assign n1810 = PKSi_62_ & PKSi_151_;
  assign n1811 = ~n1194_1 & n1810;
  assign n1812 = ~n1804 & ~n1810;
  assign n1813 = n1198_1 & n1812;
  assign n1814 = ~n1811 & ~n1813;
  assign n1107 = ~n1809 | ~n1814;
  assign n1816 = Pkey_161_ & n1170;
  assign n1817 = Pkey_169_ & n1145;
  assign n1818 = ~PKSi_50_ & ~PKSi_158_;
  assign n1819 = n1182 & n1818;
  assign n1820 = n1184 & ~n1818;
  assign n1821_1 = ~n1819 & ~n1820;
  assign n1822 = ~n1817 & n1821_1;
  assign n1823 = ~n1816 & n1822;
  assign n1824 = PKSi_50_ & PKSi_158_;
  assign n1825_1 = ~n1194_1 & n1824;
  assign n1826 = ~n1818 & ~n1824;
  assign n1827 = n1198_1 & n1826;
  assign n1828 = ~n1825_1 & ~n1827;
  assign n1111 = ~n1823 | ~n1828;
  assign n1830 = PKSi_59_ & N_N2917;
  assign n1831 = ~PKSi_59_ & ~N_N2917;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1198_1 & n1832;
  assign n1834 = ~n1194_1 & n1830;
  assign n1835 = n1182 & n1831;
  assign n1836 = n1184 & ~n1831;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = Pkey_177_ & n1145;
  assign n1839 = Pkey_169_ & n1170;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = n1837 & n1840;
  assign n1842 = ~n1834 & n1841;
  assign n1115 = n1833 | ~n1842;
  assign n1844 = Pkey_185_ & n1145;
  assign n1845 = Pkey_177_ & n1170;
  assign n1846 = ~N_N2789 & ~PKSi_147_;
  assign n1847 = n1182 & n1846;
  assign n1848 = n1184 & ~n1846;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1845 & n1849;
  assign n1851 = ~n1844 & n1850;
  assign n1852 = N_N2789 & PKSi_147_;
  assign n1853 = ~n1194_1 & n1852;
  assign n1854 = ~n1846 & ~n1852;
  assign n1855 = n1198_1 & n1854;
  assign n1856 = ~n1853 & ~n1855;
  assign n1119 = ~n1851 | ~n1856;
  assign n1858 = Pkey_185_ & n1170;
  assign n1859 = Pkey_128_ & n1145;
  assign n1860 = ~PKSi_65_ & ~PKSi_165_;
  assign n1861 = n1182 & n1860;
  assign n1862 = n1184 & ~n1860;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = ~n1859 & n1863;
  assign n1865 = ~n1858 & n1864;
  assign n1866 = PKSi_65_ & PKSi_165_;
  assign n1867 = ~n1194_1 & n1866;
  assign n1868 = ~n1860 & ~n1866;
  assign n1869 = n1198_1 & n1868;
  assign n1870 = ~n1867 & ~n1869;
  assign n1124_1 = ~n1865 | ~n1870;
  assign n1872 = Pkey_128_ & n1170;
  assign n1873 = Pkey_136_ & n1145;
  assign n1874 = ~PKSi_67_ & ~N_N2921;
  assign n1875 = n1182 & n1874;
  assign n1876 = n1184 & ~n1874;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = ~n1873 & n1877;
  assign n1879 = ~n1872 & n1878;
  assign n1880 = PKSi_67_ & N_N2921;
  assign n1881 = ~n1194_1 & n1880;
  assign n1882 = ~n1874 & ~n1880;
  assign n1883 = n1198_1 & n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n1128_1 = ~n1879 | ~n1884;
  assign n1886 = Pkey_136_ & n1170;
  assign n1887 = Pkey_144_ & n1145;
  assign n1888 = ~PKSi_57_ & ~PKSi_160_;
  assign n1889 = n1182 & n1888;
  assign n1890 = n1184 & ~n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1887 & n1891;
  assign n1893 = ~n1886 & n1892;
  assign n1894 = PKSi_57_ & PKSi_160_;
  assign n1895 = ~n1194_1 & n1894;
  assign n1896 = ~n1888 & ~n1894;
  assign n1897 = n1198_1 & n1896;
  assign n1898 = ~n1895 & ~n1897;
  assign n1132_1 = ~n1893 | ~n1898;
  assign n1900 = Pkey_144_ & n1170;
  assign n1901 = Pkey_152_ & n1145;
  assign n1902 = ~PKSi_53_ & ~PKSi_154_;
  assign n1903 = n1182 & n1902;
  assign n1904 = n1184 & ~n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1901 & n1905;
  assign n1907 = ~n1900 & n1906;
  assign n1908 = PKSi_53_ & PKSi_154_;
  assign n1909 = ~n1194_1 & n1908;
  assign n1910 = ~n1902 & ~n1908;
  assign n1911 = n1198_1 & n1910;
  assign n1912 = ~n1909 & ~n1911;
  assign n1136_1 = ~n1907 | ~n1912;
  assign n1914 = Pkey_152_ & n1170;
  assign n1915 = Pkey_160_ & n1145;
  assign n1916 = ~PKSi_63_ & ~PKSi_167_;
  assign n1917 = n1182 & n1916;
  assign n1918 = n1184 & ~n1916;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = ~n1915 & n1919;
  assign n1921 = ~n1914 & n1920;
  assign n1922 = PKSi_63_ & PKSi_167_;
  assign n1923 = ~n1194_1 & n1922;
  assign n1924 = ~n1916 & ~n1922;
  assign n1925 = n1198_1 & n1924;
  assign n1926 = ~n1923 & ~n1925;
  assign n1140_1 = ~n1921 | ~n1926;
  assign n1928 = Pkey_160_ & n1170;
  assign n1929 = Pkey_168_ & n1145;
  assign n1930 = ~PKSi_54_ & ~PKSi_146_;
  assign n1931 = n1182 & n1930;
  assign n1932 = n1184 & ~n1930;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = ~n1929 & n1933;
  assign n1935 = ~n1928 & n1934;
  assign n1936 = PKSi_54_ & PKSi_146_;
  assign n1937 = ~n1194_1 & n1936;
  assign n1938 = ~n1930 & ~n1936;
  assign n1939 = n1198_1 & n1938;
  assign n1940 = ~n1937 & ~n1939;
  assign n1144_1 = ~n1935 | ~n1940;
  assign n1942 = Pkey_168_ & n1170;
  assign n1943 = Pkey_176_ & n1145;
  assign n1944 = ~PKSi_71_ & ~PKSi_150_;
  assign n1945 = n1182 & n1944;
  assign n1946 = n1184 & ~n1944;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1943 & n1947;
  assign n1949 = ~n1942 & n1948;
  assign n1950 = PKSi_71_ & PKSi_150_;
  assign n1951 = ~n1194_1 & n1950;
  assign n1952 = ~n1944 & ~n1950;
  assign n1953 = n1198_1 & n1952;
  assign n1954 = ~n1951 & ~n1953;
  assign n1148_1 = ~n1949 | ~n1954;
  assign n1956 = Pkey_176_ & n1170;
  assign n1957 = Pkey_184_ & n1145;
  assign n1958 = ~PKSi_52_ & ~PKSi_166_;
  assign n1959 = n1182 & n1958;
  assign n1960 = n1184 & ~n1958;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1957 & n1961;
  assign n1963 = ~n1956 & n1962;
  assign n1964 = PKSi_52_ & PKSi_166_;
  assign n1965 = ~n1194_1 & n1964;
  assign n1966 = ~n1958 & ~n1964;
  assign n1967 = n1198_1 & n1966;
  assign n1968 = ~n1965 & ~n1967;
  assign n1152_1 = ~n1963 | ~n1968;
  assign n1970 = Pkey_184_ & n1170;
  assign n1971 = Pkey_99_ & n1145;
  assign n1972 = ~PKSi_31_ & ~PKSi_135_;
  assign n1973 = n1182 & n1972;
  assign n1974 = n1184 & ~n1972;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = ~n1971 & n1975;
  assign n1977 = ~n1970 & n1976;
  assign n1978 = PKSi_31_ & PKSi_135_;
  assign n1979 = ~n1194_1 & n1978;
  assign n1980 = ~n1972 & ~n1978;
  assign n1981 = n1198_1 & n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1156_1 = ~n1977 | ~n1982;
  assign n1984 = Pkey_99_ & n1170;
  assign n1985 = Pkey_107_ & n1145;
  assign n1986 = ~PKSi_44_ & ~PKSi_125_;
  assign n1987 = n1182 & n1986;
  assign n1988 = n1184 & ~n1986;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1985 & n1989;
  assign n1991 = ~n1984 & n1990;
  assign n1992 = PKSi_44_ & PKSi_125_;
  assign n1993 = ~n1194_1 & n1992;
  assign n1994 = ~n1986 & ~n1992;
  assign n1995 = n1198_1 & n1994;
  assign n1996 = ~n1993 & ~n1995;
  assign n1160_1 = ~n1991 | ~n1996;
  assign n1998 = Pkey_115_ & n1145;
  assign n1999 = Pkey_107_ & n1170;
  assign n2000 = ~PKSi_40_ & ~N_N2931;
  assign n2001 = n1182 & n2000;
  assign n2002 = n1184 & ~n2000;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = ~n1999 & n2003;
  assign n2005 = ~n1998 & n2004;
  assign n2006 = PKSi_40_ & N_N2931;
  assign n2007 = ~n1194_1 & n2006;
  assign n2008 = ~n2000 & ~n2006;
  assign n2009 = n1198_1 & n2008;
  assign n2010 = ~n2007 & ~n2009;
  assign n1164 = ~n2005 | ~n2010;
  assign n2012 = Pkey_115_ & n1170;
  assign n2013 = Pkey_123_ & n1145;
  assign n2014 = ~N_N2802 & ~PKSi_137_;
  assign n2015 = n1182 & n2014;
  assign n2016 = n1184 & ~n2014;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n2013 & n2017;
  assign n2019 = ~n2012 & n2018;
  assign n2020 = N_N2802 & PKSi_137_;
  assign n2021 = ~n1194_1 & n2020;
  assign n2022 = ~n2014 & ~n2020;
  assign n2023 = n1198_1 & n2022;
  assign n2024 = ~n2021 & ~n2023;
  assign n1168 = ~n2019 | ~n2024;
  assign n2026 = Pkey_123_ & n1170;
  assign n2027 = Pkey_66_ & n1145;
  assign n2028 = ~PKSi_27_ & ~PKSi_121_;
  assign n2029 = n1182 & n2028;
  assign n2030 = n1184 & ~n2028;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~n2027 & n2031;
  assign n2033 = ~n2026 & n2032;
  assign n2034 = PKSi_27_ & PKSi_121_;
  assign n2035 = ~n1194_1 & n2034;
  assign n2036 = ~n2028 & ~n2034;
  assign n2037 = n1198_1 & n2036;
  assign n2038 = ~n2035 & ~n2037;
  assign n1173 = ~n2033 | ~n2038;
  assign n2040 = Pkey_66_ & n1170;
  assign n2041 = Pkey_74_ & n1145;
  assign n2042 = ~PKSi_36_ & ~PKSi_128_;
  assign n2043 = n1182 & n2042;
  assign n2044 = n1184 & ~n2042;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = ~n2041 & n2045;
  assign n2047 = ~n2040 & n2046;
  assign n2048 = PKSi_36_ & PKSi_128_;
  assign n2049 = ~n1194_1 & n2048;
  assign n2050 = ~n2042 & ~n2048;
  assign n2051 = n1198_1 & n2050;
  assign n2052 = ~n2049 & ~n2051;
  assign n1177 = ~n2047 | ~n2052;
  assign n2054 = N_N2806 & PKSi_140_;
  assign n2055 = ~N_N2806 & ~PKSi_140_;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = n1198_1 & n2056;
  assign n2058 = ~n1194_1 & n2054;
  assign n2059 = n1182 & n2055;
  assign n2060 = n1184 & ~n2055;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = Pkey_74_ & n1170;
  assign n2063 = Pkey_82_ & n1145;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = n2061 & n2064;
  assign n2066 = ~n2058 & n2065;
  assign n1181 = n2057 | ~n2066;
  assign n2068 = Pkey_82_ & n1170;
  assign n2069 = Pkey_90_ & n1145;
  assign n2070 = ~PKSi_34_ & ~PKSi_133_;
  assign n2071 = n1182 & n2070;
  assign n2072 = n1184 & ~n2070;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2069 & n2073;
  assign n2075 = ~n2068 & n2074;
  assign n2076 = PKSi_34_ & PKSi_133_;
  assign n2077 = ~n1194_1 & n2076;
  assign n2078 = ~n2070 & ~n2076;
  assign n2079 = n1198_1 & n2078;
  assign n2080 = ~n2077 & ~n2079;
  assign n1186 = ~n2075 | ~n2080;
  assign n2082 = Pkey_90_ & n1170;
  assign n2083 = Pkey_98_ & n1145;
  assign n2084 = ~PKSi_45_ & ~PKSi_131_;
  assign n2085 = n1182 & n2084;
  assign n2086 = n1184 & ~n2084;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = ~n2083 & n2087;
  assign n2089 = ~n2082 & n2088;
  assign n2090 = PKSi_45_ & PKSi_131_;
  assign n2091 = ~n1194_1 & n2090;
  assign n2092 = ~n2084 & ~n2090;
  assign n2093 = n1198_1 & n2092;
  assign n2094 = ~n2091 & ~n2093;
  assign n1190 = ~n2089 | ~n2094;
  assign n2096 = Pkey_98_ & n1170;
  assign n2097 = Pkey_106_ & n1145;
  assign n2098 = ~PKSi_37_ & ~PKSi_124_;
  assign n2099 = n1182 & n2098;
  assign n2100 = n1184 & ~n2098;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = ~n2097 & n2101;
  assign n2103 = ~n2096 & n2102;
  assign n2104 = PKSi_37_ & PKSi_124_;
  assign n2105 = ~n1194_1 & n2104;
  assign n2106 = ~n2098 & ~n2104;
  assign n2107 = n1198_1 & n2106;
  assign n2108 = ~n2105 & ~n2107;
  assign n1194 = ~n2103 | ~n2108;
  assign n2110 = Pkey_114_ & n1145;
  assign n2111 = Pkey_106_ & n1170;
  assign n2112 = ~N_N2811 & ~PKSi_138_;
  assign n2113 = n1182 & n2112;
  assign n2114 = n1184 & ~n2112;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = ~n2111 & n2115;
  assign n2117 = ~n2110 & n2116;
  assign n2118 = N_N2811 & PKSi_138_;
  assign n2119 = ~n1194_1 & n2118;
  assign n2120 = ~n2112 & ~n2118;
  assign n2121 = n1198_1 & n2120;
  assign n2122 = ~n2119 & ~n2121;
  assign n1198 = ~n2117 | ~n2122;
  assign n2124 = PKSi_25_ & PKSi_129_;
  assign n2125 = ~n1194_1 & n2124;
  assign n2126 = ~PKSi_25_ & ~PKSi_129_;
  assign n2127 = ~n2124 & ~n2126;
  assign n2128 = n1198_1 & n2127;
  assign n2129 = ~n2125 & ~n2128;
  assign n2130 = Pkey_122_ & n1145;
  assign n2131 = n1184 & ~n2126;
  assign n2132 = ~n2130 & ~n2131;
  assign n2133 = Pkey_114_ & n1170;
  assign n2134 = n1182 & n2126;
  assign n2135 = ~n2133 & ~n2134;
  assign n2136 = n2132 & n2135;
  assign n1203 = ~n2129 | ~n2136;
  assign n2138 = Pkey_122_ & n1170;
  assign n2139 = Pkey_65_ & n1145;
  assign n2140 = ~PKSi_42_ & ~PKSi_132_;
  assign n2141 = n1182 & n2140;
  assign n2142 = n1184 & ~n2140;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = ~n2139 & n2143;
  assign n2145 = ~n2138 & n2144;
  assign n2146 = PKSi_42_ & PKSi_132_;
  assign n2147 = ~n1194_1 & n2146;
  assign n2148 = ~n2140 & ~n2146;
  assign n2149 = n1198_1 & n2148;
  assign n2150 = ~n2147 & ~n2149;
  assign n1207 = ~n2145 | ~n2150;
  assign n2152 = Pkey_65_ & n1170;
  assign n2153 = Pkey_73_ & n1145;
  assign n2154 = ~PKSi_32_ & ~N_N2943;
  assign n2155 = n1182 & n2154;
  assign n2156 = n1184 & ~n2154;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = ~n2153 & n2157;
  assign n2159 = ~n2152 & n2158;
  assign n2160 = PKSi_32_ & N_N2943;
  assign n2161 = ~n1194_1 & n2160;
  assign n2162 = ~n2154 & ~n2160;
  assign n2163 = n1198_1 & n2162;
  assign n2164 = ~n2161 & ~n2163;
  assign n1211 = ~n2159 | ~n2164;
  assign n2166 = Pkey_81_ & n1145;
  assign n2167 = Pkey_73_ & n1170;
  assign n2168 = ~PKSi_24_ & ~N_N2945;
  assign n2169 = n1182 & n2168;
  assign n2170 = n1184 & ~n2168;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n2167 & n2171;
  assign n2173 = ~n2166 & n2172;
  assign n2174 = PKSi_24_ & N_N2945;
  assign n2175 = ~n1194_1 & n2174;
  assign n2176 = ~n2168 & ~n2174;
  assign n2177 = n1198_1 & n2176;
  assign n2178 = ~n2175 & ~n2177;
  assign n1215 = ~n2173 | ~n2178;
  assign n2180 = Pkey_81_ & n1170;
  assign n2181 = Pkey_89_ & n1145;
  assign n2182 = ~PKSi_46_ & ~PKSi_120_;
  assign n2183 = n1182 & n2182;
  assign n2184 = n1184 & ~n2182;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = ~n2181 & n2185;
  assign n2187 = ~n2180 & n2186;
  assign n2188 = PKSi_46_ & PKSi_120_;
  assign n2189 = ~n1194_1 & n2188;
  assign n2190 = ~n2182 & ~n2188;
  assign n2191 = n1198_1 & n2190;
  assign n2192 = ~n2189 & ~n2191;
  assign n1219 = ~n2187 | ~n2192;
  assign n2194 = Pkey_89_ & n1170;
  assign n2195 = Pkey_97_ & n1145;
  assign n2196 = ~PKSi_38_ & ~PKSi_127_;
  assign n2197 = n1182 & n2196;
  assign n2198 = n1184 & ~n2196;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2195 & n2199;
  assign n2201 = ~n2194 & n2200;
  assign n2202 = PKSi_38_ & PKSi_127_;
  assign n2203 = ~n1194_1 & n2202;
  assign n2204 = ~n2196 & ~n2202;
  assign n2205 = n1198_1 & n2204;
  assign n2206 = ~n2203 & ~n2205;
  assign n1223 = ~n2201 | ~n2206;
  assign n2208 = Pkey_97_ & n1170;
  assign n2209 = Pkey_105_ & n1145;
  assign n2210 = ~PKSi_26_ & ~PKSi_134_;
  assign n2211 = n1182 & n2210;
  assign n2212 = n1184 & ~n2210;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = ~n2209 & n2213;
  assign n2215 = ~n2208 & n2214;
  assign n2216 = PKSi_26_ & PKSi_134_;
  assign n2217 = ~n1194_1 & n2216;
  assign n2218 = ~n2210 & ~n2216;
  assign n2219 = n1198_1 & n2218;
  assign n2220 = ~n2217 & ~n2219;
  assign n1227 = ~n2215 | ~n2220;
  assign n2222 = Pkey_113_ & n1145;
  assign n2223 = Pkey_105_ & n1170;
  assign n2224 = ~PKSi_35_ & ~N_N2950;
  assign n2225 = n1182 & n2224;
  assign n2226 = n1184 & ~n2224;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = ~n2223 & n2227;
  assign n2229 = ~n2222 & n2228;
  assign n2230 = PKSi_35_ & N_N2950;
  assign n2231 = ~n1194_1 & n2230;
  assign n2232 = ~n2224 & ~n2230;
  assign n2233 = n1198_1 & n2232;
  assign n2234 = ~n2231 & ~n2233;
  assign n1231 = ~n2229 | ~n2234;
  assign n2236 = Pkey_113_ & n1170;
  assign n2237 = Pkey_121_ & n1145;
  assign n2238 = ~N_N2821 & ~PKSi_123_;
  assign n2239 = n1182 & n2238;
  assign n2240 = n1184 & ~n2238;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = ~n2237 & n2241;
  assign n2243 = ~n2236 & n2242;
  assign n2244 = N_N2821 & PKSi_123_;
  assign n2245 = ~n1194_1 & n2244;
  assign n2246 = ~n2238 & ~n2244;
  assign n2247 = n1198_1 & n2246;
  assign n2248 = ~n2245 & ~n2247;
  assign n1235 = ~n2243 | ~n2248;
  assign n2250 = Pkey_121_ & n1170;
  assign n2251 = Pkey_64_ & n1145;
  assign n2252 = ~PKSi_41_ & ~PKSi_141_;
  assign n2253 = n1182 & n2252;
  assign n2254 = n1184 & ~n2252;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = ~n2251 & n2255;
  assign n2257 = ~n2250 & n2256;
  assign n2258 = PKSi_41_ & PKSi_141_;
  assign n2259 = ~n1194_1 & n2258;
  assign n2260 = ~n2252 & ~n2258;
  assign n2261 = n1198_1 & n2260;
  assign n2262 = ~n2259 & ~n2261;
  assign n1240 = ~n2257 | ~n2262;
  assign n2264 = Pkey_72_ & n1145;
  assign n2265 = Pkey_64_ & n1170;
  assign n2266 = ~PKSi_43_ & ~N_N2954;
  assign n2267 = n1182 & n2266;
  assign n2268 = n1184 & ~n2266;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = ~n2265 & n2269;
  assign n2271 = ~n2264 & n2270;
  assign n2272 = PKSi_43_ & N_N2954;
  assign n2273 = ~n1194_1 & n2272;
  assign n2274 = ~n2266 & ~n2272;
  assign n2275 = n1198_1 & n2274;
  assign n2276 = ~n2273 & ~n2275;
  assign n1244 = ~n2271 | ~n2276;
  assign n2278 = PKSi_33_ & PKSi_136_;
  assign n2279 = ~PKSi_33_ & ~PKSi_136_;
  assign n2280 = ~n2278 & ~n2279;
  assign n2281 = n1198_1 & n2280;
  assign n2282 = ~n1194_1 & n2278;
  assign n2283 = n1182 & n2279;
  assign n2284 = n1184 & ~n2279;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = Pkey_72_ & n1170;
  assign n2287 = Pkey_80_ & n1145;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = n2285 & n2288;
  assign n2290 = ~n2282 & n2289;
  assign n1248 = n2281 | ~n2290;
  assign n2292 = PKSi_29_ & PKSi_130_;
  assign n2293 = ~n1194_1 & n2292;
  assign n2294 = ~PKSi_29_ & ~PKSi_130_;
  assign n2295 = ~n2292 & ~n2294;
  assign n2296 = n1198_1 & n2295;
  assign n2297 = ~n2293 & ~n2296;
  assign n2298 = Pkey_88_ & n1145;
  assign n2299 = n1184 & ~n2294;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = Pkey_80_ & n1170;
  assign n2302 = n1182 & n2294;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = n2300 & n2303;
  assign n1252 = ~n2297 | ~n2304;
  assign n2306 = Pkey_88_ & n1170;
  assign n2307 = Pkey_96_ & n1145;
  assign n2308 = ~PKSi_39_ & ~\[282] ;
  assign n2309 = n1182 & n2308;
  assign n2310 = n1184 & ~n2308;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = ~n2307 & n2311;
  assign n2313 = ~n2306 & n2312;
  assign n2314 = PKSi_39_ & \[282] ;
  assign n2315 = ~n1194_1 & n2314;
  assign n2316 = ~n2308 & ~n2314;
  assign n2317 = n1198_1 & n2316;
  assign n2318 = ~n2315 & ~n2317;
  assign n1256 = ~n2313 | ~n2318;
  assign n2320 = Pkey_96_ & n1170;
  assign n2321 = Pkey_104_ & n1145;
  assign n2322 = ~PKSi_30_ & ~PKSi_122_;
  assign n2323 = n1182 & n2322;
  assign n2324 = n1184 & ~n2322;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n2321 & n2325;
  assign n2327 = ~n2320 & n2326;
  assign n2328 = PKSi_30_ & PKSi_122_;
  assign n2329 = ~n1194_1 & n2328;
  assign n2330 = ~n2322 & ~n2328;
  assign n2331 = n1198_1 & n2330;
  assign n2332 = ~n2329 & ~n2331;
  assign n1260 = ~n2327 | ~n2332;
  assign n2334 = Pkey_104_ & n1170;
  assign n2335 = Pkey_112_ & n1145;
  assign n2336 = ~PKSi_47_ & ~PKSi_126_;
  assign n2337 = n1182 & n2336;
  assign n2338 = n1184 & ~n2336;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = ~n2335 & n2339;
  assign n2341 = ~n2334 & n2340;
  assign n2342 = PKSi_47_ & PKSi_126_;
  assign n2343 = ~n1194_1 & n2342;
  assign n2344 = ~n2336 & ~n2342;
  assign n2345 = n1198_1 & n2344;
  assign n2346 = ~n2343 & ~n2345;
  assign n1264 = ~n2341 | ~n2346;
  assign n2348 = Pkey_112_ & n1170;
  assign n2349 = Pkey_120_ & n1145;
  assign n2350 = ~PKSi_28_ & ~PKSi_142_;
  assign n2351 = n1182 & n2350;
  assign n2352 = n1184 & ~n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n2349 & n2353;
  assign n2355 = ~n2348 & n2354;
  assign n2356 = PKSi_28_ & PKSi_142_;
  assign n2357 = ~n1194_1 & n2356;
  assign n2358 = ~n2350 & ~n2356;
  assign n2359 = n1198_1 & n2358;
  assign n2360 = ~n2357 & ~n2359;
  assign n1268 = ~n2355 | ~n2360;
  assign n2362 = Pkey_120_ & n1170;
  assign n2363 = Pkey_35_ & n1145;
  assign n2364 = ~PKSi_7_ & ~PKSi_111_;
  assign n2365 = n1182 & n2364;
  assign n2366 = n1184 & ~n2364;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n2363 & n2367;
  assign n2369 = ~n2362 & n2368;
  assign n2370 = PKSi_7_ & PKSi_111_;
  assign n2371 = ~n1194_1 & n2370;
  assign n2372 = ~n2364 & ~n2370;
  assign n2373 = n1198_1 & n2372;
  assign n2374 = ~n2371 & ~n2373;
  assign n1272 = ~n2369 | ~n2374;
  assign n2376 = Pkey_35_ & n1170;
  assign n2377 = Pkey_43_ & n1145;
  assign n2378 = ~PKSi_20_ & ~PKSi_101_;
  assign n2379 = n1182 & n2378;
  assign n2380 = n1184 & ~n2378;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = ~n2377 & n2381;
  assign n2383 = ~n2376 & n2382;
  assign n2384 = PKSi_20_ & PKSi_101_;
  assign n2385 = ~n1194_1 & n2384;
  assign n2386 = ~n2378 & ~n2384;
  assign n2387 = n1198_1 & n2386;
  assign n2388 = ~n2385 & ~n2387;
  assign n1276 = ~n2383 | ~n2388;
  assign n2390 = Pkey_51_ & n1145;
  assign n2391 = Pkey_43_ & n1170;
  assign n2392 = ~PKSi_16_ & ~N_N2964;
  assign n2393 = n1182 & n2392;
  assign n2394 = n1184 & ~n2392;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~n2391 & n2395;
  assign n2397 = ~n2390 & n2396;
  assign n2398 = PKSi_16_ & N_N2964;
  assign n2399 = ~n1194_1 & n2398;
  assign n2400 = ~n2392 & ~n2398;
  assign n2401 = n1198_1 & n2400;
  assign n2402 = ~n2399 & ~n2401;
  assign n1280 = ~n2397 | ~n2402;
  assign n2404 = Pkey_59_ & n1145;
  assign n2405 = Pkey_51_ & n1170;
  assign n2406 = ~N_N2834 & ~PKSi_113_;
  assign n2407 = n1182 & n2406;
  assign n2408 = n1184 & ~n2406;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~n2405 & n2409;
  assign n2411 = ~n2404 & n2410;
  assign n2412 = N_N2834 & PKSi_113_;
  assign n2413 = ~n1194_1 & n2412;
  assign n2414 = ~n2406 & ~n2412;
  assign n2415 = n1198_1 & n2414;
  assign n2416 = ~n2413 & ~n2415;
  assign n1284_1 = ~n2411 | ~n2416;
  assign n2418 = Pkey_59_ & n1170;
  assign n2419 = Pkey_2_ & n1145;
  assign n2420 = ~PKSi_3_ & ~PKSi_97_;
  assign n2421 = n1182 & n2420;
  assign n2422 = n1184 & ~n2420;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~n2419 & n2423;
  assign n2425 = ~n2418 & n2424;
  assign n2426 = PKSi_3_ & PKSi_97_;
  assign n2427 = ~n1194_1 & n2426;
  assign n2428 = ~n2420 & ~n2426;
  assign n2429 = n1198_1 & n2428;
  assign n2430 = ~n2427 & ~n2429;
  assign n1289_1 = ~n2425 | ~n2430;
  assign n2432 = Pkey_2_ & n1170;
  assign n2433 = Pkey_10_ & n1145;
  assign n2434 = ~PKSi_12_ & ~PKSi_104_;
  assign n2435 = n1182 & n2434;
  assign n2436 = n1184 & ~n2434;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2433 & n2437;
  assign n2439 = ~n2432 & n2438;
  assign n2440 = PKSi_12_ & PKSi_104_;
  assign n2441 = ~n1194_1 & n2440;
  assign n2442 = ~n2434 & ~n2440;
  assign n2443 = n1198_1 & n2442;
  assign n2444 = ~n2441 & ~n2443;
  assign n1293_1 = ~n2439 | ~n2444;
  assign n2446 = Pkey_10_ & n1170;
  assign n2447 = Pkey_18_ & n1145;
  assign n2448 = ~N_N2838 & ~PKSi_116_;
  assign n2449 = n1182 & n2448;
  assign n2450 = n1184 & ~n2448;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = ~n2447 & n2451;
  assign n2453 = ~n2446 & n2452;
  assign n2454 = N_N2838 & PKSi_116_;
  assign n2455 = ~n1194_1 & n2454;
  assign n2456 = ~n2448 & ~n2454;
  assign n2457 = n1198_1 & n2456;
  assign n2458 = ~n2455 & ~n2457;
  assign n1297_1 = ~n2453 | ~n2458;
  assign n2460 = Pkey_18_ & n1170;
  assign n2461 = Pkey_26_ & n1145;
  assign n2462 = ~PKSi_10_ & ~PKSi_109_;
  assign n2463 = n1182 & n2462;
  assign n2464 = n1184 & ~n2462;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~n2461 & n2465;
  assign n2467 = ~n2460 & n2466;
  assign n2468 = PKSi_10_ & PKSi_109_;
  assign n2469 = ~n1194_1 & n2468;
  assign n2470 = ~n2462 & ~n2468;
  assign n2471 = n1198_1 & n2470;
  assign n2472 = ~n2469 & ~n2471;
  assign n1302_1 = ~n2467 | ~n2472;
  assign n2474 = Pkey_26_ & n1170;
  assign n2475 = Pkey_34_ & n1145;
  assign n2476 = ~PKSi_21_ & ~PKSi_107_;
  assign n2477 = n1182 & n2476;
  assign n2478 = n1184 & ~n2476;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = ~n2475 & n2479;
  assign n2481 = ~n2474 & n2480;
  assign n2482 = PKSi_21_ & PKSi_107_;
  assign n2483 = ~n1194_1 & n2482;
  assign n2484 = ~n2476 & ~n2482;
  assign n2485 = n1198_1 & n2484;
  assign n2486 = ~n2483 & ~n2485;
  assign n1306_1 = ~n2481 | ~n2486;
  assign n2488 = PKSi_13_ & PKSi_100_;
  assign n2489 = ~n1194_1 & n2488;
  assign n2490 = ~PKSi_13_ & ~PKSi_100_;
  assign n2491 = n1198_1 & ~n2488;
  assign n2492 = ~n1184 & ~n2491;
  assign n2493 = ~n2490 & ~n2492;
  assign n2494 = Pkey_42_ & n1145;
  assign n2495 = Pkey_34_ & n1170;
  assign n2496 = n1182 & n2490;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2494 & n2497;
  assign n2499 = ~n2493 & n2498;
  assign n1310_1 = n2489 | ~n2499;
  assign n2501 = Pkey_42_ & n1170;
  assign n2502 = Pkey_50_ & n1145;
  assign n2503 = ~N_N2843 & ~PKSi_114_;
  assign n2504 = n1182 & n2503;
  assign n2505 = n1184 & ~n2503;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = ~n2502 & n2506;
  assign n2508 = ~n2501 & n2507;
  assign n2509 = N_N2843 & PKSi_114_;
  assign n2510 = ~n1194_1 & n2509;
  assign n2511 = ~n2503 & ~n2509;
  assign n2512 = n1198_1 & n2511;
  assign n2513 = ~n2510 & ~n2512;
  assign n1314_1 = ~n2508 | ~n2513;
  assign n2515 = Pkey_50_ & n1170;
  assign n2516 = Pkey_58_ & n1145;
  assign n2517 = ~PKSi_1_ & ~PKSi_105_;
  assign n2518 = n1182 & n2517;
  assign n2519 = n1184 & ~n2517;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~n2516 & n2520;
  assign n2522 = ~n2515 & n2521;
  assign n2523 = PKSi_1_ & PKSi_105_;
  assign n2524 = ~n1194_1 & n2523;
  assign n2525 = ~n2517 & ~n2523;
  assign n2526 = n1198_1 & n2525;
  assign n2527 = ~n2524 & ~n2526;
  assign n1319_1 = ~n2522 | ~n2527;
  assign n2529 = Pkey_58_ & n1170;
  assign n2530 = Pkey_1_ & n1145;
  assign n2531 = ~PKSi_18_ & ~PKSi_108_;
  assign n2532 = n1182 & n2531;
  assign n2533 = n1184 & ~n2531;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = ~n2530 & n2534;
  assign n2536 = ~n2529 & n2535;
  assign n2537 = PKSi_18_ & PKSi_108_;
  assign n2538 = ~n1194_1 & n2537;
  assign n2539 = ~n2531 & ~n2537;
  assign n2540 = n1198_1 & n2539;
  assign n2541 = ~n2538 & ~n2540;
  assign n1323_1 = ~n2536 | ~n2541;
  assign n2543 = Pkey_9_ & n1145;
  assign n2544 = Pkey_1_ & n1170;
  assign n2545 = ~PKSi_8_ & ~N_N2976;
  assign n2546 = n1182 & n2545;
  assign n2547 = n1184 & ~n2545;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = ~n2544 & n2548;
  assign n2550 = ~n2543 & n2549;
  assign n2551 = PKSi_8_ & N_N2976;
  assign n2552 = ~n1194_1 & n2551;
  assign n2553 = ~n2545 & ~n2551;
  assign n2554 = n1198_1 & n2553;
  assign n2555 = ~n2552 & ~n2554;
  assign n1327_1 = ~n2550 | ~n2555;
  assign n2557 = Pkey_9_ & n1170;
  assign n2558 = Pkey_17_ & n1145;
  assign n2559 = ~PKSi_0_ & ~PKSi_115_;
  assign n2560 = n1182 & n2559;
  assign n2561 = n1184 & ~n2559;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n2558 & n2562;
  assign n2564 = ~n2557 & n2563;
  assign n2565 = PKSi_0_ & PKSi_115_;
  assign n2566 = ~n1194_1 & n2565;
  assign n2567 = ~n2559 & ~n2565;
  assign n2568 = n1198_1 & n2567;
  assign n2569 = ~n2566 & ~n2568;
  assign n1331_1 = ~n2564 | ~n2569;
  assign n2571 = PKSi_22_ & PKSi_96_;
  assign n2572 = ~n1194_1 & n2571;
  assign n2573 = ~PKSi_22_ & ~PKSi_96_;
  assign n2574 = ~n2571 & ~n2573;
  assign n2575 = n1198_1 & n2574;
  assign n2576 = ~n2572 & ~n2575;
  assign n2577 = Pkey_25_ & n1145;
  assign n2578 = n1184 & ~n2573;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = Pkey_17_ & n1170;
  assign n2581 = n1182 & n2573;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n2579 & n2582;
  assign n1335_1 = ~n2576 | ~n2583;
  assign n2585 = Pkey_25_ & n1170;
  assign n2586 = Pkey_33_ & n1145;
  assign n2587 = ~PKSi_14_ & ~PKSi_103_;
  assign n2588 = n1182 & n2587;
  assign n2589 = n1184 & ~n2587;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2586 & n2590;
  assign n2592 = ~n2585 & n2591;
  assign n2593 = PKSi_14_ & PKSi_103_;
  assign n2594 = ~n1194_1 & n2593;
  assign n2595 = ~n2587 & ~n2593;
  assign n2596 = n1198_1 & n2595;
  assign n2597 = ~n2594 & ~n2596;
  assign n1339_1 = ~n2592 | ~n2597;
  assign n2599 = Pkey_33_ & n1170;
  assign n2600 = Pkey_41_ & n1145;
  assign n2601 = ~PKSi_2_ & ~PKSi_110_;
  assign n2602 = n1182 & n2601;
  assign n2603 = n1184 & ~n2601;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = ~n2600 & n2604;
  assign n2606 = ~n2599 & n2605;
  assign n2607 = PKSi_2_ & PKSi_110_;
  assign n2608 = ~n1194_1 & n2607;
  assign n2609 = ~n2601 & ~n2607;
  assign n2610 = n1198_1 & n2609;
  assign n2611 = ~n2608 & ~n2610;
  assign n1343_1 = ~n2606 | ~n2611;
  assign n2613 = Pkey_49_ & n1145;
  assign n2614 = Pkey_41_ & n1170;
  assign n2615 = ~PKSi_11_ & ~N_N2982;
  assign n2616 = n1182 & n2615;
  assign n2617 = n1184 & ~n2615;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2614 & n2618;
  assign n2620 = ~n2613 & n2619;
  assign n2621 = PKSi_11_ & N_N2982;
  assign n2622 = ~n1194_1 & n2621;
  assign n2623 = ~n2615 & ~n2621;
  assign n2624 = n1198_1 & n2623;
  assign n2625 = ~n2622 & ~n2624;
  assign n1347_1 = ~n2620 | ~n2625;
  assign n2627 = Pkey_57_ & n1145;
  assign n2628 = Pkey_49_ & n1170;
  assign n2629 = ~N_N2853 & ~PKSi_99_;
  assign n2630 = n1182 & n2629;
  assign n2631 = n1184 & ~n2629;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2628 & n2632;
  assign n2634 = ~n2627 & n2633;
  assign n2635 = N_N2853 & PKSi_99_;
  assign n2636 = ~n1194_1 & n2635;
  assign n2637 = ~n2629 & ~n2635;
  assign n2638 = n1198_1 & n2637;
  assign n2639 = ~n2636 & ~n2638;
  assign n1351_1 = ~n2634 | ~n2639;
  assign n2641 = PKSi_17_ & PKSi_117_;
  assign n2642 = ~PKSi_17_ & ~PKSi_117_;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = n1198_1 & n2643;
  assign n2645 = ~n1194_1 & n2641;
  assign n2646 = n1182 & n2642;
  assign n2647 = n1184 & ~n2642;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = Pkey_57_ & n1170;
  assign n2650 = Pkey_0_ & n1145;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = n2648 & n2651;
  assign n2653 = ~n2645 & n2652;
  assign n1356_1 = n2644 | ~n2653;
  assign n2655 = Pkey_8_ & n1145;
  assign n2656 = Pkey_0_ & n1170;
  assign n2657 = ~PKSi_19_ & ~N_N2986;
  assign n2658 = n1182 & n2657;
  assign n2659 = n1184 & ~n2657;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2656 & n2660;
  assign n2662 = ~n2655 & n2661;
  assign n2663 = PKSi_19_ & N_N2986;
  assign n2664 = ~n1194_1 & n2663;
  assign n2665 = ~n2657 & ~n2663;
  assign n2666 = n1198_1 & n2665;
  assign n2667 = ~n2664 & ~n2666;
  assign n1360_1 = ~n2662 | ~n2667;
  assign n2669 = Pkey_8_ & n1170;
  assign n2670 = Pkey_16_ & n1145;
  assign n2671 = ~PKSi_9_ & ~PKSi_112_;
  assign n2672 = n1182 & n2671;
  assign n2673 = n1184 & ~n2671;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = ~n2670 & n2674;
  assign n2676 = ~n2669 & n2675;
  assign n2677 = PKSi_9_ & PKSi_112_;
  assign n2678 = ~n1194_1 & n2677;
  assign n2679 = ~n2671 & ~n2677;
  assign n2680 = n1198_1 & n2679;
  assign n2681 = ~n2678 & ~n2680;
  assign n1364_1 = ~n2676 | ~n2681;
  assign n2683 = Pkey_16_ & n1170;
  assign n2684 = Pkey_24_ & n1145;
  assign n2685 = ~PKSi_5_ & ~PKSi_106_;
  assign n2686 = n1182 & n2685;
  assign n2687 = n1184 & ~n2685;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = ~n2684 & n2688;
  assign n2690 = ~n2683 & n2689;
  assign n2691 = PKSi_5_ & PKSi_106_;
  assign n2692 = ~n1194_1 & n2691;
  assign n2693 = ~n2685 & ~n2691;
  assign n2694 = n1198_1 & n2693;
  assign n2695 = ~n2692 & ~n2694;
  assign n1368_1 = ~n2690 | ~n2695;
  assign n2697 = Pkey_24_ & n1170;
  assign n2698 = Pkey_32_ & n1145;
  assign n2699 = ~PKSi_15_ & ~PKSi_119_;
  assign n2700 = n1182 & n2699;
  assign n2701 = n1184 & ~n2699;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = ~n2698 & n2702;
  assign n2704 = ~n2697 & n2703;
  assign n2705 = PKSi_15_ & PKSi_119_;
  assign n2706 = ~n1194_1 & n2705;
  assign n2707 = ~n2699 & ~n2705;
  assign n2708 = n1198_1 & n2707;
  assign n2709 = ~n2706 & ~n2708;
  assign n1372_1 = ~n2704 | ~n2709;
  assign n2711 = PKSi_6_ & PKSi_98_;
  assign n2712 = ~n1194_1 & n2711;
  assign n2713 = ~PKSi_6_ & ~PKSi_98_;
  assign n2714 = ~n2711 & ~n2713;
  assign n2715 = n1198_1 & n2714;
  assign n2716 = ~n2712 & ~n2715;
  assign n2717 = Pkey_40_ & n1145;
  assign n2718 = n1184 & ~n2713;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = Pkey_32_ & n1170;
  assign n2721 = n1182 & n2713;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n2719 & n2722;
  assign n1376_1 = ~n2716 | ~n2723;
  assign n2725 = Pkey_40_ & n1170;
  assign n2726 = Pkey_48_ & n1145;
  assign n2727 = ~PKSi_23_ & ~PKSi_102_;
  assign n2728 = n1182 & n2727;
  assign n2729 = n1184 & ~n2727;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2726 & n2730;
  assign n2732 = ~n2725 & n2731;
  assign n2733 = PKSi_23_ & PKSi_102_;
  assign n2734 = ~n1194_1 & n2733;
  assign n2735 = ~n2727 & ~n2733;
  assign n2736 = n1198_1 & n2735;
  assign n2737 = ~n2734 & ~n2736;
  assign n1380_1 = ~n2732 | ~n2737;
  assign n2739 = Pkey_48_ & n1170;
  assign n2740 = Pkey_56_ & n1145;
  assign n2741 = ~PKSi_4_ & ~PKSi_118_;
  assign n2742 = n1182 & n2741;
  assign n2743 = n1184 & ~n2741;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = ~n2740 & n2744;
  assign n2746 = ~n2739 & n2745;
  assign n2747 = PKSi_4_ & PKSi_118_;
  assign n2748 = ~n1194_1 & n2747;
  assign n2749 = ~n2741 & ~n2747;
  assign n2750 = n1198_1 & n2749;
  assign n2751 = ~n2748 & ~n2750;
  assign n1384_1 = ~n2746 | ~n2751;
  assign n2753 = n1176 & n1184;
  assign n2754 = Pkey_62_ & n1170;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = ~n1146 & ~n1197;
  assign n2757 = n1189 & ~n2756;
  assign n2758 = n1143 & ~n1192;
  assign n2759 = n1196 & n2758;
  assign n2760 = ~n1176 & n1182;
  assign n2761 = Pkey_195_ & n1145;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2759 & n2762;
  assign n2764 = ~n2757 & n2763;
  assign n1388_1 = ~n2755 | ~n2764;
  assign n2766 = n1184 & n1204;
  assign n2767 = Pkey_203_ & n1145;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = n1210 & ~n2756;
  assign n2770 = n1212 & n2758;
  assign n2771 = n1182 & ~n1204;
  assign n2772 = Pkey_195_ & n1170;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = ~n2770 & n2773;
  assign n2775 = ~n2769 & n2774;
  assign n1392_1 = ~n2768 | ~n2775;
  assign n2777 = n1184 & n1218;
  assign n2778 = Pkey_203_ & n1170;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = n1224 & ~n2756;
  assign n2781 = n1226 & n2758;
  assign n2782 = n1182 & ~n1218;
  assign n2783 = Pkey_211_ & n1145;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = ~n2781 & n2784;
  assign n2786 = ~n2780 & n2785;
  assign n1396_1 = ~n2779 | ~n2786;
  assign n2788 = n1184 & n1232;
  assign n2789 = Pkey_211_ & n1170;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = n1238 & ~n2756;
  assign n2792 = n1240_1 & n2758;
  assign n2793 = n1182 & ~n1232;
  assign n2794 = Pkey_219_ & n1145;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2792 & n2795;
  assign n2797 = ~n2791 & n2796;
  assign n1401_1 = ~n2790 | ~n2797;
  assign n2799 = n1184 & n1246;
  assign n2800 = Pkey_196_ & n1145;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n1252_1 & ~n2756;
  assign n2803 = n1254 & n2758;
  assign n2804 = n1182 & ~n1246;
  assign n2805 = Pkey_219_ & n1170;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = ~n2803 & n2806;
  assign n2808 = ~n2802 & n2807;
  assign n1405_1 = ~n2801 | ~n2808;
  assign n2810 = n1184 & n1260_1;
  assign n2811 = Pkey_196_ & n1170;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = n1266 & ~n2756;
  assign n2814 = n1268_1 & n2758;
  assign n2815 = n1182 & ~n1260_1;
  assign n2816 = Pkey_204_ & n1145;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n2814 & n2817;
  assign n2819 = ~n2813 & n2818;
  assign n1409_1 = ~n2812 | ~n2819;
  assign n2821 = n1184 & n1274;
  assign n2822 = Pkey_212_ & n1145;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n1280_1 & ~n2756;
  assign n2825 = n1282 & n2758;
  assign n2826 = n1182 & ~n1274;
  assign n2827 = Pkey_204_ & n1170;
  assign n2828 = ~n2826 & ~n2827;
  assign n2829 = ~n2825 & n2828;
  assign n2830 = ~n2824 & n2829;
  assign n1413_1 = ~n2823 | ~n2830;
  assign n2832 = n1184 & n1288;
  assign n2833 = Pkey_212_ & n1170;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = n1294 & ~n2756;
  assign n2836 = n1296 & n2758;
  assign n2837 = n1182 & ~n1288;
  assign n2838 = Pkey_220_ & n1145;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = ~n2836 & n2839;
  assign n2841 = ~n2835 & n2840;
  assign n1417_1 = ~n2834 | ~n2841;
  assign n2843 = n1184 & n1302;
  assign n2844 = Pkey_220_ & n1170;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = n1308 & ~n2756;
  assign n2847 = n1310 & n2758;
  assign n2848 = n1182 & ~n1302;
  assign n2849 = Pkey_228_ & n1145;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2847 & n2850;
  assign n2852 = ~n2846 & n2851;
  assign n1422_1 = ~n2845 | ~n2852;
  assign n2854 = n1184 & n1316;
  assign n2855 = Pkey_228_ & n1170;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = n1322 & ~n2756;
  assign n2858 = n1324 & n2758;
  assign n2859 = n1182 & ~n1316;
  assign n2860 = Pkey_172_ & n1145;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2858 & n2861;
  assign n2863 = ~n2857 & n2862;
  assign n1426_1 = ~n2856 | ~n2863;
  assign n2865 = n1328 & ~n2756;
  assign n2866 = ~n1328 & n2758;
  assign n2867 = ~n1182 & ~n2866;
  assign n2868 = ~n1330 & ~n2867;
  assign n2869 = n1184 & n1330;
  assign n2870 = Pkey_172_ & n1170;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = Pkey_244_ & n1145;
  assign n2873 = n2871 & ~n2872;
  assign n2874 = ~n2868 & n2873;
  assign n1430_1 = n2865 | ~n2874;
  assign n2876 = n1184 & n1343;
  assign n2877 = Pkey_244_ & n1170;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = n1349 & ~n2756;
  assign n2880 = n1351 & n2758;
  assign n2881 = n1182 & ~n1343;
  assign n2882 = Pkey_252_ & n1145;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = ~n2880 & n2883;
  assign n2885 = ~n2879 & n2884;
  assign n1434_1 = ~n2878 | ~n2885;
  assign n2887 = n1184 & n1357;
  assign n2888 = Pkey_252_ & n1170;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = n1363 & ~n2756;
  assign n2891 = n1365 & n2758;
  assign n2892 = n1182 & ~n1357;
  assign n2893 = Pkey_197_ & n1145;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = ~n2891 & n2894;
  assign n2896 = ~n2890 & n2895;
  assign n1438_1 = ~n2889 | ~n2896;
  assign n2898 = n1184 & n1371;
  assign n2899 = Pkey_197_ & n1170;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = n1377 & ~n2756;
  assign n2902 = n1379 & n2758;
  assign n2903 = n1182 & ~n1371;
  assign n2904 = Pkey_205_ & n1145;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = ~n2902 & n2905;
  assign n2907 = ~n2901 & n2906;
  assign n1442_1 = ~n2900 | ~n2907;
  assign n2909 = n1184 & n1385;
  assign n2910 = Pkey_213_ & n1145;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = n1391 & ~n2756;
  assign n2913 = n1393 & n2758;
  assign n2914 = n1182 & ~n1385;
  assign n2915 = Pkey_205_ & n1170;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = ~n2913 & n2916;
  assign n2918 = ~n2912 & n2917;
  assign n1447_1 = ~n2911 | ~n2918;
  assign n2920 = n1184 & n1399;
  assign n2921 = Pkey_213_ & n1170;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = n1405 & ~n2756;
  assign n2924 = n1407 & n2758;
  assign n2925 = n1182 & ~n1399;
  assign n2926 = Pkey_221_ & n1145;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = ~n2924 & n2927;
  assign n2929 = ~n2923 & n2928;
  assign n1452_1 = ~n2922 | ~n2929;
  assign n2931 = n1184 & n1413;
  assign n2932 = Pkey_221_ & n1170;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = n1419 & ~n2756;
  assign n2935 = n1421 & n2758;
  assign n2936 = n1182 & ~n1413;
  assign n2937 = Pkey_229_ & n1145;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = ~n2935 & n2938;
  assign n2940 = ~n2934 & n2939;
  assign n1457_1 = ~n2933 | ~n2940;
  assign n2942 = n1184 & n1427;
  assign n2943 = Pkey_237_ & n1145;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = n1433 & ~n2756;
  assign n2946 = n1435 & n2758;
  assign n2947 = n1182 & ~n1427;
  assign n2948 = Pkey_229_ & n1170;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = ~n2946 & n2949;
  assign n2951 = ~n2945 & n2950;
  assign n1461_1 = ~n2944 | ~n2951;
  assign n2953 = n1184 & n1441;
  assign n2954 = Pkey_245_ & n1145;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = n1447 & ~n2756;
  assign n2957 = n1449 & n2758;
  assign n2958 = n1182 & ~n1441;
  assign n2959 = Pkey_237_ & n1170;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = ~n2957 & n2960;
  assign n2962 = ~n2956 & n2961;
  assign n1465_1 = ~n2955 | ~n2962;
  assign n2964 = n1184 & n1455;
  assign n2965 = Pkey_245_ & n1170;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = n1461 & ~n2756;
  assign n2968 = n1463 & n2758;
  assign n2969 = n1182 & ~n1455;
  assign n2970 = Pkey_253_ & n1145;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = ~n2968 & n2971;
  assign n2973 = ~n2967 & n2972;
  assign n1470_1 = ~n2966 | ~n2973;
  assign n2975 = n1184 & n1469;
  assign n2976 = Pkey_253_ & n1170;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = n1475 & ~n2756;
  assign n2979 = n1477 & n2758;
  assign n2980 = n1182 & ~n1469;
  assign n2981 = Pkey_198_ & n1145;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2979 & n2982;
  assign n2984 = ~n2978 & n2983;
  assign n1474_1 = ~n2977 | ~n2984;
  assign n2986 = n1184 & n1483;
  assign n2987 = Pkey_206_ & n1145;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = n1489 & ~n2756;
  assign n2990 = n1491 & n2758;
  assign n2991 = n1182 & ~n1483;
  assign n2992 = Pkey_198_ & n1170;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = ~n2990 & n2993;
  assign n2995 = ~n2989 & n2994;
  assign n1478_1 = ~n2988 | ~n2995;
  assign n2997 = n1184 & n1497;
  assign n2998 = Pkey_214_ & n1145;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = n1503 & ~n2756;
  assign n3001 = n1505 & n2758;
  assign n3002 = n1182 & ~n1497;
  assign n3003 = Pkey_206_ & n1170;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = ~n3001 & n3004;
  assign n3006 = ~n3000 & n3005;
  assign n1483_1 = ~n2999 | ~n3006;
  assign n3008 = n1184 & n1511;
  assign n3009 = Pkey_222_ & n1145;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n1517 & ~n2756;
  assign n3012 = n1519 & n2758;
  assign n3013 = n1182 & ~n1511;
  assign n3014 = Pkey_214_ & n1170;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n3012 & n3015;
  assign n3017 = ~n3011 & n3016;
  assign n1487_1 = ~n3010 | ~n3017;
  assign n3019 = n1184 & n1525;
  assign n3020 = Pkey_222_ & n1170;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = n1531 & ~n2756;
  assign n3023 = n1533 & n2758;
  assign n3024 = n1182 & ~n1525;
  assign n3025 = Pkey_230_ & n1145;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = ~n3023 & n3026;
  assign n3028 = ~n3022 & n3027;
  assign n1491_1 = ~n3021 | ~n3028;
  assign n3030 = n1184 & n1539;
  assign n3031 = Pkey_238_ & n1145;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = n1545 & ~n2756;
  assign n3034 = n1547 & n2758;
  assign n3035 = n1182 & ~n1539;
  assign n3036 = Pkey_230_ & n1170;
  assign n3037 = ~n3035 & ~n3036;
  assign n3038 = ~n3034 & n3037;
  assign n3039 = ~n3033 & n3038;
  assign n1496_1 = ~n3032 | ~n3039;
  assign n3041 = n1184 & n1553;
  assign n3042 = Pkey_238_ & n1170;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = n1559 & ~n2756;
  assign n3045 = n1561 & n2758;
  assign n3046 = n1182 & ~n1553;
  assign n3047 = Pkey_246_ & n1145;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = ~n3045 & n3048;
  assign n3050 = ~n3044 & n3049;
  assign n1500_1 = ~n3043 | ~n3050;
  assign n3052 = n1184 & n1567;
  assign n3053 = Pkey_254_ & n1145;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = n1573 & ~n2756;
  assign n3056 = n1575 & n2758;
  assign n3057 = n1182 & ~n1567;
  assign n3058 = Pkey_246_ & n1170;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3056 & n3059;
  assign n3061 = ~n3055 & n3060;
  assign n1504_1 = ~n3054 | ~n3061;
  assign n3063 = n1184 & n1581;
  assign n3064 = Pkey_254_ & n1170;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n1587 & ~n2756;
  assign n3067 = n1589 & n2758;
  assign n3068 = n1182 & ~n1581;
  assign n3069 = Pkey_131_ & n1145;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3067 & n3070;
  assign n3072 = ~n3066 & n3071;
  assign n1508_1 = ~n3065 | ~n3072;
  assign n3074 = n1184 & n1595;
  assign n3075 = Pkey_131_ & n1170;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n1601 & ~n2756;
  assign n3078 = n1603 & n2758;
  assign n3079 = n1182 & ~n1595;
  assign n3080 = Pkey_139_ & n1145;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = ~n3078 & n3081;
  assign n3083 = ~n3077 & n3082;
  assign n1512_1 = ~n3076 | ~n3083;
  assign n3085 = n1184 & n1609;
  assign n3086 = Pkey_147_ & n1145;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n1615 & ~n2756;
  assign n3089 = n1617 & n2758;
  assign n3090 = n1182 & ~n1609;
  assign n3091 = Pkey_139_ & n1170;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = ~n3089 & n3092;
  assign n3094 = ~n3088 & n3093;
  assign n1516_1 = ~n3087 | ~n3094;
  assign n3096 = n1184 & n1623;
  assign n3097 = Pkey_155_ & n1145;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n1629 & ~n2756;
  assign n3100 = n1631 & n2758;
  assign n3101 = n1182 & ~n1623;
  assign n3102 = Pkey_147_ & n1170;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n3100 & n3103;
  assign n3105 = ~n3099 & n3104;
  assign n1521_1 = ~n3098 | ~n3105;
  assign n3107 = n1184 & n1637;
  assign n3108 = Pkey_132_ & n1145;
  assign n3109 = ~n3107 & ~n3108;
  assign n3110 = n1643 & ~n2756;
  assign n3111 = n1645 & n2758;
  assign n3112 = n1182 & ~n1637;
  assign n3113 = Pkey_155_ & n1170;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~n3111 & n3114;
  assign n3116 = ~n3110 & n3115;
  assign n1525_1 = ~n3109 | ~n3116;
  assign n3118 = n1184 & n1651;
  assign n3119 = Pkey_132_ & n1170;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = n1657 & ~n2756;
  assign n3122 = n1659 & n2758;
  assign n3123 = n1182 & ~n1651;
  assign n3124 = Pkey_140_ & n1145;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3122 & n3125;
  assign n3127 = ~n3121 & n3126;
  assign n1529_1 = ~n3120 | ~n3127;
  assign n3129 = n1184 & n1665;
  assign n3130 = Pkey_140_ & n1170;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = n1671 & ~n2756;
  assign n3133 = n1673 & n2758;
  assign n3134 = n1182 & ~n1665;
  assign n3135 = Pkey_148_ & n1145;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3133 & n3136;
  assign n3138 = ~n3132 & n3137;
  assign n1533_1 = ~n3131 | ~n3138;
  assign n3140 = n1184 & n1678;
  assign n3141 = Pkey_148_ & n1170;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = n1681 & ~n2756;
  assign n3144 = n1687 & n2758;
  assign n3145 = n1182 & ~n1678;
  assign n3146 = Pkey_156_ & n1145;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = ~n3144 & n3147;
  assign n3149 = ~n3143 & n3148;
  assign n1537_1 = ~n3142 | ~n3149;
  assign n3151 = n1184 & n1692;
  assign n3152 = Pkey_156_ & n1170;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = n1691 & ~n2756;
  assign n3155 = n1693 & n2758;
  assign n3156 = n1182 & ~n1692;
  assign n3157 = Pkey_164_ & n1145;
  assign n3158 = ~n3156 & ~n3157;
  assign n3159 = ~n3155 & n3158;
  assign n3160 = ~n3154 & n3159;
  assign n1541_1 = ~n3153 | ~n3160;
  assign n3162 = n1184 & n1707;
  assign n3163 = ~n2860 & ~n3162;
  assign n3164 = n1713 & ~n2756;
  assign n3165 = n1715 & n2758;
  assign n3166 = n1182 & ~n1707;
  assign n3167 = Pkey_164_ & n1170;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = ~n3165 & n3168;
  assign n3170 = ~n3164 & n3169;
  assign n1545_1 = ~n3163 | ~n3170;
  assign n3172 = n1719 & ~n2756;
  assign n3173 = ~n1719 & n2758;
  assign n3174 = ~n1182 & ~n3173;
  assign n3175 = ~n1721 & ~n3174;
  assign n3176 = n1184 & n1721;
  assign n3177 = Pkey_180_ & n1145;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n2870 & n3178;
  assign n3180 = ~n3175 & n3179;
  assign n1549_1 = n3172 | ~n3180;
  assign n3182 = n1184 & n1734;
  assign n3183 = Pkey_188_ & n1145;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = n1740 & ~n2756;
  assign n3186 = n1742_1 & n2758;
  assign n3187 = n1182 & ~n1734;
  assign n3188 = Pkey_180_ & n1170;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = ~n3186 & n3189;
  assign n3191 = ~n3185 & n3190;
  assign n1553_1 = ~n3184 | ~n3191;
  assign n3193 = n1184 & n1748;
  assign n3194 = Pkey_133_ & n1145;
  assign n3195 = ~n3193 & ~n3194;
  assign n3196 = n1754 & ~n2756;
  assign n3197 = n1756 & n2758;
  assign n3198 = n1182 & ~n1748;
  assign n3199 = Pkey_188_ & n1170;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = ~n3197 & n3200;
  assign n3202 = ~n3196 & n3201;
  assign n1558_1 = ~n3195 | ~n3202;
  assign n3204 = n1184 & n1762;
  assign n3205 = Pkey_141_ & n1145;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = n1768 & ~n2756;
  assign n3208 = n1770 & n2758;
  assign n3209 = n1182 & ~n1762;
  assign n3210 = Pkey_133_ & n1170;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = ~n3208 & n3211;
  assign n3213 = ~n3207 & n3212;
  assign n1562_1 = ~n3206 | ~n3213;
  assign n3215 = n1184 & n1776;
  assign n3216 = Pkey_149_ & n1145;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = n1782 & ~n2756;
  assign n3219 = n1784 & n2758;
  assign n3220 = n1182 & ~n1776;
  assign n3221 = Pkey_141_ & n1170;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~n3219 & n3222;
  assign n3224 = ~n3218 & n3223;
  assign n1566_1 = ~n3217 | ~n3224;
  assign n3226 = n1184 & n1790;
  assign n3227 = Pkey_157_ & n1145;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = n1796 & ~n2756;
  assign n3230 = n1798 & n2758;
  assign n3231 = n1182 & ~n1790;
  assign n3232 = Pkey_149_ & n1170;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = ~n3230 & n3233;
  assign n3235 = ~n3229 & n3234;
  assign n1570_1 = ~n3228 | ~n3235;
  assign n3237 = n1184 & n1804;
  assign n3238 = Pkey_157_ & n1170;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = n1810 & ~n2756;
  assign n3241 = n1812 & n2758;
  assign n3242 = n1182 & ~n1804;
  assign n3243 = Pkey_165_ & n1145;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = ~n3241 & n3244;
  assign n3246 = ~n3240 & n3245;
  assign n1574_1 = ~n3239 | ~n3246;
  assign n3248 = n1184 & n1818;
  assign n3249 = Pkey_173_ & n1145;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = n1824 & ~n2756;
  assign n3252 = n1826 & n2758;
  assign n3253 = n1182 & ~n1818;
  assign n3254 = Pkey_165_ & n1170;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3252 & n3255;
  assign n3257 = ~n3251 & n3256;
  assign n1578_1 = ~n3250 | ~n3257;
  assign n3259 = n1184 & n1831;
  assign n3260 = Pkey_173_ & n1170;
  assign n3261 = ~n3259 & ~n3260;
  assign n3262 = n1830 & ~n2756;
  assign n3263 = n1832 & n2758;
  assign n3264 = n1182 & ~n1831;
  assign n3265 = Pkey_181_ & n1145;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~n3263 & n3266;
  assign n3268 = ~n3262 & n3267;
  assign n1582_1 = ~n3261 | ~n3268;
  assign n3270 = n1184 & n1846;
  assign n3271 = Pkey_189_ & n1145;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = n1852 & ~n2756;
  assign n3274 = n1854 & n2758;
  assign n3275 = n1182 & ~n1846;
  assign n3276 = Pkey_181_ & n1170;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = ~n3274 & n3277;
  assign n3279 = ~n3273 & n3278;
  assign n1587_1 = ~n3272 | ~n3279;
  assign n3281 = n1184 & n1860;
  assign n3282 = Pkey_189_ & n1170;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = n1866 & ~n2756;
  assign n3285 = n1868 & n2758;
  assign n3286 = n1182 & ~n1860;
  assign n3287 = Pkey_134_ & n1145;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = ~n3285 & n3288;
  assign n3290 = ~n3284 & n3289;
  assign n1591_1 = ~n3283 | ~n3290;
  assign n3292 = n1184 & n1874;
  assign n3293 = Pkey_134_ & n1170;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = n1880 & ~n2756;
  assign n3296 = n1882 & n2758;
  assign n3297 = n1182 & ~n1874;
  assign n3298 = Pkey_142_ & n1145;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~n3296 & n3299;
  assign n3301 = ~n3295 & n3300;
  assign n1595_1 = ~n3294 | ~n3301;
  assign n3303 = n1184 & n1888;
  assign n3304 = Pkey_142_ & n1170;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = n1894 & ~n2756;
  assign n3307 = n1896 & n2758;
  assign n3308 = n1182 & ~n1888;
  assign n3309 = Pkey_150_ & n1145;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = ~n3307 & n3310;
  assign n3312 = ~n3306 & n3311;
  assign n1600_1 = ~n3305 | ~n3312;
  assign n3314 = n1184 & n1902;
  assign n3315 = Pkey_150_ & n1170;
  assign n3316 = ~n3314 & ~n3315;
  assign n3317 = n1908 & ~n2756;
  assign n3318 = n1910 & n2758;
  assign n3319 = n1182 & ~n1902;
  assign n3320 = Pkey_158_ & n1145;
  assign n3321 = ~n3319 & ~n3320;
  assign n3322 = ~n3318 & n3321;
  assign n3323 = ~n3317 & n3322;
  assign n1604_1 = ~n3316 | ~n3323;
  assign n3325 = n1184 & n1916;
  assign n3326 = Pkey_158_ & n1170;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = n1922 & ~n2756;
  assign n3329 = n1924 & n2758;
  assign n3330 = n1182 & ~n1916;
  assign n3331 = Pkey_166_ & n1145;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = ~n3329 & n3332;
  assign n3334 = ~n3328 & n3333;
  assign n1608_1 = ~n3327 | ~n3334;
  assign n3336 = n1184 & n1930;
  assign n3337 = Pkey_174_ & n1145;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = n1936 & ~n2756;
  assign n3340 = n1938 & n2758;
  assign n3341 = n1182 & ~n1930;
  assign n3342 = Pkey_166_ & n1170;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3340 & n3343;
  assign n3345 = ~n3339 & n3344;
  assign n1612_1 = ~n3338 | ~n3345;
  assign n3347 = n1184 & n1944;
  assign n3348 = Pkey_182_ & n1145;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = n1950 & ~n2756;
  assign n3351 = n1952 & n2758;
  assign n3352 = n1182 & ~n1944;
  assign n3353 = Pkey_174_ & n1170;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = ~n3351 & n3354;
  assign n3356 = ~n3350 & n3355;
  assign n1616_1 = ~n3349 | ~n3356;
  assign n3358 = n1184 & n1958;
  assign n3359 = Pkey_182_ & n1170;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = n1964 & ~n2756;
  assign n3362 = n1966 & n2758;
  assign n3363 = n1182 & ~n1958;
  assign n3364 = Pkey_190_ & n1145;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = ~n3362 & n3365;
  assign n3367 = ~n3361 & n3366;
  assign n1620_1 = ~n3360 | ~n3367;
  assign n3369 = n1184 & n1972;
  assign n3370 = Pkey_190_ & n1170;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = n1978 & ~n2756;
  assign n3373 = n1980 & n2758;
  assign n3374 = n1182 & ~n1972;
  assign n3375 = Pkey_67_ & n1145;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = ~n3373 & n3376;
  assign n3378 = ~n3372 & n3377;
  assign n1624_1 = ~n3371 | ~n3378;
  assign n3380 = n1184 & n1986;
  assign n3381 = Pkey_75_ & n1145;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = n1992 & ~n2756;
  assign n3384 = n1994 & n2758;
  assign n3385 = n1182 & ~n1986;
  assign n3386 = Pkey_67_ & n1170;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n3384 & n3387;
  assign n3389 = ~n3383 & n3388;
  assign n1628_1 = ~n3382 | ~n3389;
  assign n3391 = n1184 & n2000;
  assign n3392 = Pkey_75_ & n1170;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = n2006 & ~n2756;
  assign n3395 = n2008 & n2758;
  assign n3396 = n1182 & ~n2000;
  assign n3397 = Pkey_83_ & n1145;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n3395 & n3398;
  assign n3400 = ~n3394 & n3399;
  assign n1632_1 = ~n3393 | ~n3400;
  assign n3402 = n1184 & n2014;
  assign n3403 = Pkey_91_ & n1145;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n2020 & ~n2756;
  assign n3406 = n2022 & n2758;
  assign n3407 = n1182 & ~n2014;
  assign n3408 = Pkey_83_ & n1170;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~n3406 & n3409;
  assign n3411 = ~n3405 & n3410;
  assign n1637_1 = ~n3404 | ~n3411;
  assign n3413 = n1184 & n2028;
  assign n3414 = Pkey_68_ & n1145;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = n2034 & ~n2756;
  assign n3417 = n2036 & n2758;
  assign n3418 = n1182 & ~n2028;
  assign n3419 = Pkey_91_ & n1170;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = ~n3417 & n3420;
  assign n3422 = ~n3416 & n3421;
  assign n1641_1 = ~n3415 | ~n3422;
  assign n3424 = n1184 & n2042;
  assign n3425 = Pkey_76_ & n1145;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = n2048 & ~n2756;
  assign n3428 = n2050 & n2758;
  assign n3429 = n1182 & ~n2042;
  assign n3430 = Pkey_68_ & n1170;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = ~n3428 & n3431;
  assign n3433 = ~n3427 & n3432;
  assign n1645_1 = ~n3426 | ~n3433;
  assign n3435 = n1184 & n2055;
  assign n3436 = Pkey_84_ & n1145;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = n2054 & ~n2756;
  assign n3439 = n2056 & n2758;
  assign n3440 = n1182 & ~n2055;
  assign n3441 = Pkey_76_ & n1170;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = ~n3439 & n3442;
  assign n3444 = ~n3438 & n3443;
  assign n1649_1 = ~n3437 | ~n3444;
  assign n3446 = n1184 & n2070;
  assign n3447 = Pkey_92_ & n1145;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = n2076 & ~n2756;
  assign n3450 = n2078 & n2758;
  assign n3451 = n1182 & ~n2070;
  assign n3452 = Pkey_84_ & n1170;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = ~n3450 & n3453;
  assign n3455 = ~n3449 & n3454;
  assign n1653_1 = ~n3448 | ~n3455;
  assign n3457 = n1184 & n2084;
  assign n3458 = Pkey_92_ & n1170;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = n2090 & ~n2756;
  assign n3461 = n2092 & n2758;
  assign n3462 = n1182 & ~n2084;
  assign n3463 = Pkey_100_ & n1145;
  assign n3464 = ~n3462 & ~n3463;
  assign n3465 = ~n3461 & n3464;
  assign n3466 = ~n3460 & n3465;
  assign n1657_1 = ~n3459 | ~n3466;
  assign n3468 = n1182 & ~n2098;
  assign n3469 = Pkey_100_ & n1170;
  assign n3470 = ~n3468 & ~n3469;
  assign n3471 = n2104 & ~n2756;
  assign n3472 = n2106 & n2758;
  assign n3473 = n1184 & n2098;
  assign n3474 = Pkey_44_ & n1145;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = ~n3472 & n3475;
  assign n3477 = ~n3471 & n3476;
  assign n1661_1 = ~n3470 | ~n3477;
  assign n3479 = n1182 & ~n2112;
  assign n3480 = Pkey_44_ & n1170;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = n2118 & ~n2756;
  assign n3483 = n2120 & n2758;
  assign n3484 = n1184 & n2112;
  assign n3485 = Pkey_116_ & n1145;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = ~n3483 & n3486;
  assign n3488 = ~n3482 & n3487;
  assign n1665_1 = ~n3481 | ~n3488;
  assign n3490 = n1184 & n2126;
  assign n3491 = Pkey_124_ & n1145;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = n2124 & ~n2756;
  assign n3494 = n2127 & n2758;
  assign n3495 = n1182 & ~n2126;
  assign n3496 = Pkey_116_ & n1170;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = ~n3494 & n3497;
  assign n3499 = ~n3493 & n3498;
  assign n1669_1 = ~n3492 | ~n3499;
  assign n3501 = n1184 & n2140;
  assign n3502 = Pkey_124_ & n1170;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = n2146 & ~n2756;
  assign n3505 = n2148 & n2758;
  assign n3506 = n1182 & ~n2140;
  assign n3507 = Pkey_69_ & n1145;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3505 & n3508;
  assign n3510 = ~n3504 & n3509;
  assign n1673_1 = ~n3503 | ~n3510;
  assign n3512 = n1184 & n2154;
  assign n3513 = Pkey_69_ & n1170;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n2160 & ~n2756;
  assign n3516 = n2162 & n2758;
  assign n3517 = n1182 & ~n2154;
  assign n3518 = Pkey_77_ & n1145;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3516 & n3519;
  assign n3521 = ~n3515 & n3520;
  assign n1677_1 = ~n3514 | ~n3521;
  assign n3523 = n1184 & n2168;
  assign n3524 = Pkey_85_ & n1145;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = n2174 & ~n2756;
  assign n3527 = n2176 & n2758;
  assign n3528 = n1182 & ~n2168;
  assign n3529 = Pkey_77_ & n1170;
  assign n3530 = ~n3528 & ~n3529;
  assign n3531 = ~n3527 & n3530;
  assign n3532 = ~n3526 & n3531;
  assign n1682_1 = ~n3525 | ~n3532;
  assign n3534 = n1184 & n2182;
  assign n3535 = Pkey_85_ & n1170;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = n2188 & ~n2756;
  assign n3538 = n2190 & n2758;
  assign n3539 = n1182 & ~n2182;
  assign n3540 = Pkey_93_ & n1145;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = ~n3538 & n3541;
  assign n3543 = ~n3537 & n3542;
  assign n1687_1 = ~n3536 | ~n3543;
  assign n3545 = n1184 & n2196;
  assign n3546 = Pkey_101_ & n1145;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = n2202 & ~n2756;
  assign n3549 = n2204 & n2758;
  assign n3550 = n1182 & ~n2196;
  assign n3551 = Pkey_93_ & n1170;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = ~n3549 & n3552;
  assign n3554 = ~n3548 & n3553;
  assign n1691_1 = ~n3547 | ~n3554;
  assign n3556 = n1184 & n2210;
  assign n3557 = Pkey_101_ & n1170;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = n2216 & ~n2756;
  assign n3560 = n2218 & n2758;
  assign n3561 = n1182 & ~n2210;
  assign n3562 = Pkey_109_ & n1145;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n3560 & n3563;
  assign n3565 = ~n3559 & n3564;
  assign n1695_1 = ~n3558 | ~n3565;
  assign n3567 = n1184 & n2224;
  assign n3568 = Pkey_109_ & n1170;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = n2230 & ~n2756;
  assign n3571 = n2232 & n2758;
  assign n3572 = n1182 & ~n2224;
  assign n3573 = Pkey_117_ & n1145;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575 = ~n3571 & n3574;
  assign n3576 = ~n3570 & n3575;
  assign n1699_1 = ~n3569 | ~n3576;
  assign n3578 = n1184 & n2238;
  assign n3579 = Pkey_117_ & n1170;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = n2244 & ~n2756;
  assign n3582 = n2246 & n2758;
  assign n3583 = n1182 & ~n2238;
  assign n3584 = Pkey_125_ & n1145;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = ~n3582 & n3585;
  assign n3587 = ~n3581 & n3586;
  assign n1704_1 = ~n3580 | ~n3587;
  assign n3589 = n1184 & n2252;
  assign n3590 = Pkey_125_ & n1170;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = n2258 & ~n2756;
  assign n3593 = n2260 & n2758;
  assign n3594 = n1182 & ~n2252;
  assign n3595 = Pkey_70_ & n1145;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3593 & n3596;
  assign n3598 = ~n3592 & n3597;
  assign n1708_1 = ~n3591 | ~n3598;
  assign n3600 = n1184 & n2266;
  assign n3601 = Pkey_78_ & n1145;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = n2272 & ~n2756;
  assign n3604 = n2274 & n2758;
  assign n3605 = n1182 & ~n2266;
  assign n3606 = Pkey_70_ & n1170;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n3604 & n3607;
  assign n3609 = ~n3603 & n3608;
  assign n1712_1 = ~n3602 | ~n3609;
  assign n3611 = n1184 & n2279;
  assign n3612 = Pkey_86_ & n1145;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = n2278 & ~n2756;
  assign n3615 = n2280 & n2758;
  assign n3616 = n1182 & ~n2279;
  assign n3617 = Pkey_78_ & n1170;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = ~n3615 & n3618;
  assign n3620 = ~n3614 & n3619;
  assign n1717_1 = ~n3613 | ~n3620;
  assign n3622 = n1184 & n2294;
  assign n3623 = Pkey_86_ & n1170;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = n2292 & ~n2756;
  assign n3626 = n2295 & n2758;
  assign n3627 = n1182 & ~n2294;
  assign n3628 = Pkey_94_ & n1145;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = ~n3626 & n3629;
  assign n3631 = ~n3625 & n3630;
  assign n1721_1 = ~n3624 | ~n3631;
  assign n3633 = n1184 & n2308;
  assign n3634 = Pkey_94_ & n1170;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = n2314 & ~n2756;
  assign n3637 = n2316 & n2758;
  assign n3638 = n1182 & ~n2308;
  assign n3639 = Pkey_102_ & n1145;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~n3637 & n3640;
  assign n3642 = ~n3636 & n3641;
  assign n1725_1 = ~n3635 | ~n3642;
  assign n3644 = n1184 & n2322;
  assign n3645 = Pkey_110_ & n1145;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = n2328 & ~n2756;
  assign n3648 = n2330 & n2758;
  assign n3649 = n1182 & ~n2322;
  assign n3650 = Pkey_102_ & n1170;
  assign n3651 = ~n3649 & ~n3650;
  assign n3652 = ~n3648 & n3651;
  assign n3653 = ~n3647 & n3652;
  assign n1730_1 = ~n3646 | ~n3653;
  assign n3655 = n1184 & n2336;
  assign n3656 = Pkey_118_ & n1145;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = n2342 & ~n2756;
  assign n3659 = n2344 & n2758;
  assign n3660 = n1182 & ~n2336;
  assign n3661 = Pkey_110_ & n1170;
  assign n3662 = ~n3660 & ~n3661;
  assign n3663 = ~n3659 & n3662;
  assign n3664 = ~n3658 & n3663;
  assign n1734_1 = ~n3657 | ~n3664;
  assign n3666 = n1184 & n2350;
  assign n3667 = Pkey_126_ & n1145;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = n2356 & ~n2756;
  assign n3670 = n2358 & n2758;
  assign n3671 = n1182 & ~n2350;
  assign n3672 = Pkey_118_ & n1170;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = ~n3670 & n3673;
  assign n3675 = ~n3669 & n3674;
  assign n1738_1 = ~n3668 | ~n3675;
  assign n3677 = n1184 & n2364;
  assign n3678 = Pkey_126_ & n1170;
  assign n3679 = ~n3677 & ~n3678;
  assign n3680 = n2370 & ~n2756;
  assign n3681 = n2372 & n2758;
  assign n3682 = n1182 & ~n2364;
  assign n3683 = Pkey_3_ & n1145;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n3681 & n3684;
  assign n3686 = ~n3680 & n3685;
  assign n1742 = ~n3679 | ~n3686;
  assign n3688 = n1184 & n2378;
  assign n3689 = Pkey_11_ & n1145;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = n2384 & ~n2756;
  assign n3692 = n2386 & n2758;
  assign n3693 = n1182 & ~n2378;
  assign n3694 = Pkey_3_ & n1170;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = ~n3692 & n3695;
  assign n3697 = ~n3691 & n3696;
  assign n1746_1 = ~n3690 | ~n3697;
  assign n3699 = n1184 & n2392;
  assign n3700 = Pkey_19_ & n1145;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = n2398 & ~n2756;
  assign n3703 = n2400 & n2758;
  assign n3704 = n1182 & ~n2392;
  assign n3705 = Pkey_11_ & n1170;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = ~n3703 & n3706;
  assign n3708 = ~n3702 & n3707;
  assign n1750_1 = ~n3701 | ~n3708;
  assign n3710 = n1184 & n2406;
  assign n3711 = Pkey_19_ & n1170;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = n2412 & ~n2756;
  assign n3714 = n2414 & n2758;
  assign n3715 = n1182 & ~n2406;
  assign n3716 = Pkey_27_ & n1145;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = ~n3714 & n3717;
  assign n3719 = ~n3713 & n3718;
  assign n1755 = ~n3712 | ~n3719;
  assign n3721 = n1184 & n2420;
  assign n3722 = Pkey_4_ & n1145;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = n2426 & ~n2756;
  assign n3725 = n2428 & n2758;
  assign n3726 = n1182 & ~n2420;
  assign n3727 = Pkey_27_ & n1170;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n3725 & n3728;
  assign n3730 = ~n3724 & n3729;
  assign n1759 = ~n3723 | ~n3730;
  assign n3732 = n1184 & n2434;
  assign n3733 = Pkey_12_ & n1145;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = n2440 & ~n2756;
  assign n3736 = n2442 & n2758;
  assign n3737 = n1182 & ~n2434;
  assign n3738 = Pkey_4_ & n1170;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~n3736 & n3739;
  assign n3741 = ~n3735 & n3740;
  assign n1763 = ~n3734 | ~n3741;
  assign n3743 = n1184 & n2448;
  assign n3744 = Pkey_12_ & n1170;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = n2454 & ~n2756;
  assign n3747 = n2456 & n2758;
  assign n3748 = n1182 & ~n2448;
  assign n3749 = Pkey_20_ & n1145;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = ~n3747 & n3750;
  assign n3752 = ~n3746 & n3751;
  assign n1767 = ~n3745 | ~n3752;
  assign n3754 = n1184 & n2462;
  assign n3755 = Pkey_20_ & n1170;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = n2468 & ~n2756;
  assign n3758 = n2470 & n2758;
  assign n3759 = n1182 & ~n2462;
  assign n3760 = Pkey_28_ & n1145;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n3758 & n3761;
  assign n3763 = ~n3757 & n3762;
  assign n1771 = ~n3756 | ~n3763;
  assign n3765 = n1184 & n2476;
  assign n3766 = Pkey_28_ & n1170;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = n2482 & ~n2756;
  assign n3769 = n2484 & n2758;
  assign n3770 = n1182 & ~n2476;
  assign n3771 = Pkey_36_ & n1145;
  assign n3772 = ~n3770 & ~n3771;
  assign n3773 = ~n3769 & n3772;
  assign n3774 = ~n3768 & n3773;
  assign n1775 = ~n3767 | ~n3774;
  assign n3776 = n2488 & ~n2756;
  assign n3777 = ~n2488 & n2758;
  assign n3778 = ~n1182 & ~n3777;
  assign n3779 = ~n2490 & ~n3778;
  assign n3780 = Pkey_36_ & n1170;
  assign n3781 = n1184 & n2490;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~n3474 & n3782;
  assign n3784 = ~n3779 & n3783;
  assign n1779 = n3776 | ~n3784;
  assign n3786 = n1182 & ~n2503;
  assign n3787 = Pkey_52_ & n1145;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = n2509 & ~n2756;
  assign n3790 = n2511 & n2758;
  assign n3791 = n1184 & n2503;
  assign n3792 = ~n3480 & ~n3791;
  assign n3793 = ~n3790 & n3792;
  assign n3794 = ~n3789 & n3793;
  assign n1783 = ~n3788 | ~n3794;
  assign n3796 = n1184 & n2517;
  assign n3797 = Pkey_52_ & n1170;
  assign n3798 = ~n3796 & ~n3797;
  assign n3799 = n2523 & ~n2756;
  assign n3800 = n2525 & n2758;
  assign n3801 = n1182 & ~n2517;
  assign n3802 = Pkey_60_ & n1145;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = ~n3800 & n3803;
  assign n3805 = ~n3799 & n3804;
  assign n1787 = ~n3798 | ~n3805;
  assign n3807 = n1184 & n2531;
  assign n3808 = Pkey_5_ & n1145;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = n2537 & ~n2756;
  assign n3811 = n2539 & n2758;
  assign n3812 = n1182 & ~n2531;
  assign n3813 = Pkey_60_ & n1170;
  assign n3814 = ~n3812 & ~n3813;
  assign n3815 = ~n3811 & n3814;
  assign n3816 = ~n3810 & n3815;
  assign n1791 = ~n3809 | ~n3816;
  assign n3818 = n1184 & n2545;
  assign n3819 = Pkey_5_ & n1170;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = n2551 & ~n2756;
  assign n3822 = n2553 & n2758;
  assign n3823 = n1182 & ~n2545;
  assign n3824 = Pkey_13_ & n1145;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = ~n3822 & n3825;
  assign n3827 = ~n3821 & n3826;
  assign n1795 = ~n3820 | ~n3827;
  assign n3829 = n1184 & n2559;
  assign n3830 = Pkey_21_ & n1145;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n2565 & ~n2756;
  assign n3833 = n2567 & n2758;
  assign n3834 = n1182 & ~n2559;
  assign n3835 = Pkey_13_ & n1170;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3833 & n3836;
  assign n3838 = ~n3832 & n3837;
  assign n1800_1 = ~n3831 | ~n3838;
  assign n3840 = n1184 & n2573;
  assign n3841 = Pkey_29_ & n1145;
  assign n3842 = ~n3840 & ~n3841;
  assign n3843 = n2571 & ~n2756;
  assign n3844 = n2574 & n2758;
  assign n3845 = n1182 & ~n2573;
  assign n3846 = Pkey_21_ & n1170;
  assign n3847 = ~n3845 & ~n3846;
  assign n3848 = ~n3844 & n3847;
  assign n3849 = ~n3843 & n3848;
  assign n1804_1 = ~n3842 | ~n3849;
  assign n3851 = n1184 & n2587;
  assign n3852 = Pkey_37_ & n1145;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = n2593 & ~n2756;
  assign n3855 = n2595 & n2758;
  assign n3856 = n1182 & ~n2587;
  assign n3857 = Pkey_29_ & n1170;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = ~n3855 & n3858;
  assign n3860 = ~n3854 & n3859;
  assign n1808_1 = ~n3853 | ~n3860;
  assign n3862 = n1184 & n2601;
  assign n3863 = Pkey_37_ & n1170;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = n2607 & ~n2756;
  assign n3866 = n2609 & n2758;
  assign n3867 = n1182 & ~n2601;
  assign n3868 = Pkey_45_ & n1145;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3866 & n3869;
  assign n3871 = ~n3865 & n3870;
  assign n1812_1 = ~n3864 | ~n3871;
  assign n3873 = n1184 & n2615;
  assign n3874 = Pkey_53_ & n1145;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = n2621 & ~n2756;
  assign n3877 = n2623 & n2758;
  assign n3878 = n1182 & ~n2615;
  assign n3879 = Pkey_45_ & n1170;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = ~n3877 & n3880;
  assign n3882 = ~n3876 & n3881;
  assign n1816_1 = ~n3875 | ~n3882;
  assign n3884 = n1184 & n2629;
  assign n3885 = Pkey_61_ & n1145;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = n2635 & ~n2756;
  assign n3888 = n2637 & n2758;
  assign n3889 = n1182 & ~n2629;
  assign n3890 = Pkey_53_ & n1170;
  assign n3891 = ~n3889 & ~n3890;
  assign n3892 = ~n3888 & n3891;
  assign n3893 = ~n3887 & n3892;
  assign n1821 = ~n3886 | ~n3893;
  assign n3895 = n1184 & n2642;
  assign n3896 = Pkey_61_ & n1170;
  assign n3897 = ~n3895 & ~n3896;
  assign n3898 = n2641 & ~n2756;
  assign n3899 = n2643 & n2758;
  assign n3900 = n1182 & ~n2642;
  assign n3901 = Pkey_6_ & n1145;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = ~n3899 & n3902;
  assign n3904 = ~n3898 & n3903;
  assign n1825 = ~n3897 | ~n3904;
  assign n3906 = n1184 & n2657;
  assign n3907 = Pkey_6_ & n1170;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = n2663 & ~n2756;
  assign n3910 = n2665 & n2758;
  assign n3911 = n1182 & ~n2657;
  assign n3912 = Pkey_14_ & n1145;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = ~n3910 & n3913;
  assign n3915 = ~n3909 & n3914;
  assign n1829 = ~n3908 | ~n3915;
  assign n3917 = n1184 & n2671;
  assign n3918 = Pkey_14_ & n1170;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = n2677 & ~n2756;
  assign n3921 = n2679 & n2758;
  assign n3922 = n1182 & ~n2671;
  assign n3923 = Pkey_22_ & n1145;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n3921 & n3924;
  assign n3926 = ~n3920 & n3925;
  assign n1834_1 = ~n3919 | ~n3926;
  assign n3928 = n1184 & n2685;
  assign n3929 = Pkey_22_ & n1170;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n2691 & ~n2756;
  assign n3932 = n2693 & n2758;
  assign n3933 = n1182 & ~n2685;
  assign n3934 = Pkey_30_ & n1145;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = ~n3932 & n3935;
  assign n3937 = ~n3931 & n3936;
  assign n1838_1 = ~n3930 | ~n3937;
  assign n3939 = n1184 & n2699;
  assign n3940 = Pkey_30_ & n1170;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = n2705 & ~n2756;
  assign n3943 = n2707 & n2758;
  assign n3944 = n1182 & ~n2699;
  assign n3945 = Pkey_38_ & n1145;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = ~n3943 & n3946;
  assign n3948 = ~n3942 & n3947;
  assign n1842_1 = ~n3941 | ~n3948;
  assign n3950 = n1184 & n2713;
  assign n3951 = Pkey_46_ & n1145;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = n2711 & ~n2756;
  assign n3954 = n2714 & n2758;
  assign n3955 = n1182 & ~n2713;
  assign n3956 = Pkey_38_ & n1170;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3954 & n3957;
  assign n3959 = ~n3953 & n3958;
  assign n1846_1 = ~n3952 | ~n3959;
  assign n3961 = n1184 & n2727;
  assign n3962 = Pkey_54_ & n1145;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = n2733 & ~n2756;
  assign n3965 = n2735 & n2758;
  assign n3966 = n1182 & ~n2727;
  assign n3967 = Pkey_46_ & n1170;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = ~n3965 & n3968;
  assign n3970 = ~n3964 & n3969;
  assign n1850_1 = ~n3963 | ~n3970;
  assign n3972 = n1184 & n2741;
  assign n3973 = Pkey_54_ & n1170;
  assign n3974 = ~n3972 & ~n3973;
  assign n3975 = n2747 & ~n2756;
  assign n3976 = n2749 & n2758;
  assign n3977 = n1182 & ~n2741;
  assign n3978 = Pkey_62_ & n1145;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = ~n3976 & n3979;
  assign n3981 = ~n3975 & n3980;
  assign n1854_1 = ~n3974 | ~n3981;
  assign PKSi_191_ = \[234] ;
  assign PKSi_187_ = \[234] ;
  assign PKSi_181_ = \[253] ;
  assign PKSi_168_ = \[253] ;
  assign PKSi_143_ = \[282] ;
  assign PKSi_139_ = \[282] ;
  assign PKSi_90_ = \[333] ;
  assign PKSi_88_ = \[333] ;
  always @ (posedge clock) begin
    PKSi_79_ <= n922_1;
    PKSi_92_ <= n926;
    \[333]  <= n930_1;
    N_N2737 <= n935_1;
    PKSi_75_ <= n940_1;
    PKSi_84_ <= n944_1;
    N_N2741 <= n948_1;
    PKSi_82_ <= n953;
    PKSi_93_ <= n957;
    PKSi_85_ <= n961;
    N_N2746 <= n965;
    PKSi_73_ <= n970_1;
    N_N2749 <= n974_1;
    PKSi_80_ <= n979;
    PKSi_72_ <= n983;
    PKSi_94_ <= n987;
    PKSi_86_ <= n991;
    PKSi_74_ <= n995;
    PKSi_83_ <= n999;
    N_N2757 <= n1003;
    PKSi_89_ <= n1008_1;
    PKSi_91_ <= n1012_1;
    PKSi_81_ <= n1016_1;
    PKSi_77_ <= n1020_1;
    PKSi_87_ <= n1024_1;
    PKSi_78_ <= n1028_1;
    PKSi_95_ <= n1032_1;
    PKSi_76_ <= n1036_1;
    PKSi_55_ <= n1040_1;
    PKSi_68_ <= n1044_1;
    PKSi_64_ <= n1048_1;
    N_N2770 <= n1052_1;
    PKSi_51_ <= n1057;
    PKSi_60_ <= n1061;
    N_N2774 <= n1065;
    PKSi_58_ <= n1070_1;
    PKSi_69_ <= n1074_1;
    PKSi_61_ <= n1078_1;
    N_N2779 <= n1082_1;
    PKSi_49_ <= n1087;
    PKSi_66_ <= n1091;
    PKSi_56_ <= n1095;
    PKSi_48_ <= n1099;
    PKSi_70_ <= n1103;
    PKSi_62_ <= n1107;
    PKSi_50_ <= n1111;
    PKSi_59_ <= n1115;
    N_N2789 <= n1119;
    PKSi_65_ <= n1124_1;
    PKSi_67_ <= n1128_1;
    PKSi_57_ <= n1132_1;
    PKSi_53_ <= n1136_1;
    PKSi_63_ <= n1140_1;
    PKSi_54_ <= n1144_1;
    PKSi_71_ <= n1148_1;
    PKSi_52_ <= n1152_1;
    PKSi_31_ <= n1156_1;
    PKSi_44_ <= n1160_1;
    PKSi_40_ <= n1164;
    N_N2802 <= n1168;
    PKSi_27_ <= n1173;
    PKSi_36_ <= n1177;
    N_N2806 <= n1181;
    PKSi_34_ <= n1186;
    PKSi_45_ <= n1190;
    PKSi_37_ <= n1194;
    N_N2811 <= n1198;
    PKSi_25_ <= n1203;
    PKSi_42_ <= n1207;
    PKSi_32_ <= n1211;
    PKSi_24_ <= n1215;
    PKSi_46_ <= n1219;
    PKSi_38_ <= n1223;
    PKSi_26_ <= n1227;
    PKSi_35_ <= n1231;
    N_N2821 <= n1235;
    PKSi_41_ <= n1240;
    PKSi_43_ <= n1244;
    PKSi_33_ <= n1248;
    PKSi_29_ <= n1252;
    PKSi_39_ <= n1256;
    PKSi_30_ <= n1260;
    PKSi_47_ <= n1264;
    PKSi_28_ <= n1268;
    PKSi_7_ <= n1272;
    PKSi_20_ <= n1276;
    PKSi_16_ <= n1280;
    N_N2834 <= n1284_1;
    PKSi_3_ <= n1289_1;
    PKSi_12_ <= n1293_1;
    N_N2838 <= n1297_1;
    PKSi_10_ <= n1302_1;
    PKSi_21_ <= n1306_1;
    PKSi_13_ <= n1310_1;
    N_N2843 <= n1314_1;
    PKSi_1_ <= n1319_1;
    PKSi_18_ <= n1323_1;
    PKSi_8_ <= n1327_1;
    PKSi_0_ <= n1331_1;
    PKSi_22_ <= n1335_1;
    PKSi_14_ <= n1339_1;
    PKSi_2_ <= n1343_1;
    PKSi_11_ <= n1347_1;
    N_N2853 <= n1351_1;
    PKSi_17_ <= n1356_1;
    PKSi_19_ <= n1360_1;
    PKSi_9_ <= n1364_1;
    PKSi_5_ <= n1368_1;
    PKSi_15_ <= n1372_1;
    PKSi_6_ <= n1376_1;
    PKSi_23_ <= n1380_1;
    PKSi_4_ <= n1384_1;
    PKSi_183_ <= n1388_1;
    PKSi_173_ <= n1392_1;
    N_N2865 <= n1396_1;
    PKSi_185_ <= n1401_1;
    PKSi_169_ <= n1405_1;
    PKSi_176_ <= n1409_1;
    PKSi_188_ <= n1413_1;
    \[253]  <= n1417_1;
    PKSi_179_ <= n1422_1;
    PKSi_172_ <= n1426_1;
    PKSi_186_ <= n1430_1;
    PKSi_177_ <= n1434_1;
    PKSi_180_ <= n1438_1;
    N_N2877 <= n1442_1;
    N_N2879 <= n1447_1;
    N_N2881 <= n1452_1;
    PKSi_175_ <= n1457_1;
    PKSi_182_ <= n1461_1;
    N_N2885 <= n1465_1;
    PKSi_171_ <= n1470_1;
    PKSi_189_ <= n1474_1;
    N_N2889 <= n1478_1;
    PKSi_184_ <= n1483_1;
    PKSi_178_ <= n1487_1;
    \[234]  <= n1491_1;
    PKSi_170_ <= n1496_1;
    PKSi_174_ <= n1500_1;
    PKSi_190_ <= n1504_1;
    PKSi_159_ <= n1508_1;
    PKSi_149_ <= n1512_1;
    N_N2899 <= n1516_1;
    PKSi_161_ <= n1521_1;
    PKSi_145_ <= n1525_1;
    PKSi_152_ <= n1529_1;
    PKSi_164_ <= n1533_1;
    PKSi_157_ <= n1537_1;
    PKSi_155_ <= n1541_1;
    PKSi_148_ <= n1545_1;
    PKSi_162_ <= n1549_1;
    N_N2909 <= n1553_1;
    PKSi_156_ <= n1558_1;
    PKSi_153_ <= n1562_1;
    PKSi_163_ <= n1566_1;
    PKSi_144_ <= n1570_1;
    PKSi_151_ <= n1574_1;
    PKSi_158_ <= n1578_1;
    N_N2917 <= n1582_1;
    PKSi_147_ <= n1587_1;
    PKSi_165_ <= n1591_1;
    N_N2921 <= n1595_1;
    PKSi_160_ <= n1600_1;
    PKSi_154_ <= n1604_1;
    PKSi_167_ <= n1608_1;
    PKSi_146_ <= n1612_1;
    PKSi_150_ <= n1616_1;
    PKSi_166_ <= n1620_1;
    PKSi_135_ <= n1624_1;
    PKSi_125_ <= n1628_1;
    N_N2931 <= n1632_1;
    PKSi_137_ <= n1637_1;
    PKSi_121_ <= n1641_1;
    PKSi_128_ <= n1645_1;
    PKSi_140_ <= n1649_1;
    PKSi_133_ <= n1653_1;
    PKSi_131_ <= n1657_1;
    PKSi_124_ <= n1661_1;
    PKSi_138_ <= n1665_1;
    PKSi_129_ <= n1669_1;
    PKSi_132_ <= n1673_1;
    N_N2943 <= n1677_1;
    N_N2945 <= n1682_1;
    PKSi_120_ <= n1687_1;
    PKSi_127_ <= n1691_1;
    PKSi_134_ <= n1695_1;
    N_N2950 <= n1699_1;
    PKSi_123_ <= n1704_1;
    PKSi_141_ <= n1708_1;
    N_N2954 <= n1712_1;
    PKSi_136_ <= n1717_1;
    PKSi_130_ <= n1721_1;
    \[282]  <= n1725_1;
    PKSi_122_ <= n1730_1;
    PKSi_126_ <= n1734_1;
    PKSi_142_ <= n1738_1;
    PKSi_111_ <= n1742;
    PKSi_101_ <= n1746_1;
    N_N2964 <= n1750_1;
    PKSi_113_ <= n1755;
    PKSi_97_ <= n1759;
    PKSi_104_ <= n1763;
    PKSi_116_ <= n1767;
    PKSi_109_ <= n1771;
    PKSi_107_ <= n1775;
    PKSi_100_ <= n1779;
    PKSi_114_ <= n1783;
    PKSi_105_ <= n1787;
    PKSi_108_ <= n1791;
    N_N2976 <= n1795;
    PKSi_115_ <= n1800_1;
    PKSi_96_ <= n1804_1;
    PKSi_103_ <= n1808_1;
    PKSi_110_ <= n1812_1;
    N_N2982 <= n1816_1;
    PKSi_99_ <= n1821;
    PKSi_117_ <= n1825;
    N_N2986 <= n1829;
    PKSi_112_ <= n1834_1;
    PKSi_106_ <= n1838_1;
    PKSi_119_ <= n1842_1;
    PKSi_98_ <= n1846_1;
    PKSi_102_ <= n1850_1;
    PKSi_118_ <= n1854_1;
  end
endmodule


