// Benchmark "alu4" written by ABC on Sat Apr 23 20:18:09 2016

module alu4 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    z0, z1, z2, z3, z4, z5, z6, z7  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13;
  output z0, z1, z2, z3, z4, z5, z6, z7;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n46, n47, n48, n49, n50, n51,
    n52, n53, n54, n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66,
    n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925;
  assign n23 = ~x05 & ~x10;
  assign n24 = x00 & ~n23;
  assign n25 = x03 & x08;
  assign n26 = x03 & x10;
  assign n27 = ~n25 & ~n26;
  assign n28 = ~x06 & ~x10;
  assign n29 = x01 & ~n28;
  assign n30 = x02 & x10;
  assign n31 = x02 & x07;
  assign n32 = ~n30 & ~n31;
  assign n33 = ~n29 & n32;
  assign n34 = n27 & n33;
  assign n35 = ~n24 & n34;
  assign n36 = x09 & ~n35;
  assign n37 = x01 & ~x06;
  assign n38 = x00 & ~x05;
  assign n39 = x03 & ~x08;
  assign n40 = x02 & ~x07;
  assign n41 = ~n39 & ~n40;
  assign n42 = ~n38 & n41;
  assign n43 = ~n37 & n42;
  assign n44 = x10 & ~n43;
  assign z0 = n36 | n44;
  assign n46 = x04 & ~x13;
  assign n47 = ~x08 & x10;
  assign n48 = x08 & x09;
  assign n49 = ~n47 & ~n48;
  assign n50 = x03 & n49;
  assign n51 = ~x08 & ~x11;
  assign n52 = x08 & ~x12;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~x03 & n53;
  assign n55 = ~n50 & ~n54;
  assign n56 = n46 & n55;
  assign n57 = ~n46 & ~n55;
  assign z1 = ~n56 & ~n57;
  assign n59 = ~x01 & ~x06;
  assign n60 = ~x11 & n59;
  assign n61 = x12 & ~n60;
  assign n62 = ~x05 & ~x07;
  assign n63 = ~x00 & ~x05;
  assign n64 = ~x02 & ~x07;
  assign n65 = ~x03 & ~x08;
  assign n66 = ~n64 & ~n65;
  assign n67 = ~n63 & n66;
  assign n68 = ~n62 & n67;
  assign n69 = x00 & x02;
  assign n70 = x08 & n69;
  assign n71 = ~n68 & ~n70;
  assign n72 = ~x11 & n71;
  assign n73 = n61 & ~n72;
  assign n74 = x06 & x12;
  assign n75 = x07 & x09;
  assign n76 = ~x07 & x10;
  assign n77 = ~n75 & ~n76;
  assign n78 = x02 & ~n77;
  assign n79 = x02 & x03;
  assign n80 = ~n78 & ~n79;
  assign n81 = x00 & ~n80;
  assign n82 = x05 & x09;
  assign n83 = ~x01 & ~n30;
  assign n84 = n82 & ~n83;
  assign n85 = ~n81 & ~n84;
  assign n86 = n74 & ~n85;
  assign n87 = ~n73 & ~n86;
  assign n88 = ~x00 & x05;
  assign n89 = ~x07 & x11;
  assign n90 = x03 & n89;
  assign n91 = ~x08 & x11;
  assign n92 = ~x02 & x07;
  assign n93 = n91 & ~n92;
  assign n94 = ~n90 & ~n93;
  assign n95 = ~n88 & ~n94;
  assign n96 = ~x05 & x11;
  assign n97 = ~x00 & ~n96;
  assign n98 = x06 & ~x09;
  assign n99 = ~n28 & ~n98;
  assign n100 = n80 & ~n99;
  assign n101 = ~n97 & ~n100;
  assign n102 = ~n95 & ~n101;
  assign n103 = x01 & ~n102;
  assign n104 = x05 & ~x09;
  assign n105 = n24 & ~n104;
  assign n106 = x01 & ~n98;
  assign n107 = x10 & n106;
  assign n108 = ~n59 & n78;
  assign n109 = ~n107 & ~n108;
  assign n110 = x05 & x12;
  assign n111 = ~n109 & n110;
  assign n112 = ~x06 & x11;
  assign n113 = x02 & x09;
  assign n114 = ~x05 & x10;
  assign n115 = n113 & n114;
  assign n116 = ~x03 & x08;
  assign n117 = ~n92 & ~n116;
  assign n118 = ~n115 & ~n117;
  assign n119 = ~n78 & n118;
  assign n120 = n112 & ~n119;
  assign n121 = ~n88 & n120;
  assign n122 = ~n111 & ~n121;
  assign n123 = ~n105 & n122;
  assign n124 = ~n103 & n123;
  assign z2 = ~n87 | ~n124;
  assign n126 = ~x03 & n52;
  assign n127 = x03 & ~x04;
  assign n128 = ~x04 & ~n51;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n126 & ~n129;
  assign n131 = x07 & x12;
  assign n132 = ~x02 & ~x11;
  assign n133 = ~n92 & ~n132;
  assign n134 = ~n131 & ~n133;
  assign n135 = n130 & ~n134;
  assign n136 = n25 & ~n134;
  assign n137 = ~n135 & ~n136;
  assign n138 = ~n31 & n137;
  assign n139 = ~x05 & n138;
  assign n140 = ~n74 & ~n112;
  assign n141 = ~n139 & ~n140;
  assign n142 = ~x01 & ~n141;
  assign n143 = ~n82 & n142;
  assign n144 = x04 & ~x08;
  assign n145 = ~x03 & ~n128;
  assign n146 = ~n126 & ~n145;
  assign n147 = ~x07 & ~n146;
  assign n148 = ~n144 & ~n147;
  assign n149 = ~x00 & ~n148;
  assign n150 = ~x01 & n149;
  assign n151 = x00 & x05;
  assign n152 = ~x06 & n137;
  assign n153 = ~n151 & n152;
  assign n154 = ~n150 & ~n153;
  assign n155 = ~n31 & ~n154;
  assign n156 = x07 & ~x12;
  assign n157 = ~x02 & n156;
  assign n158 = ~x04 & ~n126;
  assign n159 = ~n157 & n158;
  assign n160 = ~x09 & ~n159;
  assign n161 = ~x12 & ~n79;
  assign n162 = n66 & ~n161;
  assign n163 = ~x11 & ~n162;
  assign n164 = ~x09 & n163;
  assign n165 = ~n160 & ~n164;
  assign n166 = ~x05 & ~x06;
  assign n167 = ~x11 & ~x12;
  assign n168 = ~n31 & n167;
  assign n169 = ~n79 & n168;
  assign n170 = n166 & n169;
  assign n171 = n165 & ~n170;
  assign n172 = ~n155 & n171;
  assign n173 = ~n143 & n172;
  assign n174 = ~x10 & ~n173;
  assign n175 = n41 & ~n130;
  assign n176 = ~n134 & ~n175;
  assign n177 = ~n38 & ~n176;
  assign n178 = x05 & ~x12;
  assign n179 = ~x11 & n178;
  assign n180 = ~x03 & x07;
  assign n181 = x02 & ~n180;
  assign n182 = n179 & ~n181;
  assign n183 = ~n177 & ~n182;
  assign n184 = n98 & ~n183;
  assign n185 = n97 & ~n110;
  assign n186 = x00 & ~n104;
  assign n187 = ~x02 & ~n146;
  assign n188 = ~n134 & ~n140;
  assign n189 = ~n187 & n188;
  assign n190 = ~n186 & ~n189;
  assign n191 = x07 & ~n39;
  assign n192 = ~n130 & n191;
  assign n193 = x04 & x08;
  assign n194 = ~x02 & n193;
  assign n195 = ~n179 & ~n194;
  assign n196 = ~n192 & n195;
  assign n197 = ~n38 & ~n196;
  assign n198 = ~x09 & n197;
  assign n199 = ~n190 & ~n198;
  assign n200 = ~x01 & ~n199;
  assign n201 = ~n185 & ~n200;
  assign n202 = ~n184 & n201;
  assign z3 = n174 | ~n202;
  assign n204 = x00 & ~x10;
  assign n205 = ~x09 & ~n135;
  assign n206 = n138 & n166;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~n143 & n207;
  assign n209 = n204 & ~n208;
  assign n210 = x04 & ~x10;
  assign n211 = x12 & n210;
  assign n212 = ~x09 & x11;
  assign n213 = n211 & n212;
  assign n214 = x12 & n88;
  assign n215 = ~x07 & ~x11;
  assign n216 = ~n145 & ~n215;
  assign n217 = ~x02 & ~n216;
  assign n218 = ~n29 & n217;
  assign n219 = ~n60 & ~n218;
  assign n220 = n214 & ~n219;
  assign n221 = ~n213 & ~n220;
  assign n222 = ~x02 & ~x08;
  assign n223 = n210 & n222;
  assign n224 = ~x07 & ~x10;
  assign n225 = ~n25 & n224;
  assign n226 = n129 & n225;
  assign n227 = ~n223 & ~n226;
  assign n228 = x01 & x06;
  assign n229 = n214 & ~n228;
  assign n230 = ~n227 & n229;
  assign n231 = x06 & ~x12;
  assign n232 = ~n157 & ~n231;
  assign n233 = ~n228 & ~n232;
  assign n234 = ~n25 & ~n31;
  assign n235 = ~n228 & n234;
  assign n236 = ~x04 & ~x08;
  assign n237 = ~x04 & x12;
  assign n238 = ~n236 & ~n237;
  assign n239 = n235 & n238;
  assign n240 = ~n233 & ~n239;
  assign n241 = ~n160 & n240;
  assign n242 = n23 & ~n241;
  assign n243 = x11 & n242;
  assign n244 = ~n230 & ~n243;
  assign n245 = n221 & n244;
  assign n246 = x00 & ~x09;
  assign n247 = x05 & n246;
  assign n248 = ~x01 & ~n74;
  assign n249 = ~n112 & n248;
  assign n250 = ~x11 & n231;
  assign n251 = ~n181 & n250;
  assign n252 = ~n37 & ~n176;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n249 & n253;
  assign n255 = n247 & ~n254;
  assign n256 = ~x09 & n110;
  assign n257 = ~n128 & n191;
  assign n258 = ~n194 & ~n257;
  assign n259 = ~n217 & n258;
  assign n260 = ~n37 & ~n259;
  assign n261 = n132 & n224;
  assign n262 = ~x10 & n129;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n60 & n263;
  assign n265 = ~n260 & n264;
  assign n266 = n256 & ~n265;
  assign n267 = ~n255 & ~n266;
  assign n268 = ~x00 & x11;
  assign n269 = x06 & x07;
  assign n270 = n235 & ~n269;
  assign n271 = ~x01 & n222;
  assign n272 = ~n270 & ~n271;
  assign n273 = n211 & ~n272;
  assign n274 = x07 & ~x09;
  assign n275 = ~n39 & n274;
  assign n276 = ~n158 & n275;
  assign n277 = ~x01 & n231;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~x05 & ~n278;
  assign n280 = x04 & x12;
  assign n281 = n275 & n280;
  assign n282 = ~n279 & ~n281;
  assign n283 = ~n37 & ~n282;
  assign n284 = ~x09 & n193;
  assign n285 = ~n37 & n284;
  assign n286 = ~x03 & x04;
  assign n287 = ~n126 & ~n286;
  assign n288 = ~n156 & n287;
  assign n289 = ~n106 & ~n288;
  assign n290 = ~n285 & ~n289;
  assign n291 = ~n178 & ~n290;
  assign n292 = ~x02 & n291;
  assign n293 = ~n283 & ~n292;
  assign n294 = ~n273 & n293;
  assign n295 = n268 & ~n294;
  assign n296 = n267 & ~n295;
  assign n297 = n245 & n296;
  assign n298 = ~n209 & n297;
  assign n299 = ~x13 & ~n298;
  assign n300 = x09 & x10;
  assign n301 = ~n140 & n300;
  assign n302 = ~n23 & ~n104;
  assign n303 = ~x04 & n302;
  assign n304 = ~n48 & ~n114;
  assign n305 = ~x05 & x08;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & ~n306;
  assign n308 = x03 & ~n307;
  assign n309 = x05 & ~x07;
  assign n310 = ~n76 & ~n82;
  assign n311 = ~n309 & ~n310;
  assign n312 = ~n308 & ~n311;
  assign n313 = ~n249 & ~n312;
  assign n314 = x08 & x12;
  assign n315 = ~x04 & n314;
  assign n316 = ~n59 & n315;
  assign n317 = ~x01 & x06;
  assign n318 = n236 & ~n317;
  assign n319 = x11 & n318;
  assign n320 = ~n316 & ~n319;
  assign n321 = n302 & ~n320;
  assign n322 = ~n313 & ~n321;
  assign n323 = ~n301 & n322;
  assign n324 = x02 & ~n323;
  assign n325 = ~x07 & ~x08;
  assign n326 = x01 & n303;
  assign n327 = n325 & n326;
  assign n328 = ~n300 & ~n306;
  assign n329 = x12 & ~n328;
  assign n330 = ~x06 & n300;
  assign n331 = ~n307 & ~n317;
  assign n332 = ~n330 & ~n331;
  assign n333 = ~x07 & ~n332;
  assign n334 = ~n329 & ~n333;
  assign n335 = x03 & ~n334;
  assign n336 = ~n327 & ~n335;
  assign n337 = x11 & ~n336;
  assign n338 = x09 & ~n28;
  assign n339 = ~n166 & ~n338;
  assign n340 = x01 & ~n23;
  assign n341 = ~n339 & n340;
  assign n342 = x13 & n302;
  assign n343 = n26 & n75;
  assign n344 = n74 & n343;
  assign n345 = ~n342 & ~n344;
  assign n346 = x08 & n326;
  assign n347 = ~n308 & ~n346;
  assign n348 = ~n59 & n131;
  assign n349 = ~n347 & n348;
  assign n350 = n345 & ~n349;
  assign n351 = x06 & x08;
  assign n352 = x07 & n351;
  assign n353 = x11 & ~n156;
  assign n354 = ~n52 & n353;
  assign n355 = ~n352 & ~n354;
  assign n356 = ~n231 & n303;
  assign n357 = ~n355 & n356;
  assign n358 = n350 & ~n357;
  assign n359 = ~n341 & n358;
  assign n360 = ~n337 & n359;
  assign n361 = ~n324 & n360;
  assign n362 = x00 & ~n361;
  assign n363 = ~n299 & ~n362;
  assign n364 = ~n246 & n318;
  assign n365 = ~n330 & ~n364;
  assign n366 = x11 & ~n365;
  assign n367 = ~x01 & ~n112;
  assign n368 = ~n193 & ~n210;
  assign n369 = x03 & n368;
  assign n370 = ~x00 & n369;
  assign n371 = x03 & x09;
  assign n372 = ~n144 & n371;
  assign n373 = ~n370 & ~n372;
  assign n374 = ~x00 & n76;
  assign n375 = ~n75 & ~n374;
  assign n376 = n373 & n375;
  assign n377 = ~n367 & ~n376;
  assign n378 = ~n366 & ~n377;
  assign n379 = x02 & ~n378;
  assign n380 = ~n317 & ~n373;
  assign n381 = ~x03 & ~n364;
  assign n382 = ~n365 & ~n381;
  assign n383 = ~n380 & ~n382;
  assign n384 = n89 & ~n383;
  assign n385 = ~x13 & ~n29;
  assign n386 = x09 & ~n385;
  assign n387 = x10 & n37;
  assign n388 = ~x13 & ~n387;
  assign n389 = ~x00 & ~n388;
  assign n390 = ~n386 & ~n389;
  assign n391 = ~n384 & n390;
  assign n392 = ~n379 & n391;
  assign n393 = n178 & ~n392;
  assign n394 = ~n110 & ~n204;
  assign n395 = x13 & n394;
  assign n396 = ~n247 & n395;
  assign n397 = x04 & ~n48;
  assign n398 = x03 & ~n397;
  assign n399 = ~n75 & ~n398;
  assign n400 = x02 & ~n399;
  assign n401 = ~n338 & ~n400;
  assign n402 = ~n246 & ~n401;
  assign n403 = n394 & n402;
  assign n404 = x10 & ~x12;
  assign n405 = ~n114 & ~n404;
  assign n406 = x07 & x08;
  assign n407 = n181 & ~n406;
  assign n408 = x06 & ~n407;
  assign n409 = ~n151 & ~n408;
  assign n410 = ~n405 & n409;
  assign n411 = ~n403 & ~n410;
  assign n412 = x01 & ~n411;
  assign n413 = ~x00 & ~n397;
  assign n414 = ~n64 & n413;
  assign n415 = n315 & n414;
  assign n416 = ~x08 & n26;
  assign n417 = x03 & n414;
  assign n418 = ~n416 & ~n417;
  assign n419 = n131 & ~n418;
  assign n420 = x10 & n162;
  assign n421 = ~x04 & n420;
  assign n422 = ~n419 & ~n421;
  assign n423 = ~n415 & n422;
  assign n424 = x01 & ~n423;
  assign n425 = ~x07 & n30;
  assign n426 = ~n343 & ~n425;
  assign n427 = n113 & ~n224;
  assign n428 = ~x04 & x08;
  assign n429 = ~n47 & ~n428;
  assign n430 = n66 & ~n429;
  assign n431 = ~n427 & ~n430;
  assign n432 = ~n204 & ~n431;
  assign n433 = n426 & ~n432;
  assign n434 = ~n417 & n433;
  assign n435 = n74 & ~n434;
  assign n436 = ~n424 & ~n435;
  assign n437 = ~x05 & ~n436;
  assign n438 = ~n412 & ~n437;
  assign n439 = ~n396 & n438;
  assign n440 = ~x11 & ~n439;
  assign n441 = ~n393 & ~n440;
  assign z4 = ~n363 | ~n441;
  assign n443 = ~x06 & x07;
  assign n444 = n26 & ~n284;
  assign n445 = x01 & ~x10;
  assign n446 = n428 & ~n445;
  assign n447 = ~x01 & n398;
  assign n448 = ~n446 & ~n447;
  assign n449 = ~n444 & n448;
  assign n450 = n443 & ~n449;
  assign n451 = x12 & n450;
  assign n452 = ~n26 & ~n314;
  assign n453 = ~x04 & ~x06;
  assign n454 = ~n445 & n453;
  assign n455 = ~n452 & n454;
  assign n456 = ~n76 & ~n416;
  assign n457 = ~n228 & ~n456;
  assign n458 = ~x01 & ~n399;
  assign n459 = ~n300 & ~n458;
  assign n460 = ~n457 & n459;
  assign n461 = ~n74 & ~n460;
  assign n462 = ~n455 & ~n461;
  assign n463 = x02 & ~n462;
  assign n464 = ~n74 & ~n98;
  assign n465 = x10 & n464;
  assign n466 = ~n248 & ~n465;
  assign n467 = x13 & ~n466;
  assign n468 = ~n463 & ~n467;
  assign n469 = ~n451 & n468;
  assign n470 = ~x11 & ~n469;
  assign n471 = x01 & ~x09;
  assign n472 = ~x01 & n425;
  assign n473 = ~x04 & n93;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~x13 & n474;
  assign n476 = ~n471 & ~n475;
  assign n477 = x09 & ~n144;
  assign n478 = ~x01 & n368;
  assign n479 = n89 & n300;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n477 & n480;
  assign n482 = ~n79 & ~n90;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n427 & ~n483;
  assign n485 = ~n476 & n484;
  assign n486 = n231 & ~n485;
  assign n487 = ~n470 & ~n486;
  assign n488 = ~x12 & n31;
  assign n489 = n270 & ~n488;
  assign n490 = x09 & ~n489;
  assign n491 = n210 & ~n231;
  assign n492 = ~n490 & n491;
  assign n493 = ~n284 & n288;
  assign n494 = ~x02 & ~n493;
  assign n495 = ~n276 & ~n494;
  assign n496 = n59 & ~n495;
  assign n497 = n211 & n271;
  assign n498 = ~x12 & n28;
  assign n499 = x02 & n75;
  assign n500 = n498 & ~n499;
  assign n501 = ~n117 & n500;
  assign n502 = ~n497 & ~n501;
  assign n503 = ~x02 & ~n371;
  assign n504 = ~n39 & n503;
  assign n505 = ~n275 & ~n504;
  assign n506 = n280 & ~n505;
  assign n507 = ~x01 & n506;
  assign n508 = n502 & ~n507;
  assign n509 = ~n496 & n508;
  assign n510 = ~n492 & n509;
  assign n511 = x11 & ~n510;
  assign n512 = ~n138 & ~n169;
  assign n513 = n28 & ~n512;
  assign n514 = x01 & n513;
  assign n515 = ~n217 & n227;
  assign n516 = ~x01 & ~n515;
  assign n517 = n41 & ~n128;
  assign n518 = ~x07 & n132;
  assign n519 = ~n262 & ~n518;
  assign n520 = ~n517 & n519;
  assign n521 = ~x09 & ~n520;
  assign n522 = ~n516 & ~n521;
  assign n523 = n74 & ~n522;
  assign n524 = ~x06 & x10;
  assign n525 = ~n76 & ~n368;
  assign n526 = ~n134 & ~n525;
  assign n527 = ~n524 & ~n526;
  assign n528 = ~x10 & ~n53;
  assign n529 = ~n269 & ~n528;
  assign n530 = ~n146 & ~n529;
  assign n531 = ~n527 & ~n530;
  assign n532 = ~x02 & x06;
  assign n533 = ~n39 & n532;
  assign n534 = ~n130 & n533;
  assign n535 = n531 & ~n534;
  assign n536 = n471 & ~n535;
  assign n537 = ~n523 & ~n536;
  assign n538 = ~n514 & n537;
  assign n539 = ~n511 & n538;
  assign n540 = ~x13 & ~n539;
  assign n541 = x10 & ~n215;
  assign n542 = ~n156 & n541;
  assign n543 = ~n351 & ~n542;
  assign n544 = n371 & ~n543;
  assign n545 = ~n41 & n524;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n134 & ~n546;
  assign n548 = x02 & n91;
  assign n549 = ~n90 & ~n548;
  assign n550 = ~n162 & n549;
  assign n551 = ~n354 & n550;
  assign n552 = ~x04 & ~n551;
  assign n553 = ~n427 & ~n552;
  assign n554 = ~x13 & n553;
  assign n555 = n99 & ~n554;
  assign n556 = ~n547 & ~n555;
  assign n557 = x01 & ~n556;
  assign n558 = ~n540 & ~n557;
  assign z5 = ~n487 | ~n558;
  assign n560 = n371 & n406;
  assign n561 = n132 & n371;
  assign n562 = ~x03 & ~x13;
  assign n563 = n89 & n562;
  assign n564 = ~n561 & ~n563;
  assign n565 = x08 & ~n30;
  assign n566 = ~n564 & n565;
  assign n567 = ~n91 & n562;
  assign n568 = ~n46 & ~n567;
  assign n569 = ~n444 & ~n568;
  assign n570 = x02 & ~x09;
  assign n571 = x10 & ~x11;
  assign n572 = ~n132 & ~n571;
  assign n573 = ~x07 & n572;
  assign n574 = ~n570 & ~n573;
  assign n575 = ~n569 & n574;
  assign n576 = ~n566 & ~n575;
  assign n577 = ~n560 & n576;
  assign n578 = ~x12 & ~n577;
  assign n579 = ~x13 & ~n130;
  assign n580 = n78 & ~n579;
  assign n581 = ~x13 & ~n315;
  assign n582 = ~n572 & ~n581;
  assign n583 = ~x07 & n582;
  assign n584 = ~x02 & n398;
  assign n585 = ~n444 & ~n584;
  assign n586 = n215 & ~n585;
  assign n587 = ~n583 & ~n586;
  assign n588 = ~n580 & n587;
  assign n589 = ~n578 & n588;
  assign n590 = ~n325 & ~n406;
  assign n591 = ~n300 & n590;
  assign n592 = ~n77 & ~n591;
  assign n593 = x03 & n592;
  assign n594 = n225 & n579;
  assign n595 = ~n593 & ~n594;
  assign n596 = x02 & ~n595;
  assign n597 = x09 & n25;
  assign n598 = x10 & ~n504;
  assign n599 = n46 & n89;
  assign n600 = ~n598 & n599;
  assign n601 = x12 & ~x13;
  assign n602 = ~n113 & n601;
  assign n603 = ~n128 & n602;
  assign n604 = ~n369 & n603;
  assign n605 = ~n215 & n604;
  assign n606 = ~n425 & n605;
  assign n607 = ~n600 & ~n606;
  assign n608 = ~n597 & ~n607;
  assign n609 = ~x07 & ~n528;
  assign n610 = ~n146 & ~n609;
  assign n611 = ~n525 & ~n610;
  assign n612 = ~x13 & n570;
  assign n613 = ~n611 & n612;
  assign n614 = ~n608 & ~n613;
  assign n615 = ~n596 & n614;
  assign z6 = ~n589 | ~n615;
  assign n617 = n31 & n249;
  assign n618 = ~n228 & ~n248;
  assign n619 = n37 & n157;
  assign n620 = ~n518 & ~n619;
  assign n621 = n618 & ~n620;
  assign n622 = ~n617 & ~n621;
  assign n623 = n597 & ~n622;
  assign n624 = ~x03 & ~x11;
  assign n625 = ~n31 & ~n64;
  assign n626 = ~x08 & ~n156;
  assign n627 = n618 & n626;
  assign n628 = n625 & n627;
  assign n629 = n37 & n40;
  assign n630 = ~x12 & n629;
  assign n631 = ~n628 & ~n630;
  assign n632 = n624 & ~n631;
  assign n633 = ~n623 & ~n632;
  assign n634 = x00 & ~n633;
  assign n635 = x11 & n156;
  assign n636 = n597 & n635;
  assign n637 = x02 & ~x06;
  assign n638 = ~n228 & ~n532;
  assign n639 = ~n637 & n638;
  assign n640 = n636 & n639;
  assign n641 = ~n634 & ~n640;
  assign n642 = x07 & ~n570;
  assign n643 = n112 & ~n642;
  assign n644 = ~x06 & ~x07;
  assign n645 = n69 & n644;
  assign n646 = ~n92 & n212;
  assign n647 = ~n645 & ~n646;
  assign n648 = x01 & ~n647;
  assign n649 = ~n643 & ~n648;
  assign n650 = n126 & ~n649;
  assign n651 = ~x04 & ~n650;
  assign n652 = n641 & n651;
  assign n653 = ~n48 & ~n116;
  assign n654 = n643 & n653;
  assign n655 = n39 & n645;
  assign n656 = ~n116 & n646;
  assign n657 = ~n655 & ~n656;
  assign n658 = x01 & ~n657;
  assign n659 = x00 & n66;
  assign n660 = ~x11 & ~n659;
  assign n661 = x01 & n79;
  assign n662 = n235 & ~n661;
  assign n663 = ~n660 & n662;
  assign n664 = n61 & n663;
  assign n665 = ~n658 & ~n664;
  assign n666 = ~n654 & n665;
  assign n667 = x04 & n666;
  assign n668 = ~x05 & ~n667;
  assign n669 = ~n652 & n668;
  assign n670 = n236 & n624;
  assign n671 = x04 & ~n59;
  assign n672 = ~n65 & n671;
  assign n673 = ~n670 & ~n672;
  assign n674 = ~x06 & ~n193;
  assign n675 = ~n59 & ~n64;
  assign n676 = ~n674 & n675;
  assign n677 = ~n673 & n676;
  assign n678 = x01 & x07;
  assign n679 = n129 & n678;
  assign n680 = ~n286 & n679;
  assign n681 = ~n677 & ~n680;
  assign n682 = x12 & ~n681;
  assign n683 = ~n91 & n286;
  assign n684 = n133 & ~n367;
  assign n685 = ~n130 & n684;
  assign n686 = ~n683 & n685;
  assign n687 = ~n682 & ~n686;
  assign n688 = n246 & ~n687;
  assign n689 = x01 & n670;
  assign n690 = ~n39 & ~n116;
  assign n691 = ~n351 & ~n690;
  assign n692 = n671 & n691;
  assign n693 = ~n689 & ~n692;
  assign n694 = n229 & n625;
  assign n695 = ~n693 & n694;
  assign n696 = ~n688 & ~n695;
  assign n697 = ~x00 & x12;
  assign n698 = x04 & x11;
  assign n699 = ~n272 & n698;
  assign n700 = ~n128 & ~n144;
  assign n701 = x02 & ~x03;
  assign n702 = n317 & n701;
  assign n703 = n700 & n702;
  assign n704 = x09 & ~x11;
  assign n705 = x08 & n704;
  assign n706 = n37 & n127;
  assign n707 = ~x02 & n706;
  assign n708 = n705 & n707;
  assign n709 = ~n703 & ~n708;
  assign n710 = n309 & ~n709;
  assign n711 = ~n699 & ~n710;
  assign n712 = n697 & ~n711;
  assign n713 = ~x03 & n132;
  assign n714 = ~x01 & n713;
  assign n715 = n61 & ~n714;
  assign n716 = ~n64 & n104;
  assign n717 = ~n212 & ~n716;
  assign n718 = ~x08 & n624;
  assign n719 = x04 & n718;
  assign n720 = ~n717 & ~n719;
  assign n721 = n129 & n720;
  assign n722 = n715 & n721;
  assign n723 = ~n712 & ~n722;
  assign n724 = n696 & n723;
  assign n725 = ~n669 & n724;
  assign n726 = ~x10 & ~n725;
  assign n727 = ~x06 & ~n40;
  assign n728 = ~n92 & n284;
  assign n729 = ~x04 & x09;
  assign n730 = ~n236 & ~n729;
  assign n731 = n157 & ~n730;
  assign n732 = ~n728 & ~n731;
  assign n733 = ~n27 & ~n732;
  assign n734 = ~n193 & ~n642;
  assign n735 = ~n287 & n734;
  assign n736 = ~n733 & ~n735;
  assign n737 = n727 & ~n736;
  assign n738 = n79 & n231;
  assign n739 = n592 & n738;
  assign n740 = ~x04 & n739;
  assign n741 = ~n737 & ~n740;
  assign n742 = ~x05 & ~n741;
  assign n743 = ~n506 & ~n742;
  assign n744 = n268 & ~n743;
  assign n745 = ~n193 & ~n286;
  assign n746 = n117 & n745;
  assign n747 = ~n237 & ~n746;
  assign n748 = ~n40 & n747;
  assign n749 = n112 & ~n748;
  assign n750 = x08 & n286;
  assign n751 = n47 & n127;
  assign n752 = n625 & ~n751;
  assign n753 = ~n40 & ~n112;
  assign n754 = n247 & ~n753;
  assign n755 = ~n752 & n754;
  assign n756 = ~n74 & n755;
  assign n757 = ~n750 & n756;
  assign n758 = ~n749 & n757;
  assign n759 = n180 & n700;
  assign n760 = n127 & n215;
  assign n761 = ~n49 & n760;
  assign n762 = ~n759 & ~n761;
  assign n763 = n532 & ~n762;
  assign n764 = ~x04 & ~x11;
  assign n765 = n593 & n637;
  assign n766 = n764 & n765;
  assign n767 = ~n763 & ~n766;
  assign n768 = n214 & ~n767;
  assign n769 = n41 & n698;
  assign n770 = n47 & n637;
  assign n771 = n760 & n770;
  assign n772 = ~n769 & ~n771;
  assign n773 = n256 & ~n772;
  assign n774 = ~n768 & ~n773;
  assign n775 = ~n758 & n774;
  assign n776 = ~n744 & n775;
  assign n777 = ~x01 & ~n776;
  assign n778 = ~x11 & ~n406;
  assign n779 = ~n745 & ~n778;
  assign n780 = ~n407 & n779;
  assign n781 = n26 & n64;
  assign n782 = ~n180 & ~n781;
  assign n783 = n51 & ~n782;
  assign n784 = ~x04 & n783;
  assign n785 = ~n780 & ~n784;
  assign n786 = n110 & ~n785;
  assign n787 = n697 & n769;
  assign n788 = ~n89 & n416;
  assign n789 = ~n92 & ~n215;
  assign n790 = ~n39 & n789;
  assign n791 = ~n788 & ~n790;
  assign n792 = x12 & ~n117;
  assign n793 = ~n38 & ~n792;
  assign n794 = ~n791 & n793;
  assign n795 = x02 & ~n406;
  assign n796 = ~x04 & n690;
  assign n797 = ~n795 & ~n796;
  assign n798 = x04 & ~n690;
  assign n799 = x01 & ~n97;
  assign n800 = ~n798 & n799;
  assign n801 = n797 & n800;
  assign n802 = n794 & n801;
  assign n803 = x00 & n764;
  assign n804 = n178 & n803;
  assign n805 = ~n698 & ~n803;
  assign n806 = ~n38 & ~n88;
  assign n807 = ~x08 & n806;
  assign n808 = ~n805 & n807;
  assign n809 = ~n804 & ~n808;
  assign n810 = n678 & n701;
  assign n811 = ~n809 & n810;
  assign n812 = ~n802 & ~n811;
  assign n813 = ~n787 & n812;
  assign n814 = ~n786 & n813;
  assign n815 = n98 & ~n814;
  assign n816 = ~x13 & ~n815;
  assign n817 = ~n777 & n816;
  assign n818 = ~n726 & n817;
  assign n819 = ~x10 & ~n42;
  assign n820 = ~n247 & n464;
  assign n821 = ~x09 & ~n234;
  assign n822 = ~x06 & ~n571;
  assign n823 = ~n214 & ~n822;
  assign n824 = ~n821 & n823;
  assign n825 = ~n792 & n824;
  assign n826 = x11 & ~n67;
  assign n827 = n825 & ~n826;
  assign n828 = n820 & n827;
  assign n829 = ~n819 & n828;
  assign n830 = x09 & n51;
  assign n831 = ~x05 & n443;
  assign n832 = n830 & n831;
  assign n833 = n76 & n351;
  assign n834 = n178 & n833;
  assign n835 = ~n832 & ~n834;
  assign n836 = n701 & ~n835;
  assign n837 = ~x11 & n597;
  assign n838 = ~n718 & ~n837;
  assign n839 = ~x05 & n644;
  assign n840 = ~n838 & n839;
  assign n841 = ~n50 & n167;
  assign n842 = ~n116 & ~n416;
  assign n843 = n178 & n269;
  assign n844 = ~n842 & n843;
  assign n845 = ~n841 & ~n844;
  assign n846 = ~n840 & n845;
  assign n847 = ~x02 & ~n846;
  assign n848 = n705 & n831;
  assign n849 = x06 & ~x07;
  assign n850 = n178 & n849;
  assign n851 = n47 & n850;
  assign n852 = ~n848 & ~n851;
  assign n853 = n79 & ~n852;
  assign n854 = x03 & n590;
  assign n855 = n167 & ~n854;
  assign n856 = ~n77 & n855;
  assign n857 = ~n853 & ~n856;
  assign n858 = ~n847 & n857;
  assign n859 = ~n836 & n858;
  assign n860 = ~x00 & ~n859;
  assign n861 = n404 & ~n690;
  assign n862 = x06 & n38;
  assign n863 = n625 & n862;
  assign n864 = n861 & n863;
  assign n865 = n690 & n704;
  assign n866 = ~n92 & n151;
  assign n867 = n727 & n866;
  assign n868 = n865 & n867;
  assign n869 = ~n864 & ~n868;
  assign n870 = ~n860 & n869;
  assign n871 = n41 & n82;
  assign n872 = n114 & n234;
  assign n873 = ~n871 & ~n872;
  assign n874 = n167 & ~n873;
  assign n875 = ~x01 & ~n874;
  assign n876 = n870 & n875;
  assign n877 = n806 & n830;
  assign n878 = n269 & n877;
  assign n879 = n644 & ~n806;
  assign n880 = n404 & n879;
  assign n881 = x08 & n880;
  assign n882 = ~n878 & ~n881;
  assign n883 = n701 & ~n882;
  assign n884 = x02 & n52;
  assign n885 = ~n65 & n156;
  assign n886 = ~n884 & ~n885;
  assign n887 = ~n63 & ~n886;
  assign n888 = x02 & n51;
  assign n889 = ~n116 & n215;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~n88 & ~n890;
  assign n892 = ~n887 & ~n891;
  assign n893 = n300 & ~n892;
  assign n894 = ~n883 & ~n893;
  assign n895 = ~x10 & ~n352;
  assign n896 = n24 & ~n895;
  assign n897 = x09 & n896;
  assign n898 = n63 & n269;
  assign n899 = n705 & n898;
  assign n900 = ~x08 & n879;
  assign n901 = x09 & ~n96;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n405 & ~n902;
  assign n904 = ~n899 & ~n903;
  assign n905 = ~n897 & n904;
  assign n906 = n79 & ~n905;
  assign n907 = n443 & ~n806;
  assign n908 = n861 & n907;
  assign n909 = n806 & n849;
  assign n910 = n865 & n909;
  assign n911 = ~n908 & ~n910;
  assign n912 = ~x02 & ~n911;
  assign n913 = x01 & ~n912;
  assign n914 = ~n906 & n913;
  assign n915 = n894 & n914;
  assign n916 = ~n876 & ~n915;
  assign n917 = x13 & ~n916;
  assign n918 = ~n829 & n917;
  assign n919 = ~n818 & ~n918;
  assign n920 = ~n98 & ~n730;
  assign n921 = n661 & n920;
  assign n922 = ~n105 & ~n185;
  assign n923 = ~n274 & ~n895;
  assign n924 = ~n922 & n923;
  assign n925 = n921 & n924;
  assign z7 = n919 | n925;
endmodule


