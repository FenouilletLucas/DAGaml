// Benchmark "mult_8" written by ABC on Sat Apr 23 20:18:05 2016

module mult_8 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n34, n35, n36, n37, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
    n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n492, n493, n494, n495, n496, n497, n498, n499,
    n501;
  assign po00 = pi00 & pi08;
  assign n34 = pi01 & pi08;
  assign n35 = pi00 & pi09;
  assign n36 = n34 & n35;
  assign n37 = ~n34 & ~n35;
  assign po01 = ~n36 & ~n37;
  assign n39 = pi02 & pi08;
  assign n40 = pi01 & pi09;
  assign n41 = pi00 & pi10;
  assign n42 = n40 & n41;
  assign n43 = ~n40 & ~n41;
  assign n44 = ~n42 & ~n43;
  assign n45 = ~n39 & ~n44;
  assign n46 = n39 & n44;
  assign n47 = ~n45 & ~n46;
  assign n48 = ~n36 & n47;
  assign n49 = n36 & ~n47;
  assign po02 = n48 | n49;
  assign n51 = pi03 & pi08;
  assign n52 = pi02 & pi09;
  assign n53 = n51 & n52;
  assign n54 = ~n51 & ~n52;
  assign n55 = ~n53 & ~n54;
  assign n56 = pi00 & pi11;
  assign n57 = pi01 & pi10;
  assign n58 = ~n35 & n57;
  assign n59 = n56 & ~n58;
  assign n60 = ~n56 & n58;
  assign n61 = ~n59 & ~n60;
  assign n62 = n55 & ~n61;
  assign n63 = ~n55 & n61;
  assign n64 = ~n62 & ~n63;
  assign n65 = n36 & ~n45;
  assign n66 = ~n46 & ~n65;
  assign n67 = n64 & n66;
  assign n68 = ~n64 & ~n66;
  assign po03 = n67 | n68;
  assign n70 = n56 & n57;
  assign n71 = ~n42 & ~n70;
  assign n72 = pi03 & pi09;
  assign n73 = pi04 & pi08;
  assign n74 = n72 & n73;
  assign n75 = ~n72 & ~n73;
  assign n76 = ~n74 & ~n75;
  assign n77 = pi00 & pi12;
  assign n78 = pi01 & pi11;
  assign n79 = pi02 & pi10;
  assign n80 = n78 & n79;
  assign n81 = ~n78 & ~n79;
  assign n82 = ~n80 & ~n81;
  assign n83 = n77 & ~n82;
  assign n84 = ~n77 & n82;
  assign n85 = ~n83 & ~n84;
  assign n86 = n76 & ~n85;
  assign n87 = ~n76 & n85;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n53 & n88;
  assign n90 = n53 & ~n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = n71 & n91;
  assign n93 = ~n71 & ~n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = ~n62 & n66;
  assign n96 = ~n63 & ~n95;
  assign n97 = n94 & n96;
  assign n98 = ~n94 & ~n96;
  assign po04 = ~n97 & ~n98;
  assign n100 = n53 & ~n87;
  assign n101 = ~n86 & ~n100;
  assign n102 = pi00 & pi13;
  assign n103 = pi02 & pi11;
  assign n104 = pi03 & pi10;
  assign n105 = n103 & n104;
  assign n106 = ~n103 & ~n104;
  assign n107 = ~n105 & ~n106;
  assign n108 = n102 & ~n107;
  assign n109 = ~n102 & n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = pi01 & pi12;
  assign n112 = pi04 & pi09;
  assign n113 = pi05 & pi08;
  assign n114 = n112 & n113;
  assign n115 = ~n112 & ~n113;
  assign n116 = ~n114 & ~n115;
  assign n117 = n74 & n116;
  assign n118 = ~n74 & ~n116;
  assign n119 = ~n117 & ~n118;
  assign n120 = ~n111 & n119;
  assign n121 = n111 & ~n119;
  assign n122 = ~n120 & ~n121;
  assign n123 = ~n110 & ~n122;
  assign n124 = n110 & n122;
  assign n125 = ~n123 & ~n124;
  assign n126 = n77 & ~n81;
  assign n127 = ~n80 & ~n126;
  assign n128 = ~n125 & ~n127;
  assign n129 = n125 & n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = n101 & n130;
  assign n132 = ~n101 & ~n130;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n92 & n96;
  assign n135 = ~n93 & ~n134;
  assign n136 = ~n133 & n135;
  assign n137 = n133 & ~n135;
  assign po05 = ~n136 & ~n137;
  assign n139 = pi05 & pi09;
  assign n140 = pi06 & pi08;
  assign n141 = n139 & n140;
  assign n142 = ~n139 & ~n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = pi00 & pi14;
  assign n145 = pi01 & pi13;
  assign n146 = pi04 & pi10;
  assign n147 = n145 & n146;
  assign n148 = ~n145 & ~n146;
  assign n149 = ~n147 & ~n148;
  assign n150 = ~n144 & ~n149;
  assign n151 = n144 & n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = n143 & n152;
  assign n154 = ~n143 & ~n152;
  assign n155 = ~n153 & ~n154;
  assign n156 = n102 & ~n106;
  assign n157 = ~n105 & ~n156;
  assign n158 = ~n155 & ~n157;
  assign n159 = n155 & n157;
  assign n160 = ~n158 & ~n159;
  assign n161 = n111 & ~n118;
  assign n162 = ~n117 & ~n161;
  assign n163 = n160 & n162;
  assign n164 = ~n160 & ~n162;
  assign n165 = ~n163 & ~n164;
  assign n166 = pi02 & pi12;
  assign n167 = pi03 & pi11;
  assign n168 = n114 & n167;
  assign n169 = ~n114 & ~n167;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n166 & n170;
  assign n172 = n166 & ~n170;
  assign n173 = ~n171 & ~n172;
  assign n174 = n165 & ~n173;
  assign n175 = ~n165 & n173;
  assign n176 = ~n174 & ~n175;
  assign n177 = ~n124 & ~n127;
  assign n178 = ~n123 & ~n177;
  assign n179 = n176 & ~n178;
  assign n180 = ~n176 & n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = ~n132 & n135;
  assign n183 = ~n131 & ~n182;
  assign n184 = ~n181 & n183;
  assign n185 = n181 & ~n183;
  assign po06 = n184 | n185;
  assign n187 = pi00 & pi15;
  assign n188 = pi01 & pi14;
  assign n189 = pi05 & pi10;
  assign n190 = n188 & n189;
  assign n191 = ~n188 & ~n189;
  assign n192 = ~n190 & ~n191;
  assign n193 = ~n187 & ~n192;
  assign n194 = n187 & n192;
  assign n195 = ~n193 & ~n194;
  assign n196 = n166 & ~n169;
  assign n197 = ~n168 & ~n196;
  assign n198 = ~n195 & n197;
  assign n199 = n195 & ~n197;
  assign n200 = ~n198 & ~n199;
  assign n201 = pi03 & pi12;
  assign n202 = pi02 & pi13;
  assign n203 = pi04 & pi11;
  assign n204 = n202 & n203;
  assign n205 = ~n202 & ~n203;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n201 & ~n206;
  assign n208 = n201 & n206;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~n200 & ~n209;
  assign n211 = n200 & n209;
  assign n212 = ~n210 & ~n211;
  assign n213 = ~n154 & ~n157;
  assign n214 = ~n153 & ~n213;
  assign n215 = n212 & ~n214;
  assign n216 = ~n212 & n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = pi06 & pi09;
  assign n219 = pi07 & pi08;
  assign n220 = n218 & n219;
  assign n221 = ~n218 & ~n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = n144 & ~n148;
  assign n224 = ~n147 & ~n223;
  assign n225 = n141 & ~n224;
  assign n226 = ~n141 & n224;
  assign n227 = ~n225 & ~n226;
  assign n228 = ~n222 & n227;
  assign n229 = n222 & ~n227;
  assign n230 = ~n228 & ~n229;
  assign n231 = ~n217 & ~n230;
  assign n232 = n217 & n230;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n163 & ~n173;
  assign n235 = ~n164 & ~n234;
  assign n236 = ~n233 & ~n235;
  assign n237 = n233 & n235;
  assign n238 = ~n236 & ~n237;
  assign n239 = ~n180 & n183;
  assign n240 = ~n179 & ~n239;
  assign n241 = ~n238 & ~n240;
  assign n242 = n238 & n240;
  assign po07 = n241 | n242;
  assign n244 = ~n216 & ~n230;
  assign n245 = ~n215 & ~n244;
  assign n246 = n201 & ~n205;
  assign n247 = ~n204 & ~n246;
  assign n248 = n222 & ~n226;
  assign n249 = ~n225 & ~n248;
  assign n250 = n247 & n249;
  assign n251 = ~n247 & ~n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = pi02 & pi14;
  assign n254 = pi03 & pi13;
  assign n255 = n220 & n254;
  assign n256 = ~n220 & ~n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = n253 & ~n257;
  assign n259 = ~n253 & n257;
  assign n260 = ~n258 & ~n259;
  assign n261 = n252 & ~n260;
  assign n262 = ~n252 & n260;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n199 & ~n209;
  assign n265 = ~n198 & ~n264;
  assign n266 = n263 & n265;
  assign n267 = ~n263 & ~n265;
  assign n268 = ~n266 & ~n267;
  assign n269 = pi07 & pi09;
  assign n270 = pi06 & pi10;
  assign n271 = n269 & n270;
  assign n272 = ~n269 & ~n270;
  assign n273 = ~n271 & ~n272;
  assign n274 = n187 & ~n191;
  assign n275 = ~n190 & ~n274;
  assign n276 = pi04 & pi12;
  assign n277 = pi01 & pi15;
  assign n278 = pi05 & pi11;
  assign n279 = n277 & n278;
  assign n280 = ~n277 & ~n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~n276 & ~n281;
  assign n283 = n276 & n281;
  assign n284 = ~n282 & ~n283;
  assign n285 = ~n275 & n284;
  assign n286 = n275 & ~n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~n273 & n287;
  assign n289 = n273 & ~n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n268 & ~n290;
  assign n292 = n268 & n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = n245 & n293;
  assign n295 = ~n245 & ~n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = ~n237 & ~n240;
  assign n298 = ~n236 & ~n297;
  assign n299 = ~n296 & n298;
  assign n300 = n296 & ~n298;
  assign po08 = ~n299 & ~n300;
  assign n302 = ~n266 & n290;
  assign n303 = ~n267 & ~n302;
  assign n304 = pi03 & pi14;
  assign n305 = pi04 & pi13;
  assign n306 = pi05 & pi12;
  assign n307 = n305 & n306;
  assign n308 = ~n305 & ~n306;
  assign n309 = ~n307 & ~n308;
  assign n310 = ~n304 & ~n309;
  assign n311 = n304 & n309;
  assign n312 = ~n310 & ~n311;
  assign n313 = n276 & ~n280;
  assign n314 = ~n279 & ~n313;
  assign n315 = n312 & ~n314;
  assign n316 = ~n312 & n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~n271 & n317;
  assign n319 = n271 & ~n317;
  assign n320 = ~n318 & ~n319;
  assign n321 = n253 & ~n256;
  assign n322 = ~n255 & ~n321;
  assign n323 = ~n320 & ~n322;
  assign n324 = n320 & n322;
  assign n325 = ~n323 & ~n324;
  assign n326 = pi02 & pi15;
  assign n327 = pi07 & pi10;
  assign n328 = pi06 & pi11;
  assign n329 = n327 & n328;
  assign n330 = ~n327 & ~n328;
  assign n331 = ~n329 & ~n330;
  assign n332 = n326 & ~n331;
  assign n333 = ~n326 & n331;
  assign n334 = ~n332 & ~n333;
  assign n335 = n325 & n334;
  assign n336 = ~n325 & ~n334;
  assign n337 = ~n335 & ~n336;
  assign n338 = ~n250 & ~n260;
  assign n339 = ~n251 & ~n338;
  assign n340 = n337 & n339;
  assign n341 = ~n337 & ~n339;
  assign n342 = ~n340 & ~n341;
  assign n343 = n273 & ~n286;
  assign n344 = ~n285 & ~n343;
  assign n345 = ~n342 & n344;
  assign n346 = n342 & ~n344;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~n303 & ~n347;
  assign n349 = n303 & n347;
  assign n350 = ~n348 & ~n349;
  assign n351 = ~n294 & ~n298;
  assign n352 = ~n295 & ~n351;
  assign n353 = ~n350 & n352;
  assign n354 = n350 & ~n352;
  assign po09 = ~n353 & ~n354;
  assign n356 = ~n340 & ~n344;
  assign n357 = ~n341 & ~n356;
  assign n358 = ~n324 & ~n334;
  assign n359 = ~n323 & ~n358;
  assign n360 = pi03 & pi15;
  assign n361 = pi07 & pi11;
  assign n362 = pi06 & pi12;
  assign n363 = n361 & n362;
  assign n364 = ~n361 & ~n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = n360 & ~n365;
  assign n367 = ~n360 & n365;
  assign n368 = ~n366 & ~n367;
  assign n369 = pi04 & pi14;
  assign n370 = pi05 & pi13;
  assign n371 = n326 & ~n330;
  assign n372 = ~n329 & ~n371;
  assign n373 = n370 & ~n372;
  assign n374 = ~n370 & n372;
  assign n375 = ~n373 & ~n374;
  assign n376 = n369 & ~n375;
  assign n377 = ~n369 & n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = n368 & n378;
  assign n380 = ~n368 & ~n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = ~n304 & ~n307;
  assign n383 = ~n308 & ~n382;
  assign n384 = ~n381 & ~n383;
  assign n385 = n381 & n383;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n359 & n386;
  assign n388 = n359 & ~n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = n271 & ~n316;
  assign n391 = ~n315 & ~n390;
  assign n392 = n389 & n391;
  assign n393 = ~n389 & ~n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n357 & ~n394;
  assign n396 = n357 & n394;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n348 & ~n352;
  assign n399 = ~n349 & ~n398;
  assign n400 = ~n397 & ~n399;
  assign n401 = n397 & n399;
  assign po10 = n400 | n401;
  assign n403 = ~n379 & n383;
  assign n404 = ~n380 & ~n403;
  assign n405 = pi05 & pi14;
  assign n406 = pi04 & pi15;
  assign n407 = pi07 & pi12;
  assign n408 = pi06 & pi13;
  assign n409 = n407 & n408;
  assign n410 = ~n407 & ~n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = n406 & ~n411;
  assign n413 = ~n406 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = n360 & ~n364;
  assign n416 = ~n363 & ~n415;
  assign n417 = ~n414 & ~n416;
  assign n418 = n414 & n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = n405 & ~n419;
  assign n421 = ~n405 & n419;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~n404 & ~n422;
  assign n424 = n404 & n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = n369 & ~n374;
  assign n427 = ~n373 & ~n426;
  assign n428 = ~n425 & ~n427;
  assign n429 = n425 & n427;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~n387 & n391;
  assign n432 = ~n388 & ~n431;
  assign n433 = n430 & ~n432;
  assign n434 = ~n430 & n432;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~n395 & n399;
  assign n437 = ~n396 & ~n436;
  assign n438 = ~n435 & n437;
  assign n439 = n435 & ~n437;
  assign po11 = n438 | n439;
  assign n441 = ~n423 & n427;
  assign n442 = ~n424 & ~n441;
  assign n443 = n406 & ~n410;
  assign n444 = ~n409 & ~n443;
  assign n445 = pi05 & pi15;
  assign n446 = pi07 & pi13;
  assign n447 = pi06 & pi14;
  assign n448 = ~n446 & ~n447;
  assign n449 = n446 & n447;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~n445 & ~n450;
  assign n452 = n445 & n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = n405 & ~n418;
  assign n455 = ~n417 & ~n454;
  assign n456 = ~n453 & n455;
  assign n457 = n453 & ~n455;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~n444 & ~n458;
  assign n460 = n444 & n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n442 & n461;
  assign n463 = n442 & ~n461;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~n434 & ~n437;
  assign n466 = ~n433 & ~n465;
  assign n467 = ~n464 & ~n466;
  assign n468 = n464 & n466;
  assign po12 = ~n467 & ~n468;
  assign n470 = ~n444 & ~n456;
  assign n471 = ~n457 & ~n470;
  assign n472 = pi06 & pi15;
  assign n473 = pi07 & pi14;
  assign n474 = n445 & ~n448;
  assign n475 = ~n408 & ~n474;
  assign n476 = n473 & ~n475;
  assign n477 = ~n473 & ~n474;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n472 & n478;
  assign n480 = n472 & ~n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = n471 & n481;
  assign n483 = ~n462 & n466;
  assign n484 = ~n463 & ~n483;
  assign n485 = n482 & n484;
  assign n486 = ~n471 & ~n481;
  assign n487 = n484 & ~n486;
  assign n488 = ~n482 & ~n487;
  assign n489 = ~n485 & ~n488;
  assign n490 = ~n484 & n486;
  assign po13 = n489 | n490;
  assign n492 = pi07 & pi15;
  assign n493 = n472 & ~n477;
  assign n494 = ~n476 & ~n493;
  assign n495 = ~n492 & n494;
  assign n496 = n492 & ~n494;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n488 & ~n497;
  assign n499 = n488 & n497;
  assign po14 = ~n498 & ~n499;
  assign n501 = ~n488 & ~n496;
  assign po15 = ~n495 & ~n501;
endmodule


