// Benchmark "alu4_cl" written by ABC on Tue May 16 16:07:44 2017

module alu4_cl ( 
    a, b, c, d, e, f, g, h, i, j,
    k, l, m, n, o, p  );
  input  a, b, c, d, e, f, g, h, i, j;
  output k, l, m, n, o, p;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n227, n228, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n529, n530;
  assign n17 = ~e & ~f;
  assign n18 = a & c;
  assign n19 = e & f;
  assign n20 = g & ~h;
  assign n21 = ~a & c;
  assign n22 = f & j;
  assign n23 = ~g & ~j;
  assign n24 = ~h & n23;
  assign n25 = ~f & n23;
  assign n26 = ~n24 & ~n25;
  assign n27 = a & ~c;
  assign n28 = e & ~f;
  assign n29 = ~g & ~h;
  assign n30 = ~j & n29;
  assign n31 = g & j;
  assign n32 = ~n30 & ~n31;
  assign n33 = ~a & ~c;
  assign n34 = ~f & g;
  assign n35 = e & ~j;
  assign n36 = n34 & n35;
  assign n37 = h & n36;
  assign n38 = ~e & n22;
  assign n39 = ~n20 & n38;
  assign n40 = n19 & n20;
  assign n41 = ~n39 & ~n40;
  assign n42 = ~n37 & n41;
  assign n43 = j & n18;
  assign n44 = ~g & n43;
  assign n45 = h & n44;
  assign n46 = n17 & n45;
  assign n47 = n19 & n45;
  assign n48 = ~e & n18;
  assign n49 = n20 & n48;
  assign n50 = ~f & n49;
  assign n51 = ~e & n20;
  assign n52 = n22 & n51;
  assign n53 = n21 & n52;
  assign n54 = ~e & ~n26;
  assign n55 = ~a & n54;
  assign n56 = n27 & n38;
  assign n57 = ~n32 & ~n33;
  assign n58 = n28 & n57;
  assign n59 = ~c & ~n42;
  assign n60 = ~n58 & ~n59;
  assign n61 = ~n56 & n60;
  assign n62 = ~n55 & n61;
  assign n63 = ~n53 & n62;
  assign n64 = ~n50 & n63;
  assign n65 = ~n47 & n64;
  assign n66 = ~n46 & n65;
  assign n67 = a & ~n66;
  assign n68 = e & ~g;
  assign n69 = ~e & g;
  assign n70 = ~e & h;
  assign n71 = a & ~e;
  assign n72 = ~g & ~n66;
  assign n73 = g & n66;
  assign n74 = ~n72 & ~n73;
  assign n75 = a & g;
  assign n76 = ~g & n19;
  assign n77 = n22 & n70;
  assign n78 = j & n20;
  assign n79 = n66 & n78;
  assign n80 = n17 & n79;
  assign n81 = n28 & n78;
  assign n82 = n18 & n81;
  assign n83 = n67 & n78;
  assign n84 = n19 & n83;
  assign n85 = a & n77;
  assign n86 = ~n66 & n77;
  assign n87 = ~n85 & ~n86;
  assign n88 = ~n84 & n87;
  assign n89 = ~n82 & n88;
  assign n90 = ~n80 & n89;
  assign n91 = ~g & n77;
  assign n92 = n18 & n91;
  assign n93 = n78 & n90;
  assign n94 = n28 & n93;
  assign n95 = ~n92 & ~n94;
  assign n96 = ~e & f;
  assign n97 = g & n19;
  assign n98 = ~h & j;
  assign n99 = ~n66 & n98;
  assign n100 = n34 & n99;
  assign n101 = e & n100;
  assign n102 = n95 & n101;
  assign n103 = ~g & j;
  assign n104 = h & n103;
  assign n105 = n96 & n104;
  assign n106 = ~n90 & n105;
  assign n107 = n95 & n106;
  assign n108 = n66 & n98;
  assign n109 = n34 & n108;
  assign n110 = e & n109;
  assign n111 = ~n95 & n110;
  assign n112 = n90 & n105;
  assign n113 = ~n95 & n112;
  assign n114 = ~a & n98;
  assign n115 = n34 & n114;
  assign n116 = ~n90 & n115;
  assign n117 = ~e & n116;
  assign n118 = h & j;
  assign n119 = ~n66 & n118;
  assign n120 = ~a & n119;
  assign n121 = n17 & n120;
  assign n122 = ~f & j;
  assign n123 = ~g & n122;
  assign n124 = e & n123;
  assign n125 = n21 & n124;
  assign n126 = n27 & n124;
  assign n127 = ~h & n122;
  assign n128 = n90 & n127;
  assign n129 = n71 & n128;
  assign n130 = n66 & n123;
  assign n131 = n71 & n130;
  assign n132 = h & n31;
  assign n133 = ~n66 & n132;
  assign n134 = ~a & n133;
  assign n135 = ~h & n103;
  assign n136 = ~n19 & n135;
  assign n137 = a & n136;
  assign n138 = n75 & n118;
  assign n139 = ~n19 & n138;
  assign n140 = n66 & n139;
  assign n141 = n19 & n104;
  assign n142 = n66 & n141;
  assign n143 = n97 & n98;
  assign n144 = n90 & n143;
  assign n145 = n96 & n98;
  assign n146 = ~n74 & n145;
  assign n147 = ~a & n118;
  assign n148 = n97 & n147;
  assign n149 = ~n146 & ~n148;
  assign n150 = ~n144 & n149;
  assign n151 = ~n142 & n150;
  assign n152 = ~n140 & n151;
  assign n153 = ~n137 & n152;
  assign n154 = ~n134 & n153;
  assign n155 = ~n131 & n154;
  assign n156 = ~n129 & n155;
  assign n157 = ~n126 & n156;
  assign n158 = ~n125 & n157;
  assign n159 = ~n121 & n158;
  assign n160 = ~n117 & n159;
  assign n161 = ~n113 & n160;
  assign n162 = ~n111 & n161;
  assign n163 = ~n107 & n162;
  assign n164 = ~n102 & n163;
  assign n165 = ~h & ~j;
  assign n166 = e & n165;
  assign n167 = ~f & n166;
  assign n168 = n66 & n167;
  assign n169 = ~g & n168;
  assign n170 = ~c & n165;
  assign n171 = e & n170;
  assign n172 = ~f & n171;
  assign n173 = g & n172;
  assign n174 = f & n35;
  assign n175 = g & n174;
  assign n176 = n67 & n175;
  assign n177 = ~e & ~j;
  assign n178 = f & n177;
  assign n179 = n33 & n178;
  assign n180 = n20 & n179;
  assign n181 = h & ~j;
  assign n182 = ~f & n181;
  assign n183 = n68 & n182;
  assign n184 = n21 & n183;
  assign n185 = ~n66 & n182;
  assign n186 = g & n185;
  assign n187 = f & ~j;
  assign n188 = n69 & n187;
  assign n189 = n18 & n188;
  assign n190 = f & n181;
  assign n191 = n18 & n190;
  assign n192 = c & ~j;
  assign n193 = f & n192;
  assign n194 = n70 & n193;
  assign n195 = n71 & n182;
  assign n196 = n69 & n182;
  assign n197 = n27 & n182;
  assign n198 = ~f & n177;
  assign n199 = ~n74 & n198;
  assign n200 = ~j & n72;
  assign n201 = c & n200;
  assign n202 = ~e & n201;
  assign n203 = n75 & n181;
  assign n204 = j & n76;
  assign n205 = ~h & n204;
  assign n206 = j & n164;
  assign n207 = ~i & n206;
  assign n208 = j & ~n164;
  assign n209 = i & n208;
  assign n210 = ~n207 & ~n209;
  assign n211 = ~n205 & n210;
  assign n212 = ~n203 & n211;
  assign n213 = ~n202 & n212;
  assign n214 = ~n199 & n213;
  assign n215 = ~n197 & n214;
  assign n216 = ~n196 & n215;
  assign n217 = ~n195 & n216;
  assign n218 = ~n194 & n217;
  assign n219 = ~n191 & n218;
  assign n220 = ~n189 & n219;
  assign n221 = ~n186 & n220;
  assign n222 = ~n184 & n221;
  assign n223 = ~n180 & n222;
  assign n224 = ~n176 & n223;
  assign n225 = ~n173 & n224;
  assign k = n169 | ~n225;
  assign n227 = ~b & d;
  assign n228 = b & ~d;
  assign n = b & d;
  assign n230 = ~g & n;
  assign n231 = ~b & ~d;
  assign n232 = ~f & n;
  assign n233 = n20 & n232;
  assign n234 = ~e & j;
  assign n235 = n20 & n234;
  assign n236 = ~n21 & n235;
  assign n237 = f & n236;
  assign n238 = n227 & n237;
  assign n239 = ~n21 & n234;
  assign n240 = f & n239;
  assign n241 = n228 & n240;
  assign n242 = h & n234;
  assign n243 = ~f & n242;
  assign n244 = n75 & n243;
  assign n245 = j & n230;
  assign n246 = ~e & n245;
  assign n247 = h & n246;
  assign n248 = ~f & n247;
  assign n249 = j & n231;
  assign n250 = ~e & n249;
  assign n251 = n21 & n250;
  assign n252 = f & n251;
  assign n253 = n21 & n235;
  assign n254 = n & n253;
  assign n255 = n22 & n230;
  assign n256 = e & n255;
  assign n257 = h & n256;
  assign n258 = ~b & n54;
  assign n259 = ~n32 & ~n231;
  assign n260 = n28 & n259;
  assign n261 = ~e & n233;
  assign n262 = j & n233;
  assign n263 = ~d & ~n42;
  assign n264 = ~n262 & ~n263;
  assign n265 = ~n261 & n264;
  assign n266 = ~n260 & n265;
  assign n267 = ~n258 & n266;
  assign n268 = ~n257 & n267;
  assign n269 = ~n254 & n268;
  assign n270 = ~n252 & n269;
  assign n271 = ~n248 & n270;
  assign n272 = ~n244 & n271;
  assign n273 = ~n241 & n272;
  assign n274 = ~n238 & n273;
  assign n275 = b & ~n274;
  assign n276 = b & ~e;
  assign n277 = ~n90 & ~n95;
  assign n278 = n81 & n;
  assign n279 = n78 & n274;
  assign n280 = n17 & n279;
  assign n281 = n78 & n275;
  assign n282 = n19 & n281;
  assign n283 = b & n77;
  assign n284 = n77 & ~n274;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n282 & n285;
  assign n287 = ~n280 & n286;
  assign n288 = ~n278 & n287;
  assign n289 = n77 & n230;
  assign n290 = n78 & n288;
  assign n291 = n28 & n290;
  assign n292 = ~n289 & ~n291;
  assign n293 = ~n66 & ~n95;
  assign n294 = a & ~n90;
  assign n295 = n288 & n294;
  assign n296 = ~n288 & ~n294;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n34 & ~n69;
  assign n299 = ~n17 & n298;
  assign n300 = n67 & ~n274;
  assign n301 = ~n67 & n274;
  assign n302 = ~n300 & ~n301;
  assign n303 = n66 & n274;
  assign n304 = ~f & n68;
  assign n305 = n18 & n304;
  assign n306 = n90 & n288;
  assign n307 = n19 & n306;
  assign n308 = n105 & ~n288;
  assign n309 = n292 & n308;
  assign n310 = ~n277 & n309;
  assign n311 = n105 & n288;
  assign n312 = ~n292 & n311;
  assign n313 = ~n277 & n312;
  assign n314 = n292 & n311;
  assign n315 = n277 & n314;
  assign n316 = ~n292 & n308;
  assign n317 = n277 & n316;
  assign n318 = ~h & n31;
  assign n319 = ~n274 & n318;
  assign n320 = n28 & n319;
  assign n321 = n292 & n320;
  assign n322 = ~n293 & n321;
  assign n323 = n274 & n318;
  assign n324 = n28 & n323;
  assign n325 = ~n292 & n324;
  assign n326 = ~n293 & n325;
  assign n327 = n292 & n324;
  assign n328 = n293 & n327;
  assign n329 = ~n292 & n320;
  assign n330 = n293 & n329;
  assign n331 = n19 & n132;
  assign n332 = ~b & n331;
  assign n333 = ~a & n332;
  assign n334 = n19 & n318;
  assign n335 = ~n90 & n334;
  assign n336 = ~n288 & n335;
  assign n337 = ~n297 & n318;
  assign n338 = ~b & n337;
  assign n339 = n17 & n338;
  assign n340 = n19 & n118;
  assign n341 = b & n340;
  assign n342 = n75 & n341;
  assign n343 = ~n274 & n340;
  assign n344 = n72 & n343;
  assign n345 = j & n302;
  assign n346 = h & n345;
  assign n347 = ~b & n346;
  assign n348 = ~n299 & n347;
  assign n349 = j & ~n302;
  assign n350 = h & n349;
  assign n351 = b & n350;
  assign n352 = ~n299 & n351;
  assign n353 = n145 & ~n274;
  assign n354 = ~n66 & n353;
  assign n355 = n141 & n303;
  assign n356 = n96 & n318;
  assign n357 = n303 & n356;
  assign n358 = b & n136;
  assign n359 = n96 & n135;
  assign n360 = ~n274 & n359;
  assign n361 = j & n276;
  assign n362 = ~f & n361;
  assign n363 = ~h & n362;
  assign n364 = n297 & n363;
  assign n365 = n276 & n349;
  assign n366 = ~f & n365;
  assign n367 = ~g & n366;
  assign n368 = j & n304;
  assign n369 = ~n18 & n368;
  assign n370 = n228 & n369;
  assign n371 = n227 & n369;
  assign n372 = j & n305;
  assign n373 = h & n372;
  assign n374 = n231 & n373;
  assign n375 = n307 & n318;
  assign n376 = ~h & n368;
  assign n377 = d & n376;
  assign n378 = n & n372;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n375 & n379;
  assign n381 = ~n374 & n380;
  assign n382 = ~n371 & n381;
  assign n383 = ~n370 & n382;
  assign n384 = ~n367 & n383;
  assign n385 = ~n364 & n384;
  assign n386 = ~n360 & n385;
  assign n387 = ~n358 & n386;
  assign n388 = ~n357 & n387;
  assign n389 = ~n355 & n388;
  assign n390 = ~n354 & n389;
  assign n391 = ~n352 & n390;
  assign n392 = ~n348 & n391;
  assign n393 = ~n344 & n392;
  assign n394 = ~n342 & n393;
  assign n395 = ~n339 & n394;
  assign n396 = ~n336 & n395;
  assign n397 = ~n333 & n396;
  assign n398 = ~n330 & n397;
  assign n399 = ~n328 & n398;
  assign n400 = ~n326 & n399;
  assign n401 = ~n322 & n400;
  assign n402 = ~n317 & n401;
  assign n403 = ~n315 & n402;
  assign n404 = ~n313 & n403;
  assign n405 = ~n310 & n404;
  assign n406 = ~e & ~g;
  assign n407 = ~n274 & n406;
  assign n408 = ~f & n165;
  assign n409 = ~g & n408;
  assign n410 = n274 & n409;
  assign n411 = e & n410;
  assign n412 = ~d & n165;
  assign n413 = ~f & n412;
  assign n414 = g & n413;
  assign n415 = e & n414;
  assign n416 = ~e & n187;
  assign n417 = n20 & n416;
  assign n418 = n231 & n417;
  assign n419 = g & n187;
  assign n420 = e & n419;
  assign n421 = n275 & n420;
  assign n422 = n183 & n227;
  assign n423 = g & n182;
  assign n424 = ~n274 & n423;
  assign n425 = n188 & n;
  assign n426 = n190 & n;
  assign n427 = d & ~j;
  assign n428 = f & n427;
  assign n429 = n70 & n428;
  assign n430 = n182 & n276;
  assign n431 = n182 & n228;
  assign n432 = ~f & ~j;
  assign n433 = n69 & n432;
  assign n434 = n274 & n433;
  assign n435 = b & n181;
  assign n436 = g & n435;
  assign n437 = j & n405;
  assign n438 = ~n164 & n437;
  assign n439 = ~i & n438;
  assign n440 = ~j & n407;
  assign n441 = ~f & n440;
  assign n442 = d & n440;
  assign n443 = j & ~n405;
  assign n444 = i & n443;
  assign n445 = n164 & n443;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n205 & n446;
  assign n448 = ~n442 & n447;
  assign n449 = ~n441 & n448;
  assign n450 = ~n439 & n449;
  assign n451 = ~n436 & n450;
  assign n452 = ~n196 & n451;
  assign n453 = ~n434 & n452;
  assign n454 = ~n431 & n453;
  assign n455 = ~n430 & n454;
  assign n456 = ~n429 & n455;
  assign n457 = ~n426 & n456;
  assign n458 = ~n425 & n457;
  assign n459 = ~n424 & n458;
  assign n460 = ~n422 & n459;
  assign n461 = ~n421 & n460;
  assign n462 = ~n418 & n461;
  assign n463 = ~n415 & n462;
  assign l = n411 | ~n463;
  assign m = n | n231;
  assign n466 = n34 & n98;
  assign n467 = e & n466;
  assign n468 = ~n274 & n467;
  assign n469 = n293 & n468;
  assign n470 = ~n292 & n467;
  assign n471 = n293 & n470;
  assign n472 = ~n274 & n470;
  assign n473 = n96 & n118;
  assign n474 = ~g & n473;
  assign n475 = ~n292 & n474;
  assign n476 = n277 & n475;
  assign n477 = n118 & ~n288;
  assign n478 = n96 & n477;
  assign n479 = ~g & n478;
  assign n480 = n277 & n479;
  assign n481 = ~n292 & n479;
  assign n482 = ~n288 & n466;
  assign n483 = ~e & n482;
  assign n484 = b & n483;
  assign n485 = n294 & n482;
  assign n486 = ~e & n485;
  assign n487 = n118 & ~n299;
  assign n488 = n67 & n487;
  assign n489 = ~n274 & n488;
  assign n490 = b & n487;
  assign n491 = n67 & n490;
  assign n492 = n97 & n118;
  assign n493 = ~a & n492;
  assign n494 = ~b & n493;
  assign n495 = n276 & n466;
  assign n496 = n294 & n495;
  assign n497 = j & n303;
  assign n498 = ~h & n497;
  assign n499 = n69 & n498;
  assign n500 = f & n499;
  assign n501 = n275 & n487;
  assign n502 = n118 & n304;
  assign n503 = n & n502;
  assign n504 = n118 & n305;
  assign n505 = ~n231 & n504;
  assign n506 = ~n164 & n443;
  assign n507 = ~i & n506;
  assign n508 = n98 & n307;
  assign n509 = n76 & n497;
  assign n510 = ~n205 & ~n509;
  assign n511 = ~n508 & n510;
  assign n512 = ~n507 & n511;
  assign n513 = ~n505 & n512;
  assign n514 = ~n503 & n513;
  assign n515 = ~n501 & n514;
  assign n516 = ~n500 & n515;
  assign n517 = ~n496 & n516;
  assign n518 = ~n494 & n517;
  assign n519 = ~n491 & n518;
  assign n520 = ~n489 & n519;
  assign n521 = ~n486 & n520;
  assign n522 = ~n484 & n521;
  assign n523 = ~n481 & n522;
  assign n524 = ~n480 & n523;
  assign n525 = ~n476 & n524;
  assign n526 = ~n472 & n525;
  assign n527 = ~n471 & n526;
  assign o = n469 | ~n527;
  assign n529 = n33 & m;
  assign n530 = n18 & m;
  assign p = n529 | n530;
endmodule


