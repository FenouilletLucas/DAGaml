// Benchmark "i7" written by ABC on Tue May 16 16:07:50 2017

module i7 ( 
    \V160(21) , \V160(20) , \V160(23) , \V160(22) , \V128(27) , \V160(25) ,
    \V128(26) , \V160(24) , \V128(29) , \V160(17) , \V128(28) , \V160(16) ,
    \V160(19) , \V160(18) , \V96(0) , \V96(1) , \V64(13) , \V96(2) ,
    \V64(12) , \V96(3) , \V64(15) , \V128(21) , \V96(4) , \V64(14) ,
    \V128(20) , \V96(5) , \V128(23) , \V160(11) , \V96(6) , \V128(22) ,
    \V160(10) , \V96(7) , \V64(11) , \V128(25) , \V160(13) , \V96(8) ,
    \V64(10) , \V128(24) , \V192(3) , \V160(12) , \V96(9) , \V128(17) ,
    \V192(2) , \V160(15) , \V128(16) , \V192(5) , \V160(14) , \V128(19) ,
    \V192(4) , \V128(18) , \V64(17) , \V64(16) , \V192(1) , \V64(19) ,
    \V192(0) , \V64(18) , \V64(23) , \V64(22) , \V64(25) , \V128(11) ,
    \V64(24) , \V128(10) , \V192(7) , \V128(13) , \V192(6) , \V128(12) ,
    \V192(9) , \V64(21) , \V128(15) , \V192(8) , \V64(20) , \V128(14) ,
    \V64(27) , \V64(26) , \V64(29) , \V64(28) , \V194(1) , \V160(31) ,
    \V194(0) , \V160(30) , \V64(31) , \V64(30) , \V128(3) , \V128(2) ,
    \V128(5) , \V195(0) , \V128(4) , \V128(31) , \V128(30) , \V128(1) ,
    \V128(0) , \V128(7) , \V128(6) , \V128(9) , \V128(8) , \V199(3) ,
    \V199(4) , \V199(1) , \V199(0) , \V32(0) , \V32(1) , \V32(2) ,
    \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) , \V32(15) ,
    \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) , \V32(11) ,
    \V32(10) , \V192(27) , \V192(26) , \V192(29) , \V192(28) , \V32(17) ,
    \V32(16) , \V32(19) , \V32(18) , \V32(23) , \V32(22) , \V192(21) ,
    \V32(25) , \V192(20) , \V32(24) , \V192(23) , \V192(22) , \V192(25) ,
    \V32(21) , \V192(24) , \V32(20) , \V192(17) , \V192(16) , \V192(19) ,
    \V192(18) , \V32(27) , \V96(13) , \V32(26) , \V96(12) , \V32(29) ,
    \V96(15) , \V32(28) , \V96(14) , \V192(11) , \V192(10) , \V96(11) ,
    \V192(13) , \V96(10) , \V192(12) , \V192(15) , \V32(31) , \V192(14) ,
    \V32(30) , \V96(17) , \V96(16) , \V96(19) , \V96(18) , \V96(23) ,
    \V96(22) , \V96(25) , \V96(24) , \V96(21) , \V96(20) , \V96(27) ,
    \V96(26) , \V96(29) , \V96(28) , \V192(31) , \V64(0) , \V192(30) ,
    \V96(31) , \V64(1) , \V96(30) , \V64(2) , \V64(3) , \V64(4) , \V64(5) ,
    \V64(6) , \V64(7) , \V64(8) , \V160(3) , \V64(9) , \V160(2) ,
    \V160(5) , \V160(4) , \V160(1) , \V160(0) , \V160(7) , \V160(6) ,
    \V160(9) , \V160(8) , \V160(27) , \V160(26) , \V160(29) , \V160(28) ,
    \V259(27) , \V259(26) , \V259(29) , \V259(28) , \V259(21) , \V259(20) ,
    \V259(23) , \V259(22) , \V259(25) , \V259(24) , \V259(17) , \V259(16) ,
    \V259(19) , \V259(18) , \V259(11) , \V259(10) , \V259(13) , \V259(12) ,
    \V259(15) , \V259(14) , \V259(3) , \V259(2) , \V259(5) , \V259(4) ,
    \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) , \V259(8) ,
    \V259(31) , \V259(30) , \V227(27) , \V227(26) , \V227(21) , \V227(20) ,
    \V227(23) , \V227(22) , \V227(25) , \V227(24) , \V227(17) , \V227(16) ,
    \V227(19) , \V227(18) , \V227(11) , \V227(10) , \V227(13) , \V227(12) ,
    \V227(15) , \V227(14) , \V266(3) , \V266(2) , \V266(5) , \V266(4) ,
    \V266(1) , \V266(0) , \V266(6) , \V227(3) , \V227(2) , \V227(5) ,
    \V227(4) , \V227(1) , \V227(0) , \V227(7) , \V227(6) , \V227(9) ,
    \V227(8)   );
  input  \V160(21) , \V160(20) , \V160(23) , \V160(22) , \V128(27) ,
    \V160(25) , \V128(26) , \V160(24) , \V128(29) , \V160(17) , \V128(28) ,
    \V160(16) , \V160(19) , \V160(18) , \V96(0) , \V96(1) , \V64(13) ,
    \V96(2) , \V64(12) , \V96(3) , \V64(15) , \V128(21) , \V96(4) ,
    \V64(14) , \V128(20) , \V96(5) , \V128(23) , \V160(11) , \V96(6) ,
    \V128(22) , \V160(10) , \V96(7) , \V64(11) , \V128(25) , \V160(13) ,
    \V96(8) , \V64(10) , \V128(24) , \V192(3) , \V160(12) , \V96(9) ,
    \V128(17) , \V192(2) , \V160(15) , \V128(16) , \V192(5) , \V160(14) ,
    \V128(19) , \V192(4) , \V128(18) , \V64(17) , \V64(16) , \V192(1) ,
    \V64(19) , \V192(0) , \V64(18) , \V64(23) , \V64(22) , \V64(25) ,
    \V128(11) , \V64(24) , \V128(10) , \V192(7) , \V128(13) , \V192(6) ,
    \V128(12) , \V192(9) , \V64(21) , \V128(15) , \V192(8) , \V64(20) ,
    \V128(14) , \V64(27) , \V64(26) , \V64(29) , \V64(28) , \V194(1) ,
    \V160(31) , \V194(0) , \V160(30) , \V64(31) , \V64(30) , \V128(3) ,
    \V128(2) , \V128(5) , \V195(0) , \V128(4) , \V128(31) , \V128(30) ,
    \V128(1) , \V128(0) , \V128(7) , \V128(6) , \V128(9) , \V128(8) ,
    \V199(3) , \V199(4) , \V199(1) , \V199(0) , \V32(0) , \V32(1) ,
    \V32(2) , \V32(3) , \V32(13) , \V32(4) , \V32(12) , \V32(5) ,
    \V32(15) , \V32(6) , \V32(14) , \V32(7) , \V32(8) , \V32(9) ,
    \V32(11) , \V32(10) , \V192(27) , \V192(26) , \V192(29) , \V192(28) ,
    \V32(17) , \V32(16) , \V32(19) , \V32(18) , \V32(23) , \V32(22) ,
    \V192(21) , \V32(25) , \V192(20) , \V32(24) , \V192(23) , \V192(22) ,
    \V192(25) , \V32(21) , \V192(24) , \V32(20) , \V192(17) , \V192(16) ,
    \V192(19) , \V192(18) , \V32(27) , \V96(13) , \V32(26) , \V96(12) ,
    \V32(29) , \V96(15) , \V32(28) , \V96(14) , \V192(11) , \V192(10) ,
    \V96(11) , \V192(13) , \V96(10) , \V192(12) , \V192(15) , \V32(31) ,
    \V192(14) , \V32(30) , \V96(17) , \V96(16) , \V96(19) , \V96(18) ,
    \V96(23) , \V96(22) , \V96(25) , \V96(24) , \V96(21) , \V96(20) ,
    \V96(27) , \V96(26) , \V96(29) , \V96(28) , \V192(31) , \V64(0) ,
    \V192(30) , \V96(31) , \V64(1) , \V96(30) , \V64(2) , \V64(3) ,
    \V64(4) , \V64(5) , \V64(6) , \V64(7) , \V64(8) , \V160(3) , \V64(9) ,
    \V160(2) , \V160(5) , \V160(4) , \V160(1) , \V160(0) , \V160(7) ,
    \V160(6) , \V160(9) , \V160(8) , \V160(27) , \V160(26) , \V160(29) ,
    \V160(28) ;
  output \V259(27) , \V259(26) , \V259(29) , \V259(28) , \V259(21) ,
    \V259(20) , \V259(23) , \V259(22) , \V259(25) , \V259(24) , \V259(17) ,
    \V259(16) , \V259(19) , \V259(18) , \V259(11) , \V259(10) , \V259(13) ,
    \V259(12) , \V259(15) , \V259(14) , \V259(3) , \V259(2) , \V259(5) ,
    \V259(4) , \V259(1) , \V259(0) , \V259(7) , \V259(6) , \V259(9) ,
    \V259(8) , \V259(31) , \V259(30) , \V227(27) , \V227(26) , \V227(21) ,
    \V227(20) , \V227(23) , \V227(22) , \V227(25) , \V227(24) , \V227(17) ,
    \V227(16) , \V227(19) , \V227(18) , \V227(11) , \V227(10) , \V227(13) ,
    \V227(12) , \V227(15) , \V227(14) , \V266(3) , \V266(2) , \V266(5) ,
    \V266(4) , \V266(1) , \V266(0) , \V266(6) , \V227(3) , \V227(2) ,
    \V227(5) , \V227(4) , \V227(1) , \V227(0) , \V227(7) , \V227(6) ,
    \V227(9) , \V227(8) ;
  wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n294, n295, n296, n297, n298, n299, n300, n301, n302, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n334, n335, n336, n337, n338, n339, n340, n341, n342, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n374, n375, n376, n377, n378, n379, n380, n381, n382, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n414, n415, n416, n417, n418, n419, n420, n421, n422, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n494, n495, n496, n497, n498, n499, n500, n501, n502, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n534, n535, n536, n537, n538, n539, n540, n541, n542, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n595, n596, n597,
    n598, n599, n600, n601, n602, n604, n605, n606, n607, n608, n609, n610,
    n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, n623, n624,
    n625, n626, n628, n629, n630, n631, n632, n633, n634, n636, n637, n638,
    n639, n640, n641, n642, n644, n645, n646, n647, n648, n649, n650, n652,
    n653, n654, n655, n656, n657, n658, n660, n661, n662, n663, n664, n665,
    n666, n668, n669, n670, n671, n672, n673, n674, n676, n677, n678, n679,
    n680, n681, n682, n684, n685, n686, n687, n688, n689, n690, n692, n693,
    n694, n695, n696, n697, n698, n700, n701, n702, n703, n704, n705, n706,
    n708, n709, n710, n711, n712, n713, n714, n716, n717, n718, n719, n720,
    n721, n722, n724, n725, n726, n727, n728, n729, n730, n732, n733, n734,
    n735, n736, n737, n738, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n754, n755, n756, n757, n758, n759, n760,
    n761, n763, n764, n765, n766, n768, n769, n770, n771, n773, n774, n775,
    n776, n777, n778, n779, n781, n782, n783, n784, n785, n786, n787, n789,
    n790, n792, n793, n794, n795, n796, n797, n798, n800, n801, n802, n803,
    n804, n805, n806, n808, n809, n810, n811, n812, n813, n814, n816, n817,
    n818, n819, n820, n821, n822, n824, n825, n826, n827, n828, n829, n830,
    n832, n833, n834, n835, n836, n837, n838, n840, n841, n842, n843, n844,
    n845, n846, n848, n849, n850, n851, n852, n853, n854, n856, n857, n858,
    n859, n860, n861, n862, n864, n865, n866, n867, n868, n869, n870;
  assign n267 = ~\V199(4)  & \V199(1) ;
  assign n268 = \V199(1)  & ~\V199(0) ;
  assign n269 = \V199(4)  & n268;
  assign n270 = ~\V192(23)  & n269;
  assign n271 = \V160(23)  & \V199(0) ;
  assign n272 = \V199(1)  & n271;
  assign n273 = \V199(4)  & n272;
  assign n274 = ~\V199(1)  & ~\V199(0) ;
  assign n275 = \V199(4)  & n274;
  assign n276 = \V192(23)  & n275;
  assign n277 = ~\V199(1)  & \V199(0) ;
  assign n278 = \V199(4)  & n277;
  assign n279 = \V128(23)  & n278;
  assign n280 = ~n276 & ~n279;
  assign n281 = ~n273 & n280;
  assign n282 = ~n270 & n281;
  assign \V259(27)  = n267 | ~n282;
  assign n284 = ~\V192(22)  & n269;
  assign n285 = \V160(22)  & \V199(0) ;
  assign n286 = \V199(1)  & n285;
  assign n287 = \V199(4)  & n286;
  assign n288 = \V192(22)  & n275;
  assign n289 = \V128(22)  & n278;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n287 & n290;
  assign n292 = ~n284 & n291;
  assign \V259(26)  = n267 | ~n292;
  assign n294 = ~\V192(25)  & n269;
  assign n295 = \V160(25)  & \V199(0) ;
  assign n296 = \V199(1)  & n295;
  assign n297 = \V199(4)  & n296;
  assign n298 = \V192(25)  & n275;
  assign n299 = \V128(25)  & n278;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n297 & n300;
  assign n302 = ~n294 & n301;
  assign \V259(29)  = n267 | ~n302;
  assign n304 = ~\V192(24)  & n269;
  assign n305 = \V160(24)  & \V199(0) ;
  assign n306 = \V199(1)  & n305;
  assign n307 = \V199(4)  & n306;
  assign n308 = \V192(24)  & n275;
  assign n309 = \V128(24)  & n278;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~n307 & n310;
  assign n312 = ~n304 & n311;
  assign \V259(28)  = n267 | ~n312;
  assign n314 = ~\V192(17)  & n269;
  assign n315 = \V160(17)  & \V199(0) ;
  assign n316 = \V199(1)  & n315;
  assign n317 = \V199(4)  & n316;
  assign n318 = \V192(17)  & n275;
  assign n319 = \V128(17)  & n278;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~n317 & n320;
  assign n322 = ~n314 & n321;
  assign \V259(21)  = n267 | ~n322;
  assign n324 = ~\V192(16)  & n269;
  assign n325 = \V160(16)  & \V199(0) ;
  assign n326 = \V199(1)  & n325;
  assign n327 = \V199(4)  & n326;
  assign n328 = \V192(16)  & n275;
  assign n329 = \V128(16)  & n278;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~n327 & n330;
  assign n332 = ~n324 & n331;
  assign \V259(20)  = n267 | ~n332;
  assign n334 = ~\V192(19)  & n269;
  assign n335 = \V160(19)  & \V199(0) ;
  assign n336 = \V199(1)  & n335;
  assign n337 = \V199(4)  & n336;
  assign n338 = \V192(19)  & n275;
  assign n339 = \V128(19)  & n278;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~n337 & n340;
  assign n342 = ~n334 & n341;
  assign \V259(23)  = n267 | ~n342;
  assign n344 = ~\V192(18)  & n269;
  assign n345 = \V160(18)  & \V199(0) ;
  assign n346 = \V199(1)  & n345;
  assign n347 = \V199(4)  & n346;
  assign n348 = \V192(18)  & n275;
  assign n349 = \V128(18)  & n278;
  assign n350 = ~n348 & ~n349;
  assign n351 = ~n347 & n350;
  assign n352 = ~n344 & n351;
  assign \V259(22)  = n267 | ~n352;
  assign n354 = ~\V192(21)  & n269;
  assign n355 = \V160(21)  & \V199(0) ;
  assign n356 = \V199(1)  & n355;
  assign n357 = \V199(4)  & n356;
  assign n358 = \V192(21)  & n275;
  assign n359 = \V128(21)  & n278;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~n354 & n361;
  assign \V259(25)  = n267 | ~n362;
  assign n364 = ~\V192(20)  & n269;
  assign n365 = \V160(20)  & \V199(0) ;
  assign n366 = \V199(1)  & n365;
  assign n367 = \V199(4)  & n366;
  assign n368 = \V192(20)  & n275;
  assign n369 = \V128(20)  & n278;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~n367 & n370;
  assign n372 = ~n364 & n371;
  assign \V259(24)  = n267 | ~n372;
  assign n374 = ~\V192(13)  & n269;
  assign n375 = \V160(13)  & \V199(0) ;
  assign n376 = \V199(1)  & n375;
  assign n377 = \V199(4)  & n376;
  assign n378 = \V192(13)  & n275;
  assign n379 = \V128(13)  & n278;
  assign n380 = ~n378 & ~n379;
  assign n381 = ~n377 & n380;
  assign n382 = ~n374 & n381;
  assign \V259(17)  = n267 | ~n382;
  assign n384 = ~\V192(12)  & n269;
  assign n385 = \V160(12)  & \V199(0) ;
  assign n386 = \V199(1)  & n385;
  assign n387 = \V199(4)  & n386;
  assign n388 = \V192(12)  & n275;
  assign n389 = \V128(12)  & n278;
  assign n390 = ~n388 & ~n389;
  assign n391 = ~n387 & n390;
  assign n392 = ~n384 & n391;
  assign \V259(16)  = n267 | ~n392;
  assign n394 = ~\V192(15)  & n269;
  assign n395 = \V160(15)  & \V199(0) ;
  assign n396 = \V199(1)  & n395;
  assign n397 = \V199(4)  & n396;
  assign n398 = \V192(15)  & n275;
  assign n399 = \V128(15)  & n278;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~n397 & n400;
  assign n402 = ~n394 & n401;
  assign \V259(19)  = n267 | ~n402;
  assign n404 = ~\V192(14)  & n269;
  assign n405 = \V160(14)  & \V199(0) ;
  assign n406 = \V199(1)  & n405;
  assign n407 = \V199(4)  & n406;
  assign n408 = \V192(14)  & n275;
  assign n409 = \V128(14)  & n278;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~n407 & n410;
  assign n412 = ~n404 & n411;
  assign \V259(18)  = n267 | ~n412;
  assign n414 = ~\V192(7)  & n269;
  assign n415 = \V199(0)  & \V160(7) ;
  assign n416 = \V199(1)  & n415;
  assign n417 = \V199(4)  & n416;
  assign n418 = \V192(7)  & n275;
  assign n419 = \V128(7)  & n278;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~n417 & n420;
  assign n422 = ~n414 & n421;
  assign \V259(11)  = n267 | ~n422;
  assign n424 = ~\V192(6)  & n269;
  assign n425 = \V199(0)  & \V160(6) ;
  assign n426 = \V199(1)  & n425;
  assign n427 = \V199(4)  & n426;
  assign n428 = \V192(6)  & n275;
  assign n429 = \V128(6)  & n278;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~n427 & n430;
  assign n432 = ~n424 & n431;
  assign \V259(10)  = n267 | ~n432;
  assign n434 = ~\V192(9)  & n269;
  assign n435 = \V199(0)  & \V160(9) ;
  assign n436 = \V199(1)  & n435;
  assign n437 = \V199(4)  & n436;
  assign n438 = \V192(9)  & n275;
  assign n439 = \V128(9)  & n278;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n437 & n440;
  assign n442 = ~n434 & n441;
  assign \V259(13)  = n267 | ~n442;
  assign n444 = ~\V192(8)  & n269;
  assign n445 = \V199(0)  & \V160(8) ;
  assign n446 = \V199(1)  & n445;
  assign n447 = \V199(4)  & n446;
  assign n448 = \V192(8)  & n275;
  assign n449 = \V128(8)  & n278;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~n447 & n450;
  assign n452 = ~n444 & n451;
  assign \V259(12)  = n267 | ~n452;
  assign n454 = ~\V192(11)  & n269;
  assign n455 = \V160(11)  & \V199(0) ;
  assign n456 = \V199(1)  & n455;
  assign n457 = \V199(4)  & n456;
  assign n458 = \V192(11)  & n275;
  assign n459 = \V128(11)  & n278;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n457 & n460;
  assign n462 = ~n454 & n461;
  assign \V259(15)  = n267 | ~n462;
  assign n464 = ~\V192(10)  & n269;
  assign n465 = \V160(10)  & \V199(0) ;
  assign n466 = \V199(1)  & n465;
  assign n467 = \V199(4)  & n466;
  assign n468 = \V192(10)  & n275;
  assign n469 = \V128(10)  & n278;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~n467 & n470;
  assign n472 = ~n464 & n471;
  assign \V259(14)  = n267 | ~n472;
  assign n474 = ~\V96(31)  & n269;
  assign n475 = \V64(31)  & \V199(0) ;
  assign n476 = \V199(1)  & n475;
  assign n477 = \V199(4)  & n476;
  assign n478 = \V96(31)  & n275;
  assign n479 = \V32(31)  & n278;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n477 & n480;
  assign n482 = ~n474 & n481;
  assign \V259(3)  = n267 | ~n482;
  assign n484 = ~\V96(30)  & n269;
  assign n485 = \V64(30)  & \V199(0) ;
  assign n486 = \V199(1)  & n485;
  assign n487 = \V199(4)  & n486;
  assign n488 = \V96(30)  & n275;
  assign n489 = \V32(30)  & n278;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n487 & n490;
  assign n492 = ~n484 & n491;
  assign \V259(2)  = n267 | ~n492;
  assign n494 = ~\V192(1)  & n269;
  assign n495 = \V199(0)  & \V160(1) ;
  assign n496 = \V199(1)  & n495;
  assign n497 = \V199(4)  & n496;
  assign n498 = \V192(1)  & n275;
  assign n499 = \V128(1)  & n278;
  assign n500 = ~n498 & ~n499;
  assign n501 = ~n497 & n500;
  assign n502 = ~n494 & n501;
  assign \V259(5)  = n267 | ~n502;
  assign n504 = ~\V192(0)  & n269;
  assign n505 = \V199(0)  & \V160(0) ;
  assign n506 = \V199(1)  & n505;
  assign n507 = \V199(4)  & n506;
  assign n508 = \V192(0)  & n275;
  assign n509 = \V128(0)  & n278;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n507 & n510;
  assign n512 = ~n504 & n511;
  assign \V259(4)  = n267 | ~n512;
  assign n514 = ~\V96(29)  & n269;
  assign n515 = \V64(29)  & \V199(0) ;
  assign n516 = \V199(1)  & n515;
  assign n517 = \V199(4)  & n516;
  assign n518 = \V96(29)  & n275;
  assign n519 = \V32(29)  & n278;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n517 & n520;
  assign n522 = ~n514 & n521;
  assign \V259(1)  = n267 | ~n522;
  assign n524 = ~\V96(28)  & n269;
  assign n525 = \V64(28)  & \V199(0) ;
  assign n526 = \V199(1)  & n525;
  assign n527 = \V199(4)  & n526;
  assign n528 = \V96(28)  & n275;
  assign n529 = \V32(28)  & n278;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n527 & n530;
  assign n532 = ~n524 & n531;
  assign \V259(0)  = n267 | ~n532;
  assign n534 = ~\V192(3)  & n269;
  assign n535 = \V199(0)  & \V160(3) ;
  assign n536 = \V199(1)  & n535;
  assign n537 = \V199(4)  & n536;
  assign n538 = \V192(3)  & n275;
  assign n539 = \V128(3)  & n278;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~n537 & n540;
  assign n542 = ~n534 & n541;
  assign \V259(7)  = n267 | ~n542;
  assign n544 = ~\V192(2)  & n269;
  assign n545 = \V199(0)  & \V160(2) ;
  assign n546 = \V199(1)  & n545;
  assign n547 = \V199(4)  & n546;
  assign n548 = \V192(2)  & n275;
  assign n549 = \V128(2)  & n278;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n547 & n550;
  assign n552 = ~n544 & n551;
  assign \V259(6)  = n267 | ~n552;
  assign n554 = ~\V192(5)  & n269;
  assign n555 = \V199(0)  & \V160(5) ;
  assign n556 = \V199(1)  & n555;
  assign n557 = \V199(4)  & n556;
  assign n558 = \V192(5)  & n275;
  assign n559 = \V128(5)  & n278;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n557 & n560;
  assign n562 = ~n554 & n561;
  assign \V259(9)  = n267 | ~n562;
  assign n564 = ~\V192(4)  & n269;
  assign n565 = \V199(0)  & \V160(4) ;
  assign n566 = \V199(1)  & n565;
  assign n567 = \V199(4)  & n566;
  assign n568 = \V192(4)  & n275;
  assign n569 = \V128(4)  & n278;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n567 & n570;
  assign n572 = ~n564 & n571;
  assign \V259(8)  = n267 | ~n572;
  assign n574 = ~\V192(27)  & n269;
  assign n575 = \V199(0)  & \V160(27) ;
  assign n576 = \V199(1)  & n575;
  assign n577 = \V199(4)  & n576;
  assign n578 = \V192(27)  & n275;
  assign n579 = \V128(27)  & n277;
  assign n580 = \V199(4)  & n579;
  assign n581 = ~n578 & ~n580;
  assign n582 = ~n577 & n581;
  assign n583 = ~n574 & n582;
  assign \V259(31)  = n267 | ~n583;
  assign n585 = ~\V192(26)  & n269;
  assign n586 = \V199(0)  & \V160(26) ;
  assign n587 = \V199(1)  & n586;
  assign n588 = \V199(4)  & n587;
  assign n589 = \V192(26)  & n275;
  assign n590 = \V128(26)  & n278;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n588 & n591;
  assign n593 = ~n585 & n592;
  assign \V259(30)  = n267 | ~n593;
  assign n595 = ~\V96(27)  & n268;
  assign n596 = \V64(27)  & \V199(1) ;
  assign n597 = \V199(0)  & n596;
  assign n598 = \V96(27)  & n274;
  assign n599 = ~\V199(1)  & \V32(27) ;
  assign n600 = \V199(0)  & n599;
  assign n601 = ~n598 & ~n600;
  assign n602 = ~n597 & n601;
  assign \V227(27)  = n595 | ~n602;
  assign n604 = ~\V96(26)  & n268;
  assign n605 = \V64(26)  & \V199(1) ;
  assign n606 = \V199(0)  & n605;
  assign n607 = \V96(26)  & n274;
  assign n608 = \V32(26)  & n277;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n606 & n609;
  assign \V227(26)  = n604 | ~n610;
  assign n612 = ~\V96(21)  & n268;
  assign n613 = \V64(21)  & \V199(1) ;
  assign n614 = \V199(0)  & n613;
  assign n615 = \V96(21)  & n274;
  assign n616 = \V32(21)  & n277;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~n614 & n617;
  assign \V227(21)  = n612 | ~n618;
  assign n620 = ~\V96(20)  & n268;
  assign n621 = \V64(20)  & \V199(1) ;
  assign n622 = \V199(0)  & n621;
  assign n623 = \V96(20)  & n274;
  assign n624 = \V32(20)  & n277;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n622 & n625;
  assign \V227(20)  = n620 | ~n626;
  assign n628 = ~\V96(23)  & n268;
  assign n629 = \V64(23)  & \V199(1) ;
  assign n630 = \V199(0)  & n629;
  assign n631 = \V96(23)  & n274;
  assign n632 = \V32(23)  & n277;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~n630 & n633;
  assign \V227(23)  = n628 | ~n634;
  assign n636 = ~\V96(22)  & n268;
  assign n637 = \V64(22)  & \V199(1) ;
  assign n638 = \V199(0)  & n637;
  assign n639 = \V96(22)  & n274;
  assign n640 = \V32(22)  & n277;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n638 & n641;
  assign \V227(22)  = n636 | ~n642;
  assign n644 = ~\V96(25)  & n268;
  assign n645 = \V64(25)  & \V199(1) ;
  assign n646 = \V199(0)  & n645;
  assign n647 = \V96(25)  & n274;
  assign n648 = \V32(25)  & n277;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n646 & n649;
  assign \V227(25)  = n644 | ~n650;
  assign n652 = ~\V96(24)  & n268;
  assign n653 = \V64(24)  & \V199(1) ;
  assign n654 = \V199(0)  & n653;
  assign n655 = \V96(24)  & n274;
  assign n656 = \V32(24)  & n277;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n654 & n657;
  assign \V227(24)  = n652 | ~n658;
  assign n660 = ~\V96(17)  & n268;
  assign n661 = \V64(17)  & \V199(1) ;
  assign n662 = \V199(0)  & n661;
  assign n663 = \V96(17)  & n274;
  assign n664 = \V32(17)  & n277;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~n662 & n665;
  assign \V227(17)  = n660 | ~n666;
  assign n668 = ~\V96(16)  & n268;
  assign n669 = \V64(16)  & \V199(1) ;
  assign n670 = \V199(0)  & n669;
  assign n671 = \V96(16)  & n274;
  assign n672 = \V32(16)  & n277;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n670 & n673;
  assign \V227(16)  = n668 | ~n674;
  assign n676 = ~\V96(19)  & n268;
  assign n677 = \V64(19)  & \V199(1) ;
  assign n678 = \V199(0)  & n677;
  assign n679 = \V96(19)  & n274;
  assign n680 = \V32(19)  & n277;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~n678 & n681;
  assign \V227(19)  = n676 | ~n682;
  assign n684 = ~\V96(18)  & n268;
  assign n685 = \V64(18)  & \V199(1) ;
  assign n686 = \V199(0)  & n685;
  assign n687 = \V96(18)  & n274;
  assign n688 = \V32(18)  & n277;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~n686 & n689;
  assign \V227(18)  = n684 | ~n690;
  assign n692 = ~\V96(11)  & n268;
  assign n693 = \V64(11)  & \V199(1) ;
  assign n694 = \V199(0)  & n693;
  assign n695 = \V96(11)  & n274;
  assign n696 = \V32(11)  & n277;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n694 & n697;
  assign \V227(11)  = n692 | ~n698;
  assign n700 = ~\V96(10)  & n268;
  assign n701 = \V64(10)  & \V199(1) ;
  assign n702 = \V199(0)  & n701;
  assign n703 = \V96(10)  & n274;
  assign n704 = \V32(10)  & n277;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~n702 & n705;
  assign \V227(10)  = n700 | ~n706;
  assign n708 = ~\V96(13)  & n268;
  assign n709 = \V64(13)  & \V199(1) ;
  assign n710 = \V199(0)  & n709;
  assign n711 = \V96(13)  & n274;
  assign n712 = \V32(13)  & n277;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n710 & n713;
  assign \V227(13)  = n708 | ~n714;
  assign n716 = ~\V96(12)  & n268;
  assign n717 = \V64(12)  & \V199(1) ;
  assign n718 = \V199(0)  & n717;
  assign n719 = \V96(12)  & n274;
  assign n720 = \V32(12)  & n277;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n718 & n721;
  assign \V227(12)  = n716 | ~n722;
  assign n724 = ~\V96(15)  & n268;
  assign n725 = \V64(15)  & \V199(1) ;
  assign n726 = \V199(0)  & n725;
  assign n727 = \V96(15)  & n274;
  assign n728 = \V32(15)  & n277;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n726 & n729;
  assign \V227(15)  = n724 | ~n730;
  assign n732 = ~\V96(14)  & n268;
  assign n733 = \V64(14)  & \V199(1) ;
  assign n734 = \V199(0)  & n733;
  assign n735 = \V96(14)  & n274;
  assign n736 = \V32(14)  & n277;
  assign n737 = ~n735 & ~n736;
  assign n738 = ~n734 & n737;
  assign \V227(14)  = n732 | ~n738;
  assign n740 = ~\V199(3)  & \V199(1) ;
  assign n741 = \V199(3)  & n268;
  assign n742 = ~\V192(31)  & n741;
  assign n743 = \V199(3)  & \V199(1) ;
  assign n744 = \V199(0)  & n743;
  assign n745 = \V160(31)  & n744;
  assign n746 = \V199(3)  & n274;
  assign n747 = \V192(31)  & n746;
  assign n748 = \V128(31)  & n277;
  assign n749 = \V199(3)  & n748;
  assign n750 = ~n747 & ~n749;
  assign n751 = ~n745 & n750;
  assign n752 = ~n742 & n751;
  assign \V266(3)  = n740 | ~n752;
  assign n754 = ~\V192(30)  & n741;
  assign n755 = \V160(30)  & n744;
  assign n756 = \V192(30)  & n746;
  assign n757 = \V199(3)  & n277;
  assign n758 = \V128(30)  & n757;
  assign n759 = ~n756 & ~n758;
  assign n760 = ~n755 & n759;
  assign n761 = ~n754 & n760;
  assign \V266(2)  = n740 | ~n761;
  assign n763 = ~\V194(1)  & n741;
  assign n764 = \V194(1)  & n746;
  assign n765 = ~n740 & ~n764;
  assign n766 = ~n744 & n765;
  assign \V266(5)  = n763 | ~n766;
  assign n768 = ~\V194(0)  & n741;
  assign n769 = \V194(0)  & n746;
  assign n770 = ~n740 & ~n769;
  assign n771 = ~n744 & n770;
  assign \V266(4)  = n768 | ~n771;
  assign n773 = ~\V192(29)  & n741;
  assign n774 = \V160(29)  & n744;
  assign n775 = \V192(29)  & n746;
  assign n776 = \V128(29)  & n757;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n774 & n777;
  assign n779 = ~n773 & n778;
  assign \V266(1)  = n740 | ~n779;
  assign n781 = ~\V192(28)  & n741;
  assign n782 = \V160(28)  & n744;
  assign n783 = \V192(28)  & n746;
  assign n784 = \V128(28)  & n757;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n782 & n785;
  assign n787 = ~n781 & n786;
  assign \V266(0)  = n740 | ~n787;
  assign n789 = \V195(0)  & n746;
  assign n790 = \V195(0)  & n741;
  assign \V266(6)  = n789 | n790;
  assign n792 = ~\V96(3)  & n268;
  assign n793 = \V199(1)  & \V64(3) ;
  assign n794 = \V199(0)  & n793;
  assign n795 = \V96(3)  & n274;
  assign n796 = \V32(3)  & n277;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n794 & n797;
  assign \V227(3)  = n792 | ~n798;
  assign n800 = ~\V96(2)  & n268;
  assign n801 = \V199(1)  & \V64(2) ;
  assign n802 = \V199(0)  & n801;
  assign n803 = \V96(2)  & n274;
  assign n804 = \V32(2)  & n277;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n802 & n805;
  assign \V227(2)  = n800 | ~n806;
  assign n808 = ~\V96(5)  & n268;
  assign n809 = \V199(1)  & \V64(5) ;
  assign n810 = \V199(0)  & n809;
  assign n811 = \V96(5)  & n274;
  assign n812 = \V32(5)  & n277;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n810 & n813;
  assign \V227(5)  = n808 | ~n814;
  assign n816 = ~\V96(4)  & n268;
  assign n817 = \V199(1)  & \V64(4) ;
  assign n818 = \V199(0)  & n817;
  assign n819 = \V96(4)  & n274;
  assign n820 = \V32(4)  & n277;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n818 & n821;
  assign \V227(4)  = n816 | ~n822;
  assign n824 = ~\V96(1)  & n268;
  assign n825 = \V199(1)  & \V64(1) ;
  assign n826 = \V199(0)  & n825;
  assign n827 = \V96(1)  & n274;
  assign n828 = \V32(1)  & n277;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n826 & n829;
  assign \V227(1)  = n824 | ~n830;
  assign n832 = ~\V96(0)  & n268;
  assign n833 = \V199(1)  & \V64(0) ;
  assign n834 = \V199(0)  & n833;
  assign n835 = \V96(0)  & n274;
  assign n836 = \V32(0)  & n277;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~n834 & n837;
  assign \V227(0)  = n832 | ~n838;
  assign n840 = ~\V96(7)  & n268;
  assign n841 = \V199(1)  & \V64(7) ;
  assign n842 = \V199(0)  & n841;
  assign n843 = \V96(7)  & n274;
  assign n844 = \V32(7)  & n277;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n842 & n845;
  assign \V227(7)  = n840 | ~n846;
  assign n848 = ~\V96(6)  & n268;
  assign n849 = \V199(1)  & \V64(6) ;
  assign n850 = \V199(0)  & n849;
  assign n851 = \V96(6)  & n274;
  assign n852 = \V32(6)  & n277;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n850 & n853;
  assign \V227(6)  = n848 | ~n854;
  assign n856 = ~\V96(9)  & n268;
  assign n857 = \V199(1)  & \V64(9) ;
  assign n858 = \V199(0)  & n857;
  assign n859 = \V96(9)  & n274;
  assign n860 = \V32(9)  & n277;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n858 & n861;
  assign \V227(9)  = n856 | ~n862;
  assign n864 = ~\V96(8)  & n268;
  assign n865 = \V199(1)  & \V64(8) ;
  assign n866 = \V199(0)  & n865;
  assign n867 = \V96(8)  & n274;
  assign n868 = \V32(8)  & n277;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n866 & n869;
  assign \V227(8)  = n864 | ~n870;
endmodule


