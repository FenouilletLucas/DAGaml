// Benchmark "ttt2" written by ABC on Tue May 16 16:07:53 2017

module ttt2 ( 
    a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0  );
  input  a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y;
  output z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, r0, s0, t0;
  wire n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n60,
    n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
    n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n120, n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n240, n241, n242, n243, n244, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n260, n261, n262, n263,
    n264, n265, n267, n268, n269, n270, n271, n272, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n597, n598, n599,
    n600, n602, n603, n604, n605;
  assign n46 = ~s & ~t;
  assign n47 = ~u & n46;
  assign n48 = v & n47;
  assign n49 = ~e & t;
  assign n50 = v & n49;
  assign n51 = ~e & ~s;
  assign n52 = v & n51;
  assign n53 = u & ~v;
  assign n54 = ~e & u;
  assign n55 = ~n53 & ~n54;
  assign n56 = ~n52 & n55;
  assign n57 = ~n50 & n56;
  assign n58 = ~n48 & n57;
  assign z = ~w & n58;
  assign n60 = q & w;
  assign n61 = q & ~v;
  assign n62 = ~n60 & ~n61;
  assign n63 = ~u & v;
  assign n64 = y & n53;
  assign n65 = ~n63 & ~n64;
  assign n66 = ~t & ~u;
  assign n67 = n65 & n66;
  assign n68 = ~f & n65;
  assign n69 = ~v & n65;
  assign n70 = s & n66;
  assign n71 = ~f & s;
  assign n72 = s & ~v;
  assign n73 = t & n66;
  assign n74 = t & ~v;
  assign n75 = ~f & t;
  assign n76 = ~n74 & ~n75;
  assign n77 = ~n73 & n76;
  assign n78 = ~n72 & n77;
  assign n79 = ~n71 & n78;
  assign n80 = ~n70 & n79;
  assign n81 = ~n69 & n80;
  assign n82 = ~n68 & n81;
  assign n83 = ~n67 & n82;
  assign n84 = ~v & ~y;
  assign n85 = n83 & ~n84;
  assign n86 = n62 & n85;
  assign n87 = ~s & n83;
  assign n88 = n62 & n87;
  assign n89 = t & n83;
  assign n90 = n62 & n89;
  assign n91 = ~u & n83;
  assign n92 = n62 & n91;
  assign n93 = w & ~n84;
  assign n94 = n62 & n93;
  assign n95 = ~s & w;
  assign n96 = n62 & n95;
  assign n97 = t & w;
  assign n98 = n62 & n97;
  assign n99 = ~u & w;
  assign n100 = n62 & n99;
  assign n101 = ~n98 & ~n100;
  assign n102 = ~n96 & n101;
  assign n103 = ~n94 & n102;
  assign n104 = ~n92 & n103;
  assign n105 = ~n90 & n104;
  assign n106 = ~n88 & n105;
  assign a0 = n86 | ~n106;
  assign n108 = ~v & n46;
  assign n109 = y & n108;
  assign n110 = ~u & ~v;
  assign n111 = ~g & v;
  assign n112 = ~n66 & ~n111;
  assign n113 = ~n110 & n112;
  assign n114 = ~n109 & n113;
  assign n115 = ~t & n84;
  assign n116 = s & n115;
  assign n117 = n114 & n116;
  assign n118 = ~w & n114;
  assign b0 = n117 | n118;
  assign n120 = ~v & y;
  assign n121 = q & n46;
  assign n122 = n120 & n121;
  assign n123 = ~v & ~w;
  assign n124 = ~u & n123;
  assign n125 = ~n122 & ~n124;
  assign n126 = u & v;
  assign n127 = t & ~u;
  assign n128 = t & v;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n126 & n129;
  assign n131 = ~q & w;
  assign n132 = n116 & n131;
  assign n133 = n130 & n132;
  assign n134 = n125 & n133;
  assign n135 = ~w & n131;
  assign n136 = n130 & n135;
  assign n137 = n125 & n136;
  assign n138 = ~q & n131;
  assign n139 = n130 & n138;
  assign n140 = n125 & n139;
  assign n141 = u & n116;
  assign n142 = n130 & n141;
  assign n143 = n125 & n142;
  assign n144 = t & n116;
  assign n145 = n130 & n144;
  assign n146 = n125 & n145;
  assign n147 = ~s & n116;
  assign n148 = n130 & n147;
  assign n149 = n125 & n148;
  assign n150 = u & ~w;
  assign n151 = n130 & n150;
  assign n152 = n125 & n151;
  assign n153 = t & ~w;
  assign n154 = n130 & n153;
  assign n155 = n125 & n154;
  assign n156 = ~s & ~w;
  assign n157 = n130 & n156;
  assign n158 = n125 & n157;
  assign n159 = ~q & u;
  assign n160 = n130 & n159;
  assign n161 = n125 & n160;
  assign n162 = ~q & t;
  assign n163 = n130 & n162;
  assign n164 = n125 & n163;
  assign n165 = ~q & ~s;
  assign n166 = n130 & n165;
  assign n167 = n125 & n166;
  assign n168 = h & n132;
  assign n169 = n125 & n168;
  assign n170 = h & n135;
  assign n171 = n125 & n170;
  assign n172 = h & n138;
  assign n173 = n125 & n172;
  assign n174 = h & n141;
  assign n175 = n125 & n174;
  assign n176 = h & n144;
  assign n177 = n125 & n176;
  assign n178 = h & n147;
  assign n179 = n125 & n178;
  assign n180 = h & n150;
  assign n181 = n125 & n180;
  assign n182 = h & n153;
  assign n183 = n125 & n182;
  assign n184 = h & n156;
  assign n185 = n125 & n184;
  assign n186 = h & n159;
  assign n187 = n125 & n186;
  assign n188 = h & n162;
  assign n189 = n125 & n188;
  assign n190 = h & n165;
  assign n191 = n125 & n190;
  assign n192 = w & n116;
  assign n193 = n131 & n192;
  assign n194 = n125 & n193;
  assign n195 = n125 & n131;
  assign n196 = u & w;
  assign n197 = n116 & n196;
  assign n198 = n125 & n197;
  assign n199 = n97 & n116;
  assign n200 = n125 & n199;
  assign n201 = n95 & n116;
  assign n202 = n125 & n201;
  assign n203 = w & n159;
  assign n204 = n125 & n203;
  assign n205 = w & n162;
  assign n206 = n125 & n205;
  assign n207 = w & n165;
  assign n208 = n125 & n207;
  assign n209 = ~n206 & ~n208;
  assign n210 = ~n204 & n209;
  assign n211 = ~n202 & n210;
  assign n212 = ~n200 & n211;
  assign n213 = ~n198 & n212;
  assign n214 = ~n195 & n213;
  assign n215 = ~n194 & n214;
  assign n216 = ~n191 & n215;
  assign n217 = ~n189 & n216;
  assign n218 = ~n187 & n217;
  assign n219 = ~n185 & n218;
  assign n220 = ~n183 & n219;
  assign n221 = ~n181 & n220;
  assign n222 = ~n179 & n221;
  assign n223 = ~n177 & n222;
  assign n224 = ~n175 & n223;
  assign n225 = ~n173 & n224;
  assign n226 = ~n171 & n225;
  assign n227 = ~n169 & n226;
  assign n228 = ~n167 & n227;
  assign n229 = ~n164 & n228;
  assign n230 = ~n161 & n229;
  assign n231 = ~n158 & n230;
  assign n232 = ~n155 & n231;
  assign n233 = ~n152 & n232;
  assign n234 = ~n149 & n233;
  assign n235 = ~n146 & n234;
  assign n236 = ~n143 & n235;
  assign n237 = ~n140 & n236;
  assign n238 = ~n137 & n237;
  assign c0 = n134 | ~n238;
  assign n240 = ~s & ~v;
  assign n241 = ~i & v;
  assign n242 = ~n66 & ~n241;
  assign n243 = ~n240 & n242;
  assign n244 = ~n53 & n243;
  assign d0 = ~w & n244;
  assign n246 = s & t;
  assign n247 = ~v & n246;
  assign n248 = ~j & t;
  assign n249 = v & n248;
  assign n250 = ~j & u;
  assign n251 = ~n249 & ~n250;
  assign n252 = ~n247 & n251;
  assign n253 = ~n48 & n252;
  assign n254 = ~u & ~w;
  assign n255 = n253 & n254;
  assign n256 = v & ~w;
  assign n257 = n253 & n256;
  assign e0 = n255 | n257;
  assign f0 = ~a & ~k;
  assign n260 = ~a & k;
  assign n261 = ~l & n260;
  assign n262 = ~n & n261;
  assign n263 = m & n261;
  assign n264 = l & f0;
  assign n265 = ~n263 & ~n264;
  assign g0 = n262 | ~n265;
  assign n267 = l & n260;
  assign n268 = ~m & n267;
  assign n269 = ~a & ~l;
  assign n270 = m & n269;
  assign n271 = m & f0;
  assign n272 = ~n270 & ~n271;
  assign h0 = n268 | ~n272;
  assign n274 = k & l;
  assign n275 = m & n274;
  assign n276 = n & n275;
  assign n277 = k & ~l;
  assign n278 = ~m & n277;
  assign n279 = ~a & ~n278;
  assign n280 = ~n276 & n279;
  assign n281 = l & m;
  assign n282 = k & n281;
  assign n283 = n280 & n282;
  assign n284 = n & n280;
  assign i0 = n283 | n284;
  assign n286 = ~m & n;
  assign n287 = ~l & n286;
  assign n288 = k & n287;
  assign n289 = n & o;
  assign n290 = ~x & ~n289;
  assign n291 = n288 & n290;
  assign n292 = ~a & n291;
  assign n293 = ~o & ~n289;
  assign n294 = n288 & n293;
  assign n295 = ~a & n294;
  assign n296 = m & ~x;
  assign n297 = n288 & n296;
  assign n298 = ~a & n297;
  assign n299 = l & ~x;
  assign n300 = n288 & n299;
  assign n301 = ~a & n300;
  assign n302 = ~k & ~x;
  assign n303 = n288 & n302;
  assign n304 = ~a & n303;
  assign n305 = m & ~o;
  assign n306 = n288 & n305;
  assign n307 = ~a & n306;
  assign n308 = l & ~o;
  assign n309 = n288 & n308;
  assign n310 = ~a & n309;
  assign n311 = ~k & ~o;
  assign n312 = n288 & n311;
  assign n313 = ~a & n312;
  assign n314 = o & ~x;
  assign n315 = ~n289 & n314;
  assign n316 = ~a & n315;
  assign n317 = ~o & x;
  assign n318 = ~n289 & n317;
  assign n319 = ~a & n318;
  assign n320 = m & o;
  assign n321 = ~x & n320;
  assign n322 = ~a & n321;
  assign n323 = l & o;
  assign n324 = ~x & n323;
  assign n325 = ~a & n324;
  assign n326 = ~k & o;
  assign n327 = ~x & n326;
  assign n328 = ~a & n327;
  assign n329 = x & n305;
  assign n330 = ~a & n329;
  assign n331 = x & n308;
  assign n332 = ~a & n331;
  assign n333 = x & n311;
  assign n334 = ~a & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = ~n330 & n335;
  assign n337 = ~n328 & n336;
  assign n338 = ~n325 & n337;
  assign n339 = ~n322 & n338;
  assign n340 = ~n319 & n339;
  assign n341 = ~n316 & n340;
  assign n342 = ~n313 & n341;
  assign n343 = ~n310 & n342;
  assign n344 = ~n307 & n343;
  assign n345 = ~n304 & n344;
  assign n346 = ~n301 & n345;
  assign n347 = ~n298 & n346;
  assign n348 = ~n295 & n347;
  assign j0 = n292 | ~n348;
  assign n350 = o & ~q;
  assign n351 = x & n350;
  assign n352 = r & n351;
  assign n353 = o & p;
  assign n354 = x & n353;
  assign n355 = ~o & ~p;
  assign n356 = ~a & ~n355;
  assign n357 = ~n354 & n356;
  assign n358 = ~n352 & n357;
  assign n359 = ~q & r;
  assign n360 = ~p & ~n359;
  assign n361 = ~m & n289;
  assign n362 = n288 & n360;
  assign n363 = n358 & n362;
  assign n364 = n288 & ~n361;
  assign n365 = n358 & n364;
  assign n366 = ~k & n288;
  assign n367 = n358 & n366;
  assign n368 = l & n288;
  assign n369 = n358 & n368;
  assign n370 = p & n360;
  assign n371 = n358 & n370;
  assign n372 = p & ~n361;
  assign n373 = n358 & n372;
  assign n374 = ~k & p;
  assign n375 = n358 & n374;
  assign n376 = l & p;
  assign n377 = n358 & n376;
  assign n378 = x & n360;
  assign n379 = n358 & n378;
  assign n380 = x & ~n361;
  assign n381 = n358 & n380;
  assign n382 = ~k & x;
  assign n383 = n358 & n382;
  assign n384 = l & x;
  assign n385 = n358 & n384;
  assign n386 = ~n383 & ~n385;
  assign n387 = ~n381 & n386;
  assign n388 = ~n379 & n387;
  assign n389 = ~n377 & n388;
  assign n390 = ~n375 & n389;
  assign n391 = ~n373 & n390;
  assign n392 = ~n371 & n391;
  assign n393 = ~n369 & n392;
  assign n394 = ~n367 & n393;
  assign n395 = ~n365 & n394;
  assign k0 = n363 | ~n395;
  assign n397 = ~p & ~q;
  assign n398 = ~o & ~q;
  assign n399 = ~a & ~n398;
  assign n400 = ~n397 & n399;
  assign n401 = n & n278;
  assign n402 = ~x & ~n401;
  assign n403 = n288 & n402;
  assign n404 = n400 & n403;
  assign n405 = x & n402;
  assign n406 = n400 & n405;
  assign n407 = q & n402;
  assign n408 = n400 & n407;
  assign n409 = ~q & n288;
  assign n410 = n400 & n409;
  assign n411 = ~p & n288;
  assign n412 = n400 & n411;
  assign n413 = ~o & n288;
  assign n414 = n400 & n413;
  assign n415 = ~q & x;
  assign n416 = n400 & n415;
  assign n417 = ~p & x;
  assign n418 = n400 & n417;
  assign n419 = n317 & n400;
  assign n420 = ~p & q;
  assign n421 = n400 & n420;
  assign n422 = ~o & q;
  assign n423 = n400 & n422;
  assign n424 = ~n421 & ~n423;
  assign n425 = ~n419 & n424;
  assign n426 = ~n418 & n425;
  assign n427 = ~n416 & n426;
  assign n428 = ~n414 & n427;
  assign n429 = ~n412 & n428;
  assign n430 = ~n410 & n429;
  assign n431 = ~n408 & n430;
  assign n432 = ~n406 & n431;
  assign l0 = n404 | ~n432;
  assign n434 = ~q & ~r;
  assign n435 = ~p & ~r;
  assign n436 = ~o & ~r;
  assign n437 = ~a & ~n436;
  assign n438 = ~n435 & n437;
  assign n439 = ~n434 & n438;
  assign n440 = p & q;
  assign n441 = r & n440;
  assign n442 = ~n397 & ~n441;
  assign n443 = ~x & ~n361;
  assign n444 = r & n443;
  assign n445 = n439 & n444;
  assign n446 = ~o & ~n361;
  assign n447 = r & n446;
  assign n448 = n439 & n447;
  assign n449 = r & n299;
  assign n450 = n439 & n449;
  assign n451 = r & n302;
  assign n452 = n439 & n451;
  assign n453 = r & n308;
  assign n454 = n439 & n453;
  assign n455 = r & n311;
  assign n456 = n439 & n455;
  assign n457 = ~x & n288;
  assign n458 = ~n361 & n457;
  assign n459 = n439 & n458;
  assign n460 = ~n361 & n413;
  assign n461 = n439 & n460;
  assign n462 = n317 & ~n361;
  assign n463 = n439 & n462;
  assign n464 = n300 & n439;
  assign n465 = n303 & n439;
  assign n466 = n309 & n439;
  assign n467 = n312 & n439;
  assign n468 = n331 & n439;
  assign n469 = n333 & n439;
  assign n470 = r & n442;
  assign n471 = n439 & n470;
  assign n472 = n288 & n442;
  assign n473 = n439 & n472;
  assign n474 = x & n442;
  assign n475 = n439 & n474;
  assign n476 = ~n473 & ~n475;
  assign n477 = ~n471 & n476;
  assign n478 = ~n469 & n477;
  assign n479 = ~n468 & n478;
  assign n480 = ~n467 & n479;
  assign n481 = ~n466 & n480;
  assign n482 = ~n465 & n481;
  assign n483 = ~n464 & n482;
  assign n484 = ~n463 & n483;
  assign n485 = ~n461 & n484;
  assign n486 = ~n459 & n485;
  assign n487 = ~n456 & n486;
  assign n488 = ~n454 & n487;
  assign n489 = ~n452 & n488;
  assign n490 = ~n450 & n489;
  assign n491 = ~n448 & n490;
  assign m0 = n445 | ~n491;
  assign n493 = o & ~p;
  assign n494 = n359 & n493;
  assign n495 = ~n402 & n494;
  assign n496 = r & s;
  assign n497 = ~q & n496;
  assign n498 = n402 & n495;
  assign n499 = ~a & n498;
  assign n500 = n495 & ~n497;
  assign n501 = ~a & n500;
  assign n502 = ~o & n495;
  assign n503 = ~a & n502;
  assign n504 = p & n495;
  assign n505 = ~a & n504;
  assign n506 = s & n402;
  assign n507 = ~a & n506;
  assign n508 = s & ~n497;
  assign n509 = ~a & n508;
  assign n510 = ~o & s;
  assign n511 = ~a & n510;
  assign n512 = p & s;
  assign n513 = ~a & n512;
  assign n514 = ~n511 & ~n513;
  assign n515 = ~n509 & n514;
  assign n516 = ~n507 & n515;
  assign n517 = ~n505 & n516;
  assign n518 = ~n503 & n517;
  assign n519 = ~n501 & n518;
  assign n0 = n499 | ~n519;
  assign n521 = ~x & ~n288;
  assign n522 = ~n63 & ~n521;
  assign n523 = s & ~t;
  assign n524 = r & n523;
  assign n525 = ~q & n524;
  assign n526 = o & n497;
  assign n527 = n411 & n526;
  assign n528 = n417 & n526;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~a & n493;
  assign n531 = n525 & n530;
  assign n532 = n522 & n531;
  assign n533 = ~a & t;
  assign n534 = n529 & n533;
  assign o0 = n532 | n534;
  assign n536 = ~n & ~x;
  assign n537 = ~n299 & ~n302;
  assign n538 = ~n296 & n537;
  assign n539 = ~n536 & n538;
  assign n540 = s & n127;
  assign n541 = r & n540;
  assign n542 = o & n397;
  assign n543 = r & n246;
  assign n544 = o & n543;
  assign n545 = ~q & n411;
  assign n546 = n544 & n545;
  assign n547 = ~q & n417;
  assign n548 = n544 & n547;
  assign n549 = ~n546 & ~n548;
  assign n550 = ~a & n542;
  assign n551 = n541 & n550;
  assign n552 = n539 & n551;
  assign n553 = ~a & u;
  assign n554 = n549 & n553;
  assign p0 = n552 | n554;
  assign n556 = t & n53;
  assign n557 = s & n556;
  assign n558 = ~p & n359;
  assign n559 = o & n558;
  assign n560 = r & n70;
  assign n561 = t & u;
  assign n562 = s & n561;
  assign n563 = r & n562;
  assign n564 = ~n560 & ~n563;
  assign n565 = o & ~n564;
  assign n566 = n545 & n565;
  assign n567 = n547 & n565;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~a & n539;
  assign n570 = n559 & n569;
  assign n571 = n557 & n570;
  assign n572 = ~a & v;
  assign n573 = n568 & n572;
  assign q0 = n571 | n573;
  assign n575 = ~t & u;
  assign n576 = ~s & n575;
  assign n577 = n120 & n576;
  assign n578 = ~n84 & n577;
  assign n579 = ~a & n578;
  assign n580 = ~s & n577;
  assign n581 = ~a & n580;
  assign n582 = t & n577;
  assign n583 = ~a & n582;
  assign n584 = ~u & n577;
  assign n585 = ~a & n584;
  assign n586 = ~a & n93;
  assign n587 = ~a & n95;
  assign n588 = ~a & n97;
  assign n589 = ~a & n99;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n587 & n590;
  assign n592 = ~n586 & n591;
  assign n593 = ~n585 & n592;
  assign n594 = ~n583 & n593;
  assign n595 = ~n581 & n594;
  assign r0 = n579 | ~n595;
  assign n597 = ~a & b;
  assign n598 = ~x & n597;
  assign n599 = ~a & ~b;
  assign n600 = x & n599;
  assign s0 = n598 | n600;
  assign n602 = ~a & c;
  assign n603 = ~y & n602;
  assign n604 = ~a & ~c;
  assign n605 = y & n604;
  assign t0 = n603 | n605;
endmodule


