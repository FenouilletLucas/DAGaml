// Benchmark "rca_256" written by ABC on Sat Apr 23 20:18:09 2016

module rca_256 ( 
    a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7, a8, b8,
    a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15, b15,
    a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22, b22,
    a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29, b29,
    a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36, b36,
    a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43, b43,
    a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50, b50,
    a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57, b57,
    a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64, b64,
    a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71, b71,
    a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78, b78,
    a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85, b85,
    a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92, b92,
    a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99, b99,
    a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105, b105,
    a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111, b111,
    a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117, b117,
    a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123, b123,
    a124, b124, a125, b125, a126, b126, a127, b127, a128, b128, a129, b129,
    a130, b130, a131, b131, a132, b132, a133, b133, a134, b134, a135, b135,
    a136, b136, a137, b137, a138, b138, a139, b139, a140, b140, a141, b141,
    a142, b142, a143, b143, a144, b144, a145, b145, a146, b146, a147, b147,
    a148, b148, a149, b149, a150, b150, a151, b151, a152, b152, a153, b153,
    a154, b154, a155, b155, a156, b156, a157, b157, a158, b158, a159, b159,
    a160, b160, a161, b161, a162, b162, a163, b163, a164, b164, a165, b165,
    a166, b166, a167, b167, a168, b168, a169, b169, a170, b170, a171, b171,
    a172, b172, a173, b173, a174, b174, a175, b175, a176, b176, a177, b177,
    a178, b178, a179, b179, a180, b180, a181, b181, a182, b182, a183, b183,
    a184, b184, a185, b185, a186, b186, a187, b187, a188, b188, a189, b189,
    a190, b190, a191, b191, a192, b192, a193, b193, a194, b194, a195, b195,
    a196, b196, a197, b197, a198, b198, a199, b199, a200, b200, a201, b201,
    a202, b202, a203, b203, a204, b204, a205, b205, a206, b206, a207, b207,
    a208, b208, a209, b209, a210, b210, a211, b211, a212, b212, a213, b213,
    a214, b214, a215, b215, a216, b216, a217, b217, a218, b218, a219, b219,
    a220, b220, a221, b221, a222, b222, a223, b223, a224, b224, a225, b225,
    a226, b226, a227, b227, a228, b228, a229, b229, a230, b230, a231, b231,
    a232, b232, a233, b233, a234, b234, a235, b235, a236, b236, a237, b237,
    a238, b238, a239, b239, a240, b240, a241, b241, a242, b242, a243, b243,
    a244, b244, a245, b245, a246, b246, a247, b247, a248, b248, a249, b249,
    a250, b250, a251, b251, a252, b252, a253, b253, a254, b254, a255, b255,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128, s129, s130, s131, s132, s133, s134, s135,
    s136, s137, s138, s139, s140, s141, s142, s143, s144, s145, s146, s147,
    s148, s149, s150, s151, s152, s153, s154, s155, s156, s157, s158, s159,
    s160, s161, s162, s163, s164, s165, s166, s167, s168, s169, s170, s171,
    s172, s173, s174, s175, s176, s177, s178, s179, s180, s181, s182, s183,
    s184, s185, s186, s187, s188, s189, s190, s191, s192, s193, s194, s195,
    s196, s197, s198, s199, s200, s201, s202, s203, s204, s205, s206, s207,
    s208, s209, s210, s211, s212, s213, s214, s215, s216, s217, s218, s219,
    s220, s221, s222, s223, s224, s225, s226, s227, s228, s229, s230, s231,
    s232, s233, s234, s235, s236, s237, s238, s239, s240, s241, s242, s243,
    s244, s245, s246, s247, s248, s249, s250, s251, s252, s253, s254, s255,
    s256  );
  input  a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7,
    a8, b8, a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15,
    b15, a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22,
    b22, a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29,
    b29, a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36,
    b36, a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43,
    b43, a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50,
    b50, a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57,
    b57, a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64,
    b64, a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71,
    b71, a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78,
    b78, a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85,
    b85, a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92,
    b92, a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99,
    b99, a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105,
    b105, a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111,
    b111, a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117,
    b117, a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123,
    b123, a124, b124, a125, b125, a126, b126, a127, b127, a128, b128, a129,
    b129, a130, b130, a131, b131, a132, b132, a133, b133, a134, b134, a135,
    b135, a136, b136, a137, b137, a138, b138, a139, b139, a140, b140, a141,
    b141, a142, b142, a143, b143, a144, b144, a145, b145, a146, b146, a147,
    b147, a148, b148, a149, b149, a150, b150, a151, b151, a152, b152, a153,
    b153, a154, b154, a155, b155, a156, b156, a157, b157, a158, b158, a159,
    b159, a160, b160, a161, b161, a162, b162, a163, b163, a164, b164, a165,
    b165, a166, b166, a167, b167, a168, b168, a169, b169, a170, b170, a171,
    b171, a172, b172, a173, b173, a174, b174, a175, b175, a176, b176, a177,
    b177, a178, b178, a179, b179, a180, b180, a181, b181, a182, b182, a183,
    b183, a184, b184, a185, b185, a186, b186, a187, b187, a188, b188, a189,
    b189, a190, b190, a191, b191, a192, b192, a193, b193, a194, b194, a195,
    b195, a196, b196, a197, b197, a198, b198, a199, b199, a200, b200, a201,
    b201, a202, b202, a203, b203, a204, b204, a205, b205, a206, b206, a207,
    b207, a208, b208, a209, b209, a210, b210, a211, b211, a212, b212, a213,
    b213, a214, b214, a215, b215, a216, b216, a217, b217, a218, b218, a219,
    b219, a220, b220, a221, b221, a222, b222, a223, b223, a224, b224, a225,
    b225, a226, b226, a227, b227, a228, b228, a229, b229, a230, b230, a231,
    b231, a232, b232, a233, b233, a234, b234, a235, b235, a236, b236, a237,
    b237, a238, b238, a239, b239, a240, b240, a241, b241, a242, b242, a243,
    b243, a244, b244, a245, b245, a246, b246, a247, b247, a248, b248, a249,
    b249, a250, b250, a251, b251, a252, b252, a253, b253, a254, b254, a255,
    b255;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128, s129, s130, s131, s132, s133, s134, s135,
    s136, s137, s138, s139, s140, s141, s142, s143, s144, s145, s146, s147,
    s148, s149, s150, s151, s152, s153, s154, s155, s156, s157, s158, s159,
    s160, s161, s162, s163, s164, s165, s166, s167, s168, s169, s170, s171,
    s172, s173, s174, s175, s176, s177, s178, s179, s180, s181, s182, s183,
    s184, s185, s186, s187, s188, s189, s190, s191, s192, s193, s194, s195,
    s196, s197, s198, s199, s200, s201, s202, s203, s204, s205, s206, s207,
    s208, s209, s210, s211, s212, s213, s214, s215, s216, s217, s218, s219,
    s220, s221, s222, s223, s224, s225, s226, s227, s228, s229, s230, s231,
    s232, s233, s234, s235, s236, s237, s238, s239, s240, s241, s242, s243,
    s244, s245, s246, s247, s248, s249, s250, s251, s252, s253, s254, s255,
    s256;
  wire n770, n771, n773, n774, n775, n776, n777, n779, n780, n781, n782,
    n783, n784, n786, n787, n788, n789, n790, n791, n793, n794, n795, n796,
    n797, n798, n800, n801, n802, n803, n804, n805, n807, n808, n809, n810,
    n811, n812, n814, n815, n816, n817, n818, n819, n821, n822, n823, n824,
    n825, n826, n828, n829, n830, n831, n832, n833, n835, n836, n837, n838,
    n839, n840, n842, n843, n844, n845, n846, n847, n849, n850, n851, n852,
    n853, n854, n856, n857, n858, n859, n860, n861, n863, n864, n865, n866,
    n867, n868, n870, n871, n872, n873, n874, n875, n877, n878, n879, n880,
    n881, n882, n884, n885, n886, n887, n888, n889, n891, n892, n893, n894,
    n895, n896, n898, n899, n900, n901, n902, n903, n905, n906, n907, n908,
    n909, n910, n912, n913, n914, n915, n916, n917, n919, n920, n921, n922,
    n923, n924, n926, n927, n928, n929, n930, n931, n933, n934, n935, n936,
    n937, n938, n940, n941, n942, n943, n944, n945, n947, n948, n949, n950,
    n951, n952, n954, n955, n956, n957, n958, n959, n961, n962, n963, n964,
    n965, n966, n968, n969, n970, n971, n972, n973, n975, n976, n977, n978,
    n979, n980, n982, n983, n984, n985, n986, n987, n989, n990, n991, n992,
    n993, n994, n996, n997, n998, n999, n1000, n1001, n1003, n1004, n1005,
    n1006, n1007, n1008, n1010, n1011, n1012, n1013, n1014, n1015, n1017,
    n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028,
    n1029, n1031, n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1040,
    n1041, n1042, n1043, n1045, n1046, n1047, n1048, n1049, n1050, n1052,
    n1053, n1054, n1055, n1056, n1057, n1059, n1060, n1061, n1062, n1063,
    n1064, n1066, n1067, n1068, n1069, n1070, n1071, n1073, n1074, n1075,
    n1076, n1077, n1078, n1080, n1081, n1082, n1083, n1084, n1085, n1087,
    n1088, n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1097, n1098,
    n1099, n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109, n1110,
    n1111, n1112, n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1122,
    n1123, n1124, n1125, n1126, n1127, n1129, n1130, n1131, n1132, n1133,
    n1134, n1136, n1137, n1138, n1139, n1140, n1141, n1143, n1144, n1145,
    n1146, n1147, n1148, n1150, n1151, n1152, n1153, n1154, n1155, n1157,
    n1158, n1159, n1160, n1161, n1162, n1164, n1165, n1166, n1167, n1168,
    n1169, n1171, n1172, n1173, n1174, n1175, n1176, n1178, n1179, n1180,
    n1181, n1182, n1183, n1185, n1186, n1187, n1188, n1189, n1190, n1192,
    n1193, n1194, n1195, n1196, n1197, n1199, n1200, n1201, n1202, n1203,
    n1204, n1206, n1207, n1208, n1209, n1210, n1211, n1213, n1214, n1215,
    n1216, n1217, n1218, n1220, n1221, n1222, n1223, n1224, n1225, n1227,
    n1228, n1229, n1230, n1231, n1232, n1234, n1235, n1236, n1237, n1238,
    n1239, n1241, n1242, n1243, n1244, n1245, n1246, n1248, n1249, n1250,
    n1251, n1252, n1253, n1255, n1256, n1257, n1258, n1259, n1260, n1262,
    n1263, n1264, n1265, n1266, n1267, n1269, n1270, n1271, n1272, n1273,
    n1274, n1276, n1277, n1278, n1279, n1280, n1281, n1283, n1284, n1285,
    n1286, n1287, n1288, n1290, n1291, n1292, n1293, n1294, n1295, n1297,
    n1298, n1299, n1300, n1301, n1302, n1304, n1305, n1306, n1307, n1308,
    n1309, n1311, n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320,
    n1321, n1322, n1323, n1325, n1326, n1327, n1328, n1329, n1330, n1332,
    n1333, n1334, n1335, n1336, n1337, n1339, n1340, n1341, n1342, n1343,
    n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1353, n1354, n1355,
    n1356, n1357, n1358, n1360, n1361, n1362, n1363, n1364, n1365, n1367,
    n1368, n1369, n1370, n1371, n1372, n1374, n1375, n1376, n1377, n1378,
    n1379, n1381, n1382, n1383, n1384, n1385, n1386, n1388, n1389, n1390,
    n1391, n1392, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1402,
    n1403, n1404, n1405, n1406, n1407, n1409, n1410, n1411, n1412, n1413,
    n1414, n1416, n1417, n1418, n1419, n1420, n1421, n1423, n1424, n1425,
    n1426, n1427, n1428, n1430, n1431, n1432, n1433, n1434, n1435, n1437,
    n1438, n1439, n1440, n1441, n1442, n1444, n1445, n1446, n1447, n1448,
    n1449, n1451, n1452, n1453, n1454, n1455, n1456, n1458, n1459, n1460,
    n1461, n1462, n1463, n1465, n1466, n1467, n1468, n1469, n1470, n1472,
    n1473, n1474, n1475, n1476, n1477, n1479, n1480, n1481, n1482, n1483,
    n1484, n1486, n1487, n1488, n1489, n1490, n1491, n1493, n1494, n1495,
    n1496, n1497, n1498, n1500, n1501, n1502, n1503, n1504, n1505, n1507,
    n1508, n1509, n1510, n1511, n1512, n1514, n1515, n1516, n1517, n1518,
    n1519, n1521, n1522, n1523, n1524, n1525, n1526, n1528, n1529, n1530,
    n1531, n1532, n1533, n1535, n1536, n1537, n1538, n1539, n1540, n1542,
    n1543, n1544, n1545, n1546, n1547, n1549, n1550, n1551, n1552, n1553,
    n1554, n1556, n1557, n1558, n1559, n1560, n1561, n1563, n1564, n1565,
    n1566, n1567, n1568, n1570, n1571, n1572, n1573, n1574, n1575, n1577,
    n1578, n1579, n1580, n1581, n1582, n1584, n1585, n1586, n1587, n1588,
    n1589, n1591, n1592, n1593, n1594, n1595, n1596, n1598, n1599, n1600,
    n1601, n1602, n1603, n1605, n1606, n1607, n1608, n1609, n1610, n1612,
    n1613, n1614, n1615, n1616, n1617, n1619, n1620, n1621, n1622, n1623,
    n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1633, n1634, n1635,
    n1636, n1637, n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1647,
    n1648, n1649, n1650, n1651, n1652, n1654, n1655, n1656, n1657, n1658,
    n1659, n1661, n1662, n1663, n1664, n1665, n1666, n1668, n1669, n1670,
    n1671, n1672, n1673, n1675, n1676, n1677, n1678, n1679, n1680, n1682,
    n1683, n1684, n1685, n1686, n1687, n1689, n1690, n1691, n1692, n1693,
    n1694, n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704, n1705,
    n1706, n1707, n1708, n1710, n1711, n1712, n1713, n1714, n1715, n1717,
    n1718, n1719, n1720, n1721, n1722, n1724, n1725, n1726, n1727, n1728,
    n1729, n1731, n1732, n1733, n1734, n1735, n1736, n1738, n1739, n1740,
    n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1749, n1750, n1752,
    n1753, n1754, n1755, n1756, n1757, n1759, n1760, n1761, n1762, n1763,
    n1764, n1766, n1767, n1768, n1769, n1770, n1771, n1773, n1774, n1775,
    n1776, n1777, n1778, n1780, n1781, n1782, n1783, n1784, n1785, n1787,
    n1788, n1789, n1790, n1791, n1792, n1794, n1795, n1796, n1797, n1798,
    n1799, n1801, n1802, n1803, n1804, n1805, n1806, n1808, n1809, n1810,
    n1811, n1812, n1813, n1815, n1816, n1817, n1818, n1819, n1820, n1822,
    n1823, n1824, n1825, n1826, n1827, n1829, n1830, n1831, n1832, n1833,
    n1834, n1836, n1837, n1838, n1839, n1840, n1841, n1843, n1844, n1845,
    n1846, n1847, n1848, n1850, n1851, n1852, n1853, n1854, n1855, n1857,
    n1858, n1859, n1860, n1861, n1862, n1864, n1865, n1866, n1867, n1868,
    n1869, n1871, n1872, n1873, n1874, n1875, n1876, n1878, n1879, n1880,
    n1881, n1882, n1883, n1885, n1886, n1887, n1888, n1889, n1890, n1892,
    n1893, n1894, n1895, n1896, n1897, n1899, n1900, n1901, n1902, n1903,
    n1904, n1906, n1907, n1908, n1909, n1910, n1911, n1913, n1914, n1915,
    n1916, n1917, n1918, n1920, n1921, n1922, n1923, n1924, n1925, n1927,
    n1928, n1929, n1930, n1931, n1932, n1934, n1935, n1936, n1937, n1938,
    n1939, n1941, n1942, n1943, n1944, n1945, n1946, n1948, n1949, n1950,
    n1951, n1952, n1953, n1955, n1956, n1957, n1958, n1959, n1960, n1962,
    n1963, n1964, n1965, n1966, n1967, n1969, n1970, n1971, n1972, n1973,
    n1974, n1976, n1977, n1978, n1979, n1980, n1981, n1983, n1984, n1985,
    n1986, n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1995, n1997,
    n1998, n1999, n2000, n2001, n2002, n2004, n2005, n2006, n2007, n2008,
    n2009, n2011, n2012, n2013, n2014, n2015, n2016, n2018, n2019, n2020,
    n2021, n2022, n2023, n2025, n2026, n2027, n2028, n2029, n2030, n2032,
    n2033, n2034, n2035, n2036, n2037, n2039, n2040, n2041, n2042, n2043,
    n2044, n2046, n2047, n2048, n2049, n2050, n2051, n2053, n2054, n2055,
    n2056, n2057, n2058, n2060, n2061, n2062, n2063, n2064, n2065, n2067,
    n2068, n2069, n2070, n2071, n2072, n2074, n2075, n2076, n2077, n2078,
    n2079, n2081, n2082, n2083, n2084, n2085, n2086, n2088, n2089, n2090,
    n2091, n2092, n2093, n2095, n2096, n2097, n2098, n2099, n2100, n2102,
    n2103, n2104, n2105, n2106, n2107, n2109, n2110, n2111, n2112, n2113,
    n2114, n2116, n2117, n2118, n2119, n2120, n2121, n2123, n2124, n2125,
    n2126, n2127, n2128, n2130, n2131, n2132, n2133, n2134, n2135, n2137,
    n2138, n2139, n2140, n2141, n2142, n2144, n2145, n2146, n2147, n2148,
    n2149, n2151, n2152, n2153, n2154, n2155, n2156, n2158, n2159, n2160,
    n2161, n2162, n2163, n2165, n2166, n2167, n2168, n2169, n2170, n2172,
    n2173, n2174, n2175, n2176, n2177, n2179, n2180, n2181, n2182, n2183,
    n2184, n2186, n2187, n2188, n2189, n2190, n2191, n2193, n2194, n2195,
    n2196, n2197, n2198, n2200, n2201, n2202, n2203, n2204, n2205, n2207,
    n2208, n2209, n2210, n2211, n2212, n2214, n2215, n2216, n2217, n2218,
    n2219, n2221, n2222, n2223, n2224, n2225, n2226, n2228, n2229, n2230,
    n2231, n2232, n2233, n2235, n2236, n2237, n2238, n2239, n2240, n2242,
    n2243, n2244, n2245, n2246, n2247, n2249, n2250, n2251, n2252, n2253,
    n2254, n2256, n2257, n2258, n2259, n2260, n2261, n2263, n2264, n2265,
    n2266, n2267, n2268, n2270, n2271, n2272, n2273, n2274, n2275, n2277,
    n2278, n2279, n2280, n2281, n2282, n2284, n2285, n2286, n2287, n2288,
    n2289, n2291, n2292, n2293, n2294, n2295, n2296, n2298, n2299, n2300,
    n2301, n2302, n2303, n2305, n2306, n2307, n2308, n2309, n2310, n2312,
    n2313, n2314, n2315, n2316, n2317, n2319, n2320, n2321, n2322, n2323,
    n2324, n2326, n2327, n2328, n2329, n2330, n2331, n2333, n2334, n2335,
    n2336, n2337, n2338, n2340, n2341, n2342, n2343, n2344, n2345, n2347,
    n2348, n2349, n2350, n2351, n2352, n2354, n2355, n2356, n2357, n2358,
    n2359, n2361, n2362, n2363, n2364, n2365, n2366, n2368, n2369, n2370,
    n2371, n2372, n2373, n2375, n2376, n2377, n2378, n2379, n2380, n2382,
    n2383, n2384, n2385, n2386, n2387, n2389, n2390, n2391, n2392, n2393,
    n2394, n2396, n2397, n2398, n2399, n2400, n2401, n2403, n2404, n2405,
    n2406, n2407, n2408, n2410, n2411, n2412, n2413, n2414, n2415, n2417,
    n2418, n2419, n2420, n2421, n2422, n2424, n2425, n2426, n2427, n2428,
    n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2438, n2439, n2440,
    n2441, n2442, n2443, n2445, n2446, n2447, n2448, n2449, n2450, n2452,
    n2453, n2454, n2455, n2456, n2457, n2459, n2460, n2461, n2462, n2463,
    n2464, n2466, n2467, n2468, n2469, n2470, n2471, n2473, n2474, n2475,
    n2476, n2477, n2478, n2480, n2481, n2482, n2483, n2484, n2485, n2487,
    n2488, n2489, n2490, n2491, n2492, n2494, n2495, n2496, n2497, n2498,
    n2499, n2501, n2502, n2503, n2504, n2505, n2506, n2508, n2509, n2510,
    n2511, n2512, n2513, n2515, n2516, n2517, n2518, n2519, n2520, n2522,
    n2523, n2524, n2525, n2526, n2527, n2529, n2530, n2531, n2532, n2533,
    n2534, n2536, n2537, n2538, n2539, n2540, n2541, n2543, n2544, n2545,
    n2546, n2547, n2548, n2550, n2551, n2552, n2553, n2554, n2555;
  assign n770 = a0 & b0;
  assign n771 = ~a0 & ~b0;
  assign s0 = ~n770 & ~n771;
  assign n773 = a1 & b1;
  assign n774 = ~a1 & ~b1;
  assign n775 = ~n773 & ~n774;
  assign n776 = n770 & n775;
  assign n777 = ~n770 & ~n775;
  assign s1 = ~n776 & ~n777;
  assign n779 = ~n773 & ~n776;
  assign n780 = a2 & b2;
  assign n781 = ~a2 & ~b2;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n779 & n782;
  assign n784 = n779 & ~n782;
  assign s2 = ~n783 & ~n784;
  assign n786 = ~n780 & ~n783;
  assign n787 = a3 & b3;
  assign n788 = ~a3 & ~b3;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~n786 & n789;
  assign n791 = n786 & ~n789;
  assign s3 = ~n790 & ~n791;
  assign n793 = ~n787 & ~n790;
  assign n794 = a4 & b4;
  assign n795 = ~a4 & ~b4;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~n793 & n796;
  assign n798 = n793 & ~n796;
  assign s4 = ~n797 & ~n798;
  assign n800 = ~n794 & ~n797;
  assign n801 = a5 & b5;
  assign n802 = ~a5 & ~b5;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n800 & n803;
  assign n805 = n800 & ~n803;
  assign s5 = ~n804 & ~n805;
  assign n807 = ~n801 & ~n804;
  assign n808 = a6 & b6;
  assign n809 = ~a6 & ~b6;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n807 & n810;
  assign n812 = n807 & ~n810;
  assign s6 = ~n811 & ~n812;
  assign n814 = ~n808 & ~n811;
  assign n815 = a7 & b7;
  assign n816 = ~a7 & ~b7;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~n814 & n817;
  assign n819 = n814 & ~n817;
  assign s7 = ~n818 & ~n819;
  assign n821 = ~n815 & ~n818;
  assign n822 = a8 & b8;
  assign n823 = ~a8 & ~b8;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n821 & n824;
  assign n826 = n821 & ~n824;
  assign s8 = ~n825 & ~n826;
  assign n828 = ~n822 & ~n825;
  assign n829 = a9 & b9;
  assign n830 = ~a9 & ~b9;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n828 & n831;
  assign n833 = n828 & ~n831;
  assign s9 = ~n832 & ~n833;
  assign n835 = ~n829 & ~n832;
  assign n836 = a10 & b10;
  assign n837 = ~a10 & ~b10;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n835 & n838;
  assign n840 = n835 & ~n838;
  assign s10 = ~n839 & ~n840;
  assign n842 = ~n836 & ~n839;
  assign n843 = a11 & b11;
  assign n844 = ~a11 & ~b11;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n842 & n845;
  assign n847 = n842 & ~n845;
  assign s11 = ~n846 & ~n847;
  assign n849 = ~n843 & ~n846;
  assign n850 = a12 & b12;
  assign n851 = ~a12 & ~b12;
  assign n852 = ~n850 & ~n851;
  assign n853 = ~n849 & n852;
  assign n854 = n849 & ~n852;
  assign s12 = ~n853 & ~n854;
  assign n856 = ~n850 & ~n853;
  assign n857 = a13 & b13;
  assign n858 = ~a13 & ~b13;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n856 & n859;
  assign n861 = n856 & ~n859;
  assign s13 = ~n860 & ~n861;
  assign n863 = ~n857 & ~n860;
  assign n864 = a14 & b14;
  assign n865 = ~a14 & ~b14;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n863 & n866;
  assign n868 = n863 & ~n866;
  assign s14 = ~n867 & ~n868;
  assign n870 = ~n864 & ~n867;
  assign n871 = a15 & b15;
  assign n872 = ~a15 & ~b15;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n870 & n873;
  assign n875 = n870 & ~n873;
  assign s15 = ~n874 & ~n875;
  assign n877 = ~n871 & ~n874;
  assign n878 = a16 & b16;
  assign n879 = ~a16 & ~b16;
  assign n880 = ~n878 & ~n879;
  assign n881 = ~n877 & n880;
  assign n882 = n877 & ~n880;
  assign s16 = ~n881 & ~n882;
  assign n884 = ~n878 & ~n881;
  assign n885 = a17 & b17;
  assign n886 = ~a17 & ~b17;
  assign n887 = ~n885 & ~n886;
  assign n888 = ~n884 & n887;
  assign n889 = n884 & ~n887;
  assign s17 = ~n888 & ~n889;
  assign n891 = ~n885 & ~n888;
  assign n892 = a18 & b18;
  assign n893 = ~a18 & ~b18;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n891 & n894;
  assign n896 = n891 & ~n894;
  assign s18 = ~n895 & ~n896;
  assign n898 = ~n892 & ~n895;
  assign n899 = a19 & b19;
  assign n900 = ~a19 & ~b19;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n898 & n901;
  assign n903 = n898 & ~n901;
  assign s19 = ~n902 & ~n903;
  assign n905 = ~n899 & ~n902;
  assign n906 = a20 & b20;
  assign n907 = ~a20 & ~b20;
  assign n908 = ~n906 & ~n907;
  assign n909 = ~n905 & n908;
  assign n910 = n905 & ~n908;
  assign s20 = ~n909 & ~n910;
  assign n912 = ~n906 & ~n909;
  assign n913 = a21 & b21;
  assign n914 = ~a21 & ~b21;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n912 & n915;
  assign n917 = n912 & ~n915;
  assign s21 = ~n916 & ~n917;
  assign n919 = ~n913 & ~n916;
  assign n920 = a22 & b22;
  assign n921 = ~a22 & ~b22;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n919 & n922;
  assign n924 = n919 & ~n922;
  assign s22 = ~n923 & ~n924;
  assign n926 = ~n920 & ~n923;
  assign n927 = a23 & b23;
  assign n928 = ~a23 & ~b23;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n926 & n929;
  assign n931 = n926 & ~n929;
  assign s23 = ~n930 & ~n931;
  assign n933 = ~n927 & ~n930;
  assign n934 = a24 & b24;
  assign n935 = ~a24 & ~b24;
  assign n936 = ~n934 & ~n935;
  assign n937 = ~n933 & n936;
  assign n938 = n933 & ~n936;
  assign s24 = ~n937 & ~n938;
  assign n940 = ~n934 & ~n937;
  assign n941 = a25 & b25;
  assign n942 = ~a25 & ~b25;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n940 & n943;
  assign n945 = n940 & ~n943;
  assign s25 = ~n944 & ~n945;
  assign n947 = ~n941 & ~n944;
  assign n948 = a26 & b26;
  assign n949 = ~a26 & ~b26;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n947 & n950;
  assign n952 = n947 & ~n950;
  assign s26 = ~n951 & ~n952;
  assign n954 = ~n948 & ~n951;
  assign n955 = a27 & b27;
  assign n956 = ~a27 & ~b27;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n954 & n957;
  assign n959 = n954 & ~n957;
  assign s27 = ~n958 & ~n959;
  assign n961 = ~n955 & ~n958;
  assign n962 = a28 & b28;
  assign n963 = ~a28 & ~b28;
  assign n964 = ~n962 & ~n963;
  assign n965 = ~n961 & n964;
  assign n966 = n961 & ~n964;
  assign s28 = ~n965 & ~n966;
  assign n968 = ~n962 & ~n965;
  assign n969 = a29 & b29;
  assign n970 = ~a29 & ~b29;
  assign n971 = ~n969 & ~n970;
  assign n972 = ~n968 & n971;
  assign n973 = n968 & ~n971;
  assign s29 = ~n972 & ~n973;
  assign n975 = ~n969 & ~n972;
  assign n976 = a30 & b30;
  assign n977 = ~a30 & ~b30;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n975 & n978;
  assign n980 = n975 & ~n978;
  assign s30 = ~n979 & ~n980;
  assign n982 = ~n976 & ~n979;
  assign n983 = a31 & b31;
  assign n984 = ~a31 & ~b31;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n982 & n985;
  assign n987 = n982 & ~n985;
  assign s31 = ~n986 & ~n987;
  assign n989 = ~n983 & ~n986;
  assign n990 = a32 & b32;
  assign n991 = ~a32 & ~b32;
  assign n992 = ~n990 & ~n991;
  assign n993 = ~n989 & n992;
  assign n994 = n989 & ~n992;
  assign s32 = ~n993 & ~n994;
  assign n996 = ~n990 & ~n993;
  assign n997 = a33 & b33;
  assign n998 = ~a33 & ~b33;
  assign n999 = ~n997 & ~n998;
  assign n1000 = ~n996 & n999;
  assign n1001 = n996 & ~n999;
  assign s33 = ~n1000 & ~n1001;
  assign n1003 = ~n997 & ~n1000;
  assign n1004 = a34 & b34;
  assign n1005 = ~a34 & ~b34;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1003 & n1006;
  assign n1008 = n1003 & ~n1006;
  assign s34 = ~n1007 & ~n1008;
  assign n1010 = ~n1004 & ~n1007;
  assign n1011 = a35 & b35;
  assign n1012 = ~a35 & ~b35;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1010 & n1013;
  assign n1015 = n1010 & ~n1013;
  assign s35 = ~n1014 & ~n1015;
  assign n1017 = ~n1011 & ~n1014;
  assign n1018 = a36 & b36;
  assign n1019 = ~a36 & ~b36;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~n1017 & n1020;
  assign n1022 = n1017 & ~n1020;
  assign s36 = ~n1021 & ~n1022;
  assign n1024 = ~n1018 & ~n1021;
  assign n1025 = a37 & b37;
  assign n1026 = ~a37 & ~b37;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~n1024 & n1027;
  assign n1029 = n1024 & ~n1027;
  assign s37 = ~n1028 & ~n1029;
  assign n1031 = ~n1025 & ~n1028;
  assign n1032 = a38 & b38;
  assign n1033 = ~a38 & ~b38;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1031 & n1034;
  assign n1036 = n1031 & ~n1034;
  assign s38 = ~n1035 & ~n1036;
  assign n1038 = ~n1032 & ~n1035;
  assign n1039 = a39 & b39;
  assign n1040 = ~a39 & ~b39;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = ~n1038 & n1041;
  assign n1043 = n1038 & ~n1041;
  assign s39 = ~n1042 & ~n1043;
  assign n1045 = ~n1039 & ~n1042;
  assign n1046 = a40 & b40;
  assign n1047 = ~a40 & ~b40;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1045 & n1048;
  assign n1050 = n1045 & ~n1048;
  assign s40 = ~n1049 & ~n1050;
  assign n1052 = ~n1046 & ~n1049;
  assign n1053 = a41 & b41;
  assign n1054 = ~a41 & ~b41;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1052 & n1055;
  assign n1057 = n1052 & ~n1055;
  assign s41 = ~n1056 & ~n1057;
  assign n1059 = ~n1053 & ~n1056;
  assign n1060 = a42 & b42;
  assign n1061 = ~a42 & ~b42;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1059 & n1062;
  assign n1064 = n1059 & ~n1062;
  assign s42 = ~n1063 & ~n1064;
  assign n1066 = ~n1060 & ~n1063;
  assign n1067 = a43 & b43;
  assign n1068 = ~a43 & ~b43;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~n1066 & n1069;
  assign n1071 = n1066 & ~n1069;
  assign s43 = ~n1070 & ~n1071;
  assign n1073 = ~n1067 & ~n1070;
  assign n1074 = a44 & b44;
  assign n1075 = ~a44 & ~b44;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = ~n1073 & n1076;
  assign n1078 = n1073 & ~n1076;
  assign s44 = ~n1077 & ~n1078;
  assign n1080 = ~n1074 & ~n1077;
  assign n1081 = a45 & b45;
  assign n1082 = ~a45 & ~b45;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1080 & n1083;
  assign n1085 = n1080 & ~n1083;
  assign s45 = ~n1084 & ~n1085;
  assign n1087 = ~n1081 & ~n1084;
  assign n1088 = a46 & b46;
  assign n1089 = ~a46 & ~b46;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~n1087 & n1090;
  assign n1092 = n1087 & ~n1090;
  assign s46 = ~n1091 & ~n1092;
  assign n1094 = ~n1088 & ~n1091;
  assign n1095 = a47 & b47;
  assign n1096 = ~a47 & ~b47;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n1094 & n1097;
  assign n1099 = n1094 & ~n1097;
  assign s47 = ~n1098 & ~n1099;
  assign n1101 = ~n1095 & ~n1098;
  assign n1102 = a48 & b48;
  assign n1103 = ~a48 & ~b48;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n1101 & n1104;
  assign n1106 = n1101 & ~n1104;
  assign s48 = ~n1105 & ~n1106;
  assign n1108 = ~n1102 & ~n1105;
  assign n1109 = a49 & b49;
  assign n1110 = ~a49 & ~b49;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1108 & n1111;
  assign n1113 = n1108 & ~n1111;
  assign s49 = ~n1112 & ~n1113;
  assign n1115 = ~n1109 & ~n1112;
  assign n1116 = a50 & b50;
  assign n1117 = ~a50 & ~b50;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1115 & n1118;
  assign n1120 = n1115 & ~n1118;
  assign s50 = ~n1119 & ~n1120;
  assign n1122 = ~n1116 & ~n1119;
  assign n1123 = a51 & b51;
  assign n1124 = ~a51 & ~b51;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1122 & n1125;
  assign n1127 = n1122 & ~n1125;
  assign s51 = ~n1126 & ~n1127;
  assign n1129 = ~n1123 & ~n1126;
  assign n1130 = a52 & b52;
  assign n1131 = ~a52 & ~b52;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1129 & n1132;
  assign n1134 = n1129 & ~n1132;
  assign s52 = ~n1133 & ~n1134;
  assign n1136 = ~n1130 & ~n1133;
  assign n1137 = a53 & b53;
  assign n1138 = ~a53 & ~b53;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1136 & n1139;
  assign n1141 = n1136 & ~n1139;
  assign s53 = ~n1140 & ~n1141;
  assign n1143 = ~n1137 & ~n1140;
  assign n1144 = a54 & b54;
  assign n1145 = ~a54 & ~b54;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1143 & n1146;
  assign n1148 = n1143 & ~n1146;
  assign s54 = ~n1147 & ~n1148;
  assign n1150 = ~n1144 & ~n1147;
  assign n1151 = a55 & b55;
  assign n1152 = ~a55 & ~b55;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1150 & n1153;
  assign n1155 = n1150 & ~n1153;
  assign s55 = ~n1154 & ~n1155;
  assign n1157 = ~n1151 & ~n1154;
  assign n1158 = a56 & b56;
  assign n1159 = ~a56 & ~b56;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1157 & n1160;
  assign n1162 = n1157 & ~n1160;
  assign s56 = ~n1161 & ~n1162;
  assign n1164 = ~n1158 & ~n1161;
  assign n1165 = a57 & b57;
  assign n1166 = ~a57 & ~b57;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1164 & n1167;
  assign n1169 = n1164 & ~n1167;
  assign s57 = ~n1168 & ~n1169;
  assign n1171 = ~n1165 & ~n1168;
  assign n1172 = a58 & b58;
  assign n1173 = ~a58 & ~b58;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1171 & n1174;
  assign n1176 = n1171 & ~n1174;
  assign s58 = ~n1175 & ~n1176;
  assign n1178 = ~n1172 & ~n1175;
  assign n1179 = a59 & b59;
  assign n1180 = ~a59 & ~b59;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1178 & n1181;
  assign n1183 = n1178 & ~n1181;
  assign s59 = ~n1182 & ~n1183;
  assign n1185 = ~n1179 & ~n1182;
  assign n1186 = a60 & b60;
  assign n1187 = ~a60 & ~b60;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n1185 & n1188;
  assign n1190 = n1185 & ~n1188;
  assign s60 = ~n1189 & ~n1190;
  assign n1192 = ~n1186 & ~n1189;
  assign n1193 = a61 & b61;
  assign n1194 = ~a61 & ~b61;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = ~n1192 & n1195;
  assign n1197 = n1192 & ~n1195;
  assign s61 = ~n1196 & ~n1197;
  assign n1199 = ~n1193 & ~n1196;
  assign n1200 = a62 & b62;
  assign n1201 = ~a62 & ~b62;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1199 & n1202;
  assign n1204 = n1199 & ~n1202;
  assign s62 = ~n1203 & ~n1204;
  assign n1206 = ~n1200 & ~n1203;
  assign n1207 = a63 & b63;
  assign n1208 = ~a63 & ~b63;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n1206 & n1209;
  assign n1211 = n1206 & ~n1209;
  assign s63 = ~n1210 & ~n1211;
  assign n1213 = ~n1207 & ~n1210;
  assign n1214 = a64 & b64;
  assign n1215 = ~a64 & ~b64;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1213 & n1216;
  assign n1218 = n1213 & ~n1216;
  assign s64 = ~n1217 & ~n1218;
  assign n1220 = ~n1214 & ~n1217;
  assign n1221 = a65 & b65;
  assign n1222 = ~a65 & ~b65;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1220 & n1223;
  assign n1225 = n1220 & ~n1223;
  assign s65 = ~n1224 & ~n1225;
  assign n1227 = ~n1221 & ~n1224;
  assign n1228 = a66 & b66;
  assign n1229 = ~a66 & ~b66;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n1227 & n1230;
  assign n1232 = n1227 & ~n1230;
  assign s66 = ~n1231 & ~n1232;
  assign n1234 = ~n1228 & ~n1231;
  assign n1235 = a67 & b67;
  assign n1236 = ~a67 & ~b67;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~n1234 & n1237;
  assign n1239 = n1234 & ~n1237;
  assign s67 = ~n1238 & ~n1239;
  assign n1241 = ~n1235 & ~n1238;
  assign n1242 = a68 & b68;
  assign n1243 = ~a68 & ~b68;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1241 & n1244;
  assign n1246 = n1241 & ~n1244;
  assign s68 = ~n1245 & ~n1246;
  assign n1248 = ~n1242 & ~n1245;
  assign n1249 = a69 & b69;
  assign n1250 = ~a69 & ~b69;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1248 & n1251;
  assign n1253 = n1248 & ~n1251;
  assign s69 = ~n1252 & ~n1253;
  assign n1255 = ~n1249 & ~n1252;
  assign n1256 = a70 & b70;
  assign n1257 = ~a70 & ~b70;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n1255 & n1258;
  assign n1260 = n1255 & ~n1258;
  assign s70 = ~n1259 & ~n1260;
  assign n1262 = ~n1256 & ~n1259;
  assign n1263 = a71 & b71;
  assign n1264 = ~a71 & ~b71;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1262 & n1265;
  assign n1267 = n1262 & ~n1265;
  assign s71 = ~n1266 & ~n1267;
  assign n1269 = ~n1263 & ~n1266;
  assign n1270 = a72 & b72;
  assign n1271 = ~a72 & ~b72;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1269 & n1272;
  assign n1274 = n1269 & ~n1272;
  assign s72 = ~n1273 & ~n1274;
  assign n1276 = ~n1270 & ~n1273;
  assign n1277 = a73 & b73;
  assign n1278 = ~a73 & ~b73;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1276 & n1279;
  assign n1281 = n1276 & ~n1279;
  assign s73 = ~n1280 & ~n1281;
  assign n1283 = ~n1277 & ~n1280;
  assign n1284 = a74 & b74;
  assign n1285 = ~a74 & ~b74;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1283 & n1286;
  assign n1288 = n1283 & ~n1286;
  assign s74 = ~n1287 & ~n1288;
  assign n1290 = ~n1284 & ~n1287;
  assign n1291 = a75 & b75;
  assign n1292 = ~a75 & ~b75;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1290 & n1293;
  assign n1295 = n1290 & ~n1293;
  assign s75 = ~n1294 & ~n1295;
  assign n1297 = ~n1291 & ~n1294;
  assign n1298 = a76 & b76;
  assign n1299 = ~a76 & ~b76;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = ~n1297 & n1300;
  assign n1302 = n1297 & ~n1300;
  assign s76 = ~n1301 & ~n1302;
  assign n1304 = ~n1298 & ~n1301;
  assign n1305 = a77 & b77;
  assign n1306 = ~a77 & ~b77;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1304 & n1307;
  assign n1309 = n1304 & ~n1307;
  assign s77 = ~n1308 & ~n1309;
  assign n1311 = ~n1305 & ~n1308;
  assign n1312 = a78 & b78;
  assign n1313 = ~a78 & ~b78;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1311 & n1314;
  assign n1316 = n1311 & ~n1314;
  assign s78 = ~n1315 & ~n1316;
  assign n1318 = ~n1312 & ~n1315;
  assign n1319 = a79 & b79;
  assign n1320 = ~a79 & ~b79;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = ~n1318 & n1321;
  assign n1323 = n1318 & ~n1321;
  assign s79 = ~n1322 & ~n1323;
  assign n1325 = ~n1319 & ~n1322;
  assign n1326 = a80 & b80;
  assign n1327 = ~a80 & ~b80;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1325 & n1328;
  assign n1330 = n1325 & ~n1328;
  assign s80 = ~n1329 & ~n1330;
  assign n1332 = ~n1326 & ~n1329;
  assign n1333 = a81 & b81;
  assign n1334 = ~a81 & ~b81;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1332 & n1335;
  assign n1337 = n1332 & ~n1335;
  assign s81 = ~n1336 & ~n1337;
  assign n1339 = ~n1333 & ~n1336;
  assign n1340 = a82 & b82;
  assign n1341 = ~a82 & ~b82;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = ~n1339 & n1342;
  assign n1344 = n1339 & ~n1342;
  assign s82 = ~n1343 & ~n1344;
  assign n1346 = ~n1340 & ~n1343;
  assign n1347 = a83 & b83;
  assign n1348 = ~a83 & ~b83;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1346 & n1349;
  assign n1351 = n1346 & ~n1349;
  assign s83 = ~n1350 & ~n1351;
  assign n1353 = ~n1347 & ~n1350;
  assign n1354 = a84 & b84;
  assign n1355 = ~a84 & ~b84;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = ~n1353 & n1356;
  assign n1358 = n1353 & ~n1356;
  assign s84 = ~n1357 & ~n1358;
  assign n1360 = ~n1354 & ~n1357;
  assign n1361 = a85 & b85;
  assign n1362 = ~a85 & ~b85;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = ~n1360 & n1363;
  assign n1365 = n1360 & ~n1363;
  assign s85 = ~n1364 & ~n1365;
  assign n1367 = ~n1361 & ~n1364;
  assign n1368 = a86 & b86;
  assign n1369 = ~a86 & ~b86;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1367 & n1370;
  assign n1372 = n1367 & ~n1370;
  assign s86 = ~n1371 & ~n1372;
  assign n1374 = ~n1368 & ~n1371;
  assign n1375 = a87 & b87;
  assign n1376 = ~a87 & ~b87;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = ~n1374 & n1377;
  assign n1379 = n1374 & ~n1377;
  assign s87 = ~n1378 & ~n1379;
  assign n1381 = ~n1375 & ~n1378;
  assign n1382 = a88 & b88;
  assign n1383 = ~a88 & ~b88;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1381 & n1384;
  assign n1386 = n1381 & ~n1384;
  assign s88 = ~n1385 & ~n1386;
  assign n1388 = ~n1382 & ~n1385;
  assign n1389 = a89 & b89;
  assign n1390 = ~a89 & ~b89;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1388 & n1391;
  assign n1393 = n1388 & ~n1391;
  assign s89 = ~n1392 & ~n1393;
  assign n1395 = ~n1389 & ~n1392;
  assign n1396 = a90 & b90;
  assign n1397 = ~a90 & ~b90;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1395 & n1398;
  assign n1400 = n1395 & ~n1398;
  assign s90 = ~n1399 & ~n1400;
  assign n1402 = ~n1396 & ~n1399;
  assign n1403 = a91 & b91;
  assign n1404 = ~a91 & ~b91;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1402 & n1405;
  assign n1407 = n1402 & ~n1405;
  assign s91 = ~n1406 & ~n1407;
  assign n1409 = ~n1403 & ~n1406;
  assign n1410 = a92 & b92;
  assign n1411 = ~a92 & ~b92;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~n1409 & n1412;
  assign n1414 = n1409 & ~n1412;
  assign s92 = ~n1413 & ~n1414;
  assign n1416 = ~n1410 & ~n1413;
  assign n1417 = a93 & b93;
  assign n1418 = ~a93 & ~b93;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~n1416 & n1419;
  assign n1421 = n1416 & ~n1419;
  assign s93 = ~n1420 & ~n1421;
  assign n1423 = ~n1417 & ~n1420;
  assign n1424 = a94 & b94;
  assign n1425 = ~a94 & ~b94;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n1423 & n1426;
  assign n1428 = n1423 & ~n1426;
  assign s94 = ~n1427 & ~n1428;
  assign n1430 = ~n1424 & ~n1427;
  assign n1431 = a95 & b95;
  assign n1432 = ~a95 & ~b95;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = n1430 & ~n1433;
  assign s95 = ~n1434 & ~n1435;
  assign n1437 = ~n1431 & ~n1434;
  assign n1438 = a96 & b96;
  assign n1439 = ~a96 & ~b96;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1437 & n1440;
  assign n1442 = n1437 & ~n1440;
  assign s96 = ~n1441 & ~n1442;
  assign n1444 = ~n1438 & ~n1441;
  assign n1445 = a97 & b97;
  assign n1446 = ~a97 & ~b97;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1444 & n1447;
  assign n1449 = n1444 & ~n1447;
  assign s97 = ~n1448 & ~n1449;
  assign n1451 = ~n1445 & ~n1448;
  assign n1452 = a98 & b98;
  assign n1453 = ~a98 & ~b98;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1451 & n1454;
  assign n1456 = n1451 & ~n1454;
  assign s98 = ~n1455 & ~n1456;
  assign n1458 = ~n1452 & ~n1455;
  assign n1459 = a99 & b99;
  assign n1460 = ~a99 & ~b99;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1458 & n1461;
  assign n1463 = n1458 & ~n1461;
  assign s99 = ~n1462 & ~n1463;
  assign n1465 = ~n1459 & ~n1462;
  assign n1466 = a100 & b100;
  assign n1467 = ~a100 & ~b100;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = ~n1465 & n1468;
  assign n1470 = n1465 & ~n1468;
  assign s100 = ~n1469 & ~n1470;
  assign n1472 = ~n1466 & ~n1469;
  assign n1473 = a101 & b101;
  assign n1474 = ~a101 & ~b101;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n1472 & n1475;
  assign n1477 = n1472 & ~n1475;
  assign s101 = ~n1476 & ~n1477;
  assign n1479 = ~n1473 & ~n1476;
  assign n1480 = a102 & b102;
  assign n1481 = ~a102 & ~b102;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1479 & n1482;
  assign n1484 = n1479 & ~n1482;
  assign s102 = ~n1483 & ~n1484;
  assign n1486 = ~n1480 & ~n1483;
  assign n1487 = a103 & b103;
  assign n1488 = ~a103 & ~b103;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1486 & n1489;
  assign n1491 = n1486 & ~n1489;
  assign s103 = ~n1490 & ~n1491;
  assign n1493 = ~n1487 & ~n1490;
  assign n1494 = a104 & b104;
  assign n1495 = ~a104 & ~b104;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1493 & n1496;
  assign n1498 = n1493 & ~n1496;
  assign s104 = ~n1497 & ~n1498;
  assign n1500 = ~n1494 & ~n1497;
  assign n1501 = a105 & b105;
  assign n1502 = ~a105 & ~b105;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~n1500 & n1503;
  assign n1505 = n1500 & ~n1503;
  assign s105 = ~n1504 & ~n1505;
  assign n1507 = ~n1501 & ~n1504;
  assign n1508 = a106 & b106;
  assign n1509 = ~a106 & ~b106;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1507 & n1510;
  assign n1512 = n1507 & ~n1510;
  assign s106 = ~n1511 & ~n1512;
  assign n1514 = ~n1508 & ~n1511;
  assign n1515 = a107 & b107;
  assign n1516 = ~a107 & ~b107;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1514 & n1517;
  assign n1519 = n1514 & ~n1517;
  assign s107 = ~n1518 & ~n1519;
  assign n1521 = ~n1515 & ~n1518;
  assign n1522 = a108 & b108;
  assign n1523 = ~a108 & ~b108;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1521 & n1524;
  assign n1526 = n1521 & ~n1524;
  assign s108 = ~n1525 & ~n1526;
  assign n1528 = ~n1522 & ~n1525;
  assign n1529 = a109 & b109;
  assign n1530 = ~a109 & ~b109;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n1528 & n1531;
  assign n1533 = n1528 & ~n1531;
  assign s109 = ~n1532 & ~n1533;
  assign n1535 = ~n1529 & ~n1532;
  assign n1536 = a110 & b110;
  assign n1537 = ~a110 & ~b110;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1535 & n1538;
  assign n1540 = n1535 & ~n1538;
  assign s110 = ~n1539 & ~n1540;
  assign n1542 = ~n1536 & ~n1539;
  assign n1543 = a111 & b111;
  assign n1544 = ~a111 & ~b111;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~n1542 & n1545;
  assign n1547 = n1542 & ~n1545;
  assign s111 = ~n1546 & ~n1547;
  assign n1549 = ~n1543 & ~n1546;
  assign n1550 = a112 & b112;
  assign n1551 = ~a112 & ~b112;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1549 & n1552;
  assign n1554 = n1549 & ~n1552;
  assign s112 = ~n1553 & ~n1554;
  assign n1556 = ~n1550 & ~n1553;
  assign n1557 = a113 & b113;
  assign n1558 = ~a113 & ~b113;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1556 & n1559;
  assign n1561 = n1556 & ~n1559;
  assign s113 = ~n1560 & ~n1561;
  assign n1563 = ~n1557 & ~n1560;
  assign n1564 = a114 & b114;
  assign n1565 = ~a114 & ~b114;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = ~n1563 & n1566;
  assign n1568 = n1563 & ~n1566;
  assign s114 = ~n1567 & ~n1568;
  assign n1570 = ~n1564 & ~n1567;
  assign n1571 = a115 & b115;
  assign n1572 = ~a115 & ~b115;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1570 & n1573;
  assign n1575 = n1570 & ~n1573;
  assign s115 = ~n1574 & ~n1575;
  assign n1577 = ~n1571 & ~n1574;
  assign n1578 = a116 & b116;
  assign n1579 = ~a116 & ~b116;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1577 & n1580;
  assign n1582 = n1577 & ~n1580;
  assign s116 = ~n1581 & ~n1582;
  assign n1584 = ~n1578 & ~n1581;
  assign n1585 = a117 & b117;
  assign n1586 = ~a117 & ~b117;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = ~n1584 & n1587;
  assign n1589 = n1584 & ~n1587;
  assign s117 = ~n1588 & ~n1589;
  assign n1591 = ~n1585 & ~n1588;
  assign n1592 = a118 & b118;
  assign n1593 = ~a118 & ~b118;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1591 & n1594;
  assign n1596 = n1591 & ~n1594;
  assign s118 = ~n1595 & ~n1596;
  assign n1598 = ~n1592 & ~n1595;
  assign n1599 = a119 & b119;
  assign n1600 = ~a119 & ~b119;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = ~n1598 & n1601;
  assign n1603 = n1598 & ~n1601;
  assign s119 = ~n1602 & ~n1603;
  assign n1605 = ~n1599 & ~n1602;
  assign n1606 = a120 & b120;
  assign n1607 = ~a120 & ~b120;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = ~n1605 & n1608;
  assign n1610 = n1605 & ~n1608;
  assign s120 = ~n1609 & ~n1610;
  assign n1612 = ~n1606 & ~n1609;
  assign n1613 = a121 & b121;
  assign n1614 = ~a121 & ~b121;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = n1612 & ~n1615;
  assign s121 = ~n1616 & ~n1617;
  assign n1619 = ~n1613 & ~n1616;
  assign n1620 = a122 & b122;
  assign n1621 = ~a122 & ~b122;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = ~n1619 & n1622;
  assign n1624 = n1619 & ~n1622;
  assign s122 = ~n1623 & ~n1624;
  assign n1626 = ~n1620 & ~n1623;
  assign n1627 = a123 & b123;
  assign n1628 = ~a123 & ~b123;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~n1626 & n1629;
  assign n1631 = n1626 & ~n1629;
  assign s123 = ~n1630 & ~n1631;
  assign n1633 = ~n1627 & ~n1630;
  assign n1634 = a124 & b124;
  assign n1635 = ~a124 & ~b124;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1633 & n1636;
  assign n1638 = n1633 & ~n1636;
  assign s124 = ~n1637 & ~n1638;
  assign n1640 = ~n1634 & ~n1637;
  assign n1641 = a125 & b125;
  assign n1642 = ~a125 & ~b125;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1640 & n1643;
  assign n1645 = n1640 & ~n1643;
  assign s125 = ~n1644 & ~n1645;
  assign n1647 = ~n1641 & ~n1644;
  assign n1648 = a126 & b126;
  assign n1649 = ~a126 & ~b126;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~n1647 & n1650;
  assign n1652 = n1647 & ~n1650;
  assign s126 = ~n1651 & ~n1652;
  assign n1654 = ~n1648 & ~n1651;
  assign n1655 = a127 & b127;
  assign n1656 = ~a127 & ~b127;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = ~n1654 & n1657;
  assign n1659 = n1654 & ~n1657;
  assign s127 = ~n1658 & ~n1659;
  assign n1661 = ~n1655 & ~n1658;
  assign n1662 = a128 & b128;
  assign n1663 = ~a128 & ~b128;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1661 & n1664;
  assign n1666 = n1661 & ~n1664;
  assign s128 = ~n1665 & ~n1666;
  assign n1668 = ~n1662 & ~n1665;
  assign n1669 = a129 & b129;
  assign n1670 = ~a129 & ~b129;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1668 & n1671;
  assign n1673 = n1668 & ~n1671;
  assign s129 = ~n1672 & ~n1673;
  assign n1675 = ~n1669 & ~n1672;
  assign n1676 = a130 & b130;
  assign n1677 = ~a130 & ~b130;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1675 & n1678;
  assign n1680 = n1675 & ~n1678;
  assign s130 = ~n1679 & ~n1680;
  assign n1682 = ~n1676 & ~n1679;
  assign n1683 = a131 & b131;
  assign n1684 = ~a131 & ~b131;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1682 & n1685;
  assign n1687 = n1682 & ~n1685;
  assign s131 = ~n1686 & ~n1687;
  assign n1689 = ~n1683 & ~n1686;
  assign n1690 = a132 & b132;
  assign n1691 = ~a132 & ~b132;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1689 & n1692;
  assign n1694 = n1689 & ~n1692;
  assign s132 = ~n1693 & ~n1694;
  assign n1696 = ~n1690 & ~n1693;
  assign n1697 = a133 & b133;
  assign n1698 = ~a133 & ~b133;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1696 & n1699;
  assign n1701 = n1696 & ~n1699;
  assign s133 = ~n1700 & ~n1701;
  assign n1703 = ~n1697 & ~n1700;
  assign n1704 = a134 & b134;
  assign n1705 = ~a134 & ~b134;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1703 & n1706;
  assign n1708 = n1703 & ~n1706;
  assign s134 = ~n1707 & ~n1708;
  assign n1710 = ~n1704 & ~n1707;
  assign n1711 = a135 & b135;
  assign n1712 = ~a135 & ~b135;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = ~n1710 & n1713;
  assign n1715 = n1710 & ~n1713;
  assign s135 = ~n1714 & ~n1715;
  assign n1717 = ~n1711 & ~n1714;
  assign n1718 = a136 & b136;
  assign n1719 = ~a136 & ~b136;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~n1717 & n1720;
  assign n1722 = n1717 & ~n1720;
  assign s136 = ~n1721 & ~n1722;
  assign n1724 = ~n1718 & ~n1721;
  assign n1725 = a137 & b137;
  assign n1726 = ~a137 & ~b137;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1724 & n1727;
  assign n1729 = n1724 & ~n1727;
  assign s137 = ~n1728 & ~n1729;
  assign n1731 = ~n1725 & ~n1728;
  assign n1732 = a138 & b138;
  assign n1733 = ~a138 & ~b138;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~n1731 & n1734;
  assign n1736 = n1731 & ~n1734;
  assign s138 = ~n1735 & ~n1736;
  assign n1738 = ~n1732 & ~n1735;
  assign n1739 = a139 & b139;
  assign n1740 = ~a139 & ~b139;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1738 & n1741;
  assign n1743 = n1738 & ~n1741;
  assign s139 = ~n1742 & ~n1743;
  assign n1745 = ~n1739 & ~n1742;
  assign n1746 = a140 & b140;
  assign n1747 = ~a140 & ~b140;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = ~n1745 & n1748;
  assign n1750 = n1745 & ~n1748;
  assign s140 = ~n1749 & ~n1750;
  assign n1752 = ~n1746 & ~n1749;
  assign n1753 = a141 & b141;
  assign n1754 = ~a141 & ~b141;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n1752 & n1755;
  assign n1757 = n1752 & ~n1755;
  assign s141 = ~n1756 & ~n1757;
  assign n1759 = ~n1753 & ~n1756;
  assign n1760 = a142 & b142;
  assign n1761 = ~a142 & ~b142;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1759 & n1762;
  assign n1764 = n1759 & ~n1762;
  assign s142 = ~n1763 & ~n1764;
  assign n1766 = ~n1760 & ~n1763;
  assign n1767 = a143 & b143;
  assign n1768 = ~a143 & ~b143;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = ~n1766 & n1769;
  assign n1771 = n1766 & ~n1769;
  assign s143 = ~n1770 & ~n1771;
  assign n1773 = ~n1767 & ~n1770;
  assign n1774 = a144 & b144;
  assign n1775 = ~a144 & ~b144;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = ~n1773 & n1776;
  assign n1778 = n1773 & ~n1776;
  assign s144 = ~n1777 & ~n1778;
  assign n1780 = ~n1774 & ~n1777;
  assign n1781 = a145 & b145;
  assign n1782 = ~a145 & ~b145;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1780 & n1783;
  assign n1785 = n1780 & ~n1783;
  assign s145 = ~n1784 & ~n1785;
  assign n1787 = ~n1781 & ~n1784;
  assign n1788 = a146 & b146;
  assign n1789 = ~a146 & ~b146;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1787 & n1790;
  assign n1792 = n1787 & ~n1790;
  assign s146 = ~n1791 & ~n1792;
  assign n1794 = ~n1788 & ~n1791;
  assign n1795 = a147 & b147;
  assign n1796 = ~a147 & ~b147;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n1794 & n1797;
  assign n1799 = n1794 & ~n1797;
  assign s147 = ~n1798 & ~n1799;
  assign n1801 = ~n1795 & ~n1798;
  assign n1802 = a148 & b148;
  assign n1803 = ~a148 & ~b148;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1801 & n1804;
  assign n1806 = n1801 & ~n1804;
  assign s148 = ~n1805 & ~n1806;
  assign n1808 = ~n1802 & ~n1805;
  assign n1809 = a149 & b149;
  assign n1810 = ~a149 & ~b149;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n1808 & n1811;
  assign n1813 = n1808 & ~n1811;
  assign s149 = ~n1812 & ~n1813;
  assign n1815 = ~n1809 & ~n1812;
  assign n1816 = a150 & b150;
  assign n1817 = ~a150 & ~b150;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1815 & n1818;
  assign n1820 = n1815 & ~n1818;
  assign s150 = ~n1819 & ~n1820;
  assign n1822 = ~n1816 & ~n1819;
  assign n1823 = a151 & b151;
  assign n1824 = ~a151 & ~b151;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = ~n1822 & n1825;
  assign n1827 = n1822 & ~n1825;
  assign s151 = ~n1826 & ~n1827;
  assign n1829 = ~n1823 & ~n1826;
  assign n1830 = a152 & b152;
  assign n1831 = ~a152 & ~b152;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1829 & n1832;
  assign n1834 = n1829 & ~n1832;
  assign s152 = ~n1833 & ~n1834;
  assign n1836 = ~n1830 & ~n1833;
  assign n1837 = a153 & b153;
  assign n1838 = ~a153 & ~b153;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~n1836 & n1839;
  assign n1841 = n1836 & ~n1839;
  assign s153 = ~n1840 & ~n1841;
  assign n1843 = ~n1837 & ~n1840;
  assign n1844 = a154 & b154;
  assign n1845 = ~a154 & ~b154;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = ~n1843 & n1846;
  assign n1848 = n1843 & ~n1846;
  assign s154 = ~n1847 & ~n1848;
  assign n1850 = ~n1844 & ~n1847;
  assign n1851 = a155 & b155;
  assign n1852 = ~a155 & ~b155;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = ~n1850 & n1853;
  assign n1855 = n1850 & ~n1853;
  assign s155 = ~n1854 & ~n1855;
  assign n1857 = ~n1851 & ~n1854;
  assign n1858 = a156 & b156;
  assign n1859 = ~a156 & ~b156;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & n1860;
  assign n1862 = n1857 & ~n1860;
  assign s156 = ~n1861 & ~n1862;
  assign n1864 = ~n1858 & ~n1861;
  assign n1865 = a157 & b157;
  assign n1866 = ~a157 & ~b157;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = ~n1864 & n1867;
  assign n1869 = n1864 & ~n1867;
  assign s157 = ~n1868 & ~n1869;
  assign n1871 = ~n1865 & ~n1868;
  assign n1872 = a158 & b158;
  assign n1873 = ~a158 & ~b158;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1871 & n1874;
  assign n1876 = n1871 & ~n1874;
  assign s158 = ~n1875 & ~n1876;
  assign n1878 = ~n1872 & ~n1875;
  assign n1879 = a159 & b159;
  assign n1880 = ~a159 & ~b159;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~n1878 & n1881;
  assign n1883 = n1878 & ~n1881;
  assign s159 = ~n1882 & ~n1883;
  assign n1885 = ~n1879 & ~n1882;
  assign n1886 = a160 & b160;
  assign n1887 = ~a160 & ~b160;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = ~n1885 & n1888;
  assign n1890 = n1885 & ~n1888;
  assign s160 = ~n1889 & ~n1890;
  assign n1892 = ~n1886 & ~n1889;
  assign n1893 = a161 & b161;
  assign n1894 = ~a161 & ~b161;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = ~n1892 & n1895;
  assign n1897 = n1892 & ~n1895;
  assign s161 = ~n1896 & ~n1897;
  assign n1899 = ~n1893 & ~n1896;
  assign n1900 = a162 & b162;
  assign n1901 = ~a162 & ~b162;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = ~n1899 & n1902;
  assign n1904 = n1899 & ~n1902;
  assign s162 = ~n1903 & ~n1904;
  assign n1906 = ~n1900 & ~n1903;
  assign n1907 = a163 & b163;
  assign n1908 = ~a163 & ~b163;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = ~n1906 & n1909;
  assign n1911 = n1906 & ~n1909;
  assign s163 = ~n1910 & ~n1911;
  assign n1913 = ~n1907 & ~n1910;
  assign n1914 = a164 & b164;
  assign n1915 = ~a164 & ~b164;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1913 & n1916;
  assign n1918 = n1913 & ~n1916;
  assign s164 = ~n1917 & ~n1918;
  assign n1920 = ~n1914 & ~n1917;
  assign n1921 = a165 & b165;
  assign n1922 = ~a165 & ~b165;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~n1920 & n1923;
  assign n1925 = n1920 & ~n1923;
  assign s165 = ~n1924 & ~n1925;
  assign n1927 = ~n1921 & ~n1924;
  assign n1928 = a166 & b166;
  assign n1929 = ~a166 & ~b166;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = ~n1927 & n1930;
  assign n1932 = n1927 & ~n1930;
  assign s166 = ~n1931 & ~n1932;
  assign n1934 = ~n1928 & ~n1931;
  assign n1935 = a167 & b167;
  assign n1936 = ~a167 & ~b167;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = ~n1934 & n1937;
  assign n1939 = n1934 & ~n1937;
  assign s167 = ~n1938 & ~n1939;
  assign n1941 = ~n1935 & ~n1938;
  assign n1942 = a168 & b168;
  assign n1943 = ~a168 & ~b168;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1941 & n1944;
  assign n1946 = n1941 & ~n1944;
  assign s168 = ~n1945 & ~n1946;
  assign n1948 = ~n1942 & ~n1945;
  assign n1949 = a169 & b169;
  assign n1950 = ~a169 & ~b169;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n1948 & n1951;
  assign n1953 = n1948 & ~n1951;
  assign s169 = ~n1952 & ~n1953;
  assign n1955 = ~n1949 & ~n1952;
  assign n1956 = a170 & b170;
  assign n1957 = ~a170 & ~b170;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = ~n1955 & n1958;
  assign n1960 = n1955 & ~n1958;
  assign s170 = ~n1959 & ~n1960;
  assign n1962 = ~n1956 & ~n1959;
  assign n1963 = a171 & b171;
  assign n1964 = ~a171 & ~b171;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n1962 & n1965;
  assign n1967 = n1962 & ~n1965;
  assign s171 = ~n1966 & ~n1967;
  assign n1969 = ~n1963 & ~n1966;
  assign n1970 = a172 & b172;
  assign n1971 = ~a172 & ~b172;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & n1972;
  assign n1974 = n1969 & ~n1972;
  assign s172 = ~n1973 & ~n1974;
  assign n1976 = ~n1970 & ~n1973;
  assign n1977 = a173 & b173;
  assign n1978 = ~a173 & ~b173;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~n1976 & n1979;
  assign n1981 = n1976 & ~n1979;
  assign s173 = ~n1980 & ~n1981;
  assign n1983 = ~n1977 & ~n1980;
  assign n1984 = a174 & b174;
  assign n1985 = ~a174 & ~b174;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n1983 & n1986;
  assign n1988 = n1983 & ~n1986;
  assign s174 = ~n1987 & ~n1988;
  assign n1990 = ~n1984 & ~n1987;
  assign n1991 = a175 & b175;
  assign n1992 = ~a175 & ~b175;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n1990 & n1993;
  assign n1995 = n1990 & ~n1993;
  assign s175 = ~n1994 & ~n1995;
  assign n1997 = ~n1991 & ~n1994;
  assign n1998 = a176 & b176;
  assign n1999 = ~a176 & ~b176;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~n1997 & n2000;
  assign n2002 = n1997 & ~n2000;
  assign s176 = ~n2001 & ~n2002;
  assign n2004 = ~n1998 & ~n2001;
  assign n2005 = a177 & b177;
  assign n2006 = ~a177 & ~b177;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = ~n2004 & n2007;
  assign n2009 = n2004 & ~n2007;
  assign s177 = ~n2008 & ~n2009;
  assign n2011 = ~n2005 & ~n2008;
  assign n2012 = a178 & b178;
  assign n2013 = ~a178 & ~b178;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n2011 & n2014;
  assign n2016 = n2011 & ~n2014;
  assign s178 = ~n2015 & ~n2016;
  assign n2018 = ~n2012 & ~n2015;
  assign n2019 = a179 & b179;
  assign n2020 = ~a179 & ~b179;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = ~n2018 & n2021;
  assign n2023 = n2018 & ~n2021;
  assign s179 = ~n2022 & ~n2023;
  assign n2025 = ~n2019 & ~n2022;
  assign n2026 = a180 & b180;
  assign n2027 = ~a180 & ~b180;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = ~n2025 & n2028;
  assign n2030 = n2025 & ~n2028;
  assign s180 = ~n2029 & ~n2030;
  assign n2032 = ~n2026 & ~n2029;
  assign n2033 = a181 & b181;
  assign n2034 = ~a181 & ~b181;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = ~n2032 & n2035;
  assign n2037 = n2032 & ~n2035;
  assign s181 = ~n2036 & ~n2037;
  assign n2039 = ~n2033 & ~n2036;
  assign n2040 = a182 & b182;
  assign n2041 = ~a182 & ~b182;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = ~n2039 & n2042;
  assign n2044 = n2039 & ~n2042;
  assign s182 = ~n2043 & ~n2044;
  assign n2046 = ~n2040 & ~n2043;
  assign n2047 = a183 & b183;
  assign n2048 = ~a183 & ~b183;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = ~n2046 & n2049;
  assign n2051 = n2046 & ~n2049;
  assign s183 = ~n2050 & ~n2051;
  assign n2053 = ~n2047 & ~n2050;
  assign n2054 = a184 & b184;
  assign n2055 = ~a184 & ~b184;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~n2053 & n2056;
  assign n2058 = n2053 & ~n2056;
  assign s184 = ~n2057 & ~n2058;
  assign n2060 = ~n2054 & ~n2057;
  assign n2061 = a185 & b185;
  assign n2062 = ~a185 & ~b185;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2060 & n2063;
  assign n2065 = n2060 & ~n2063;
  assign s185 = ~n2064 & ~n2065;
  assign n2067 = ~n2061 & ~n2064;
  assign n2068 = a186 & b186;
  assign n2069 = ~a186 & ~b186;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2067 & n2070;
  assign n2072 = n2067 & ~n2070;
  assign s186 = ~n2071 & ~n2072;
  assign n2074 = ~n2068 & ~n2071;
  assign n2075 = a187 & b187;
  assign n2076 = ~a187 & ~b187;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = ~n2074 & n2077;
  assign n2079 = n2074 & ~n2077;
  assign s187 = ~n2078 & ~n2079;
  assign n2081 = ~n2075 & ~n2078;
  assign n2082 = a188 & b188;
  assign n2083 = ~a188 & ~b188;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = ~n2081 & n2084;
  assign n2086 = n2081 & ~n2084;
  assign s188 = ~n2085 & ~n2086;
  assign n2088 = ~n2082 & ~n2085;
  assign n2089 = a189 & b189;
  assign n2090 = ~a189 & ~b189;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = n2088 & ~n2091;
  assign s189 = ~n2092 & ~n2093;
  assign n2095 = ~n2089 & ~n2092;
  assign n2096 = a190 & b190;
  assign n2097 = ~a190 & ~b190;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2095 & n2098;
  assign n2100 = n2095 & ~n2098;
  assign s190 = ~n2099 & ~n2100;
  assign n2102 = ~n2096 & ~n2099;
  assign n2103 = a191 & b191;
  assign n2104 = ~a191 & ~b191;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = ~n2102 & n2105;
  assign n2107 = n2102 & ~n2105;
  assign s191 = ~n2106 & ~n2107;
  assign n2109 = ~n2103 & ~n2106;
  assign n2110 = a192 & b192;
  assign n2111 = ~a192 & ~b192;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~n2109 & n2112;
  assign n2114 = n2109 & ~n2112;
  assign s192 = ~n2113 & ~n2114;
  assign n2116 = ~n2110 & ~n2113;
  assign n2117 = a193 & b193;
  assign n2118 = ~a193 & ~b193;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~n2116 & n2119;
  assign n2121 = n2116 & ~n2119;
  assign s193 = ~n2120 & ~n2121;
  assign n2123 = ~n2117 & ~n2120;
  assign n2124 = a194 & b194;
  assign n2125 = ~a194 & ~b194;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2123 & n2126;
  assign n2128 = n2123 & ~n2126;
  assign s194 = ~n2127 & ~n2128;
  assign n2130 = ~n2124 & ~n2127;
  assign n2131 = a195 & b195;
  assign n2132 = ~a195 & ~b195;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = ~n2130 & n2133;
  assign n2135 = n2130 & ~n2133;
  assign s195 = ~n2134 & ~n2135;
  assign n2137 = ~n2131 & ~n2134;
  assign n2138 = a196 & b196;
  assign n2139 = ~a196 & ~b196;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = ~n2137 & n2140;
  assign n2142 = n2137 & ~n2140;
  assign s196 = ~n2141 & ~n2142;
  assign n2144 = ~n2138 & ~n2141;
  assign n2145 = a197 & b197;
  assign n2146 = ~a197 & ~b197;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2144 & n2147;
  assign n2149 = n2144 & ~n2147;
  assign s197 = ~n2148 & ~n2149;
  assign n2151 = ~n2145 & ~n2148;
  assign n2152 = a198 & b198;
  assign n2153 = ~a198 & ~b198;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = ~n2151 & n2154;
  assign n2156 = n2151 & ~n2154;
  assign s198 = ~n2155 & ~n2156;
  assign n2158 = ~n2152 & ~n2155;
  assign n2159 = a199 & b199;
  assign n2160 = ~a199 & ~b199;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n2158 & n2161;
  assign n2163 = n2158 & ~n2161;
  assign s199 = ~n2162 & ~n2163;
  assign n2165 = ~n2159 & ~n2162;
  assign n2166 = a200 & b200;
  assign n2167 = ~a200 & ~b200;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~n2165 & n2168;
  assign n2170 = n2165 & ~n2168;
  assign s200 = ~n2169 & ~n2170;
  assign n2172 = ~n2166 & ~n2169;
  assign n2173 = a201 & b201;
  assign n2174 = ~a201 & ~b201;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = ~n2172 & n2175;
  assign n2177 = n2172 & ~n2175;
  assign s201 = ~n2176 & ~n2177;
  assign n2179 = ~n2173 & ~n2176;
  assign n2180 = a202 & b202;
  assign n2181 = ~a202 & ~b202;
  assign n2182 = ~n2180 & ~n2181;
  assign n2183 = ~n2179 & n2182;
  assign n2184 = n2179 & ~n2182;
  assign s202 = ~n2183 & ~n2184;
  assign n2186 = ~n2180 & ~n2183;
  assign n2187 = a203 & b203;
  assign n2188 = ~a203 & ~b203;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = ~n2186 & n2189;
  assign n2191 = n2186 & ~n2189;
  assign s203 = ~n2190 & ~n2191;
  assign n2193 = ~n2187 & ~n2190;
  assign n2194 = a204 & b204;
  assign n2195 = ~a204 & ~b204;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = ~n2193 & n2196;
  assign n2198 = n2193 & ~n2196;
  assign s204 = ~n2197 & ~n2198;
  assign n2200 = ~n2194 & ~n2197;
  assign n2201 = a205 & b205;
  assign n2202 = ~a205 & ~b205;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = ~n2200 & n2203;
  assign n2205 = n2200 & ~n2203;
  assign s205 = ~n2204 & ~n2205;
  assign n2207 = ~n2201 & ~n2204;
  assign n2208 = a206 & b206;
  assign n2209 = ~a206 & ~b206;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = ~n2207 & n2210;
  assign n2212 = n2207 & ~n2210;
  assign s206 = ~n2211 & ~n2212;
  assign n2214 = ~n2208 & ~n2211;
  assign n2215 = a207 & b207;
  assign n2216 = ~a207 & ~b207;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2214 & n2217;
  assign n2219 = n2214 & ~n2217;
  assign s207 = ~n2218 & ~n2219;
  assign n2221 = ~n2215 & ~n2218;
  assign n2222 = a208 & b208;
  assign n2223 = ~a208 & ~b208;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~n2221 & n2224;
  assign n2226 = n2221 & ~n2224;
  assign s208 = ~n2225 & ~n2226;
  assign n2228 = ~n2222 & ~n2225;
  assign n2229 = a209 & b209;
  assign n2230 = ~a209 & ~b209;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = ~n2228 & n2231;
  assign n2233 = n2228 & ~n2231;
  assign s209 = ~n2232 & ~n2233;
  assign n2235 = ~n2229 & ~n2232;
  assign n2236 = a210 & b210;
  assign n2237 = ~a210 & ~b210;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n2235 & n2238;
  assign n2240 = n2235 & ~n2238;
  assign s210 = ~n2239 & ~n2240;
  assign n2242 = ~n2236 & ~n2239;
  assign n2243 = a211 & b211;
  assign n2244 = ~a211 & ~b211;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = ~n2242 & n2245;
  assign n2247 = n2242 & ~n2245;
  assign s211 = ~n2246 & ~n2247;
  assign n2249 = ~n2243 & ~n2246;
  assign n2250 = a212 & b212;
  assign n2251 = ~a212 & ~b212;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = ~n2249 & n2252;
  assign n2254 = n2249 & ~n2252;
  assign s212 = ~n2253 & ~n2254;
  assign n2256 = ~n2250 & ~n2253;
  assign n2257 = a213 & b213;
  assign n2258 = ~a213 & ~b213;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2256 & n2259;
  assign n2261 = n2256 & ~n2259;
  assign s213 = ~n2260 & ~n2261;
  assign n2263 = ~n2257 & ~n2260;
  assign n2264 = a214 & b214;
  assign n2265 = ~a214 & ~b214;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n2263 & n2266;
  assign n2268 = n2263 & ~n2266;
  assign s214 = ~n2267 & ~n2268;
  assign n2270 = ~n2264 & ~n2267;
  assign n2271 = a215 & b215;
  assign n2272 = ~a215 & ~b215;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2270 & n2273;
  assign n2275 = n2270 & ~n2273;
  assign s215 = ~n2274 & ~n2275;
  assign n2277 = ~n2271 & ~n2274;
  assign n2278 = a216 & b216;
  assign n2279 = ~a216 & ~b216;
  assign n2280 = ~n2278 & ~n2279;
  assign n2281 = ~n2277 & n2280;
  assign n2282 = n2277 & ~n2280;
  assign s216 = ~n2281 & ~n2282;
  assign n2284 = ~n2278 & ~n2281;
  assign n2285 = a217 & b217;
  assign n2286 = ~a217 & ~b217;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = ~n2284 & n2287;
  assign n2289 = n2284 & ~n2287;
  assign s217 = ~n2288 & ~n2289;
  assign n2291 = ~n2285 & ~n2288;
  assign n2292 = a218 & b218;
  assign n2293 = ~a218 & ~b218;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n2291 & n2294;
  assign n2296 = n2291 & ~n2294;
  assign s218 = ~n2295 & ~n2296;
  assign n2298 = ~n2292 & ~n2295;
  assign n2299 = a219 & b219;
  assign n2300 = ~a219 & ~b219;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = n2298 & ~n2301;
  assign s219 = ~n2302 & ~n2303;
  assign n2305 = ~n2299 & ~n2302;
  assign n2306 = a220 & b220;
  assign n2307 = ~a220 & ~b220;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n2305 & n2308;
  assign n2310 = n2305 & ~n2308;
  assign s220 = ~n2309 & ~n2310;
  assign n2312 = ~n2306 & ~n2309;
  assign n2313 = a221 & b221;
  assign n2314 = ~a221 & ~b221;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n2312 & n2315;
  assign n2317 = n2312 & ~n2315;
  assign s221 = ~n2316 & ~n2317;
  assign n2319 = ~n2313 & ~n2316;
  assign n2320 = a222 & b222;
  assign n2321 = ~a222 & ~b222;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = ~n2319 & n2322;
  assign n2324 = n2319 & ~n2322;
  assign s222 = ~n2323 & ~n2324;
  assign n2326 = ~n2320 & ~n2323;
  assign n2327 = a223 & b223;
  assign n2328 = ~a223 & ~b223;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = ~n2326 & n2329;
  assign n2331 = n2326 & ~n2329;
  assign s223 = ~n2330 & ~n2331;
  assign n2333 = ~n2327 & ~n2330;
  assign n2334 = a224 & b224;
  assign n2335 = ~a224 & ~b224;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = ~n2333 & n2336;
  assign n2338 = n2333 & ~n2336;
  assign s224 = ~n2337 & ~n2338;
  assign n2340 = ~n2334 & ~n2337;
  assign n2341 = a225 & b225;
  assign n2342 = ~a225 & ~b225;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = ~n2340 & n2343;
  assign n2345 = n2340 & ~n2343;
  assign s225 = ~n2344 & ~n2345;
  assign n2347 = ~n2341 & ~n2344;
  assign n2348 = a226 & b226;
  assign n2349 = ~a226 & ~b226;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~n2347 & n2350;
  assign n2352 = n2347 & ~n2350;
  assign s226 = ~n2351 & ~n2352;
  assign n2354 = ~n2348 & ~n2351;
  assign n2355 = a227 & b227;
  assign n2356 = ~a227 & ~b227;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = ~n2354 & n2357;
  assign n2359 = n2354 & ~n2357;
  assign s227 = ~n2358 & ~n2359;
  assign n2361 = ~n2355 & ~n2358;
  assign n2362 = a228 & b228;
  assign n2363 = ~a228 & ~b228;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = ~n2361 & n2364;
  assign n2366 = n2361 & ~n2364;
  assign s228 = ~n2365 & ~n2366;
  assign n2368 = ~n2362 & ~n2365;
  assign n2369 = a229 & b229;
  assign n2370 = ~a229 & ~b229;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n2368 & n2371;
  assign n2373 = n2368 & ~n2371;
  assign s229 = ~n2372 & ~n2373;
  assign n2375 = ~n2369 & ~n2372;
  assign n2376 = a230 & b230;
  assign n2377 = ~a230 & ~b230;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = ~n2375 & n2378;
  assign n2380 = n2375 & ~n2378;
  assign s230 = ~n2379 & ~n2380;
  assign n2382 = ~n2376 & ~n2379;
  assign n2383 = a231 & b231;
  assign n2384 = ~a231 & ~b231;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = ~n2382 & n2385;
  assign n2387 = n2382 & ~n2385;
  assign s231 = ~n2386 & ~n2387;
  assign n2389 = ~n2383 & ~n2386;
  assign n2390 = a232 & b232;
  assign n2391 = ~a232 & ~b232;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2389 & n2392;
  assign n2394 = n2389 & ~n2392;
  assign s232 = ~n2393 & ~n2394;
  assign n2396 = ~n2390 & ~n2393;
  assign n2397 = a233 & b233;
  assign n2398 = ~a233 & ~b233;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = ~n2396 & n2399;
  assign n2401 = n2396 & ~n2399;
  assign s233 = ~n2400 & ~n2401;
  assign n2403 = ~n2397 & ~n2400;
  assign n2404 = a234 & b234;
  assign n2405 = ~a234 & ~b234;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~n2403 & n2406;
  assign n2408 = n2403 & ~n2406;
  assign s234 = ~n2407 & ~n2408;
  assign n2410 = ~n2404 & ~n2407;
  assign n2411 = a235 & b235;
  assign n2412 = ~a235 & ~b235;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2410 & n2413;
  assign n2415 = n2410 & ~n2413;
  assign s235 = ~n2414 & ~n2415;
  assign n2417 = ~n2411 & ~n2414;
  assign n2418 = a236 & b236;
  assign n2419 = ~a236 & ~b236;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = ~n2417 & n2420;
  assign n2422 = n2417 & ~n2420;
  assign s236 = ~n2421 & ~n2422;
  assign n2424 = ~n2418 & ~n2421;
  assign n2425 = a237 & b237;
  assign n2426 = ~a237 & ~b237;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = ~n2424 & n2427;
  assign n2429 = n2424 & ~n2427;
  assign s237 = ~n2428 & ~n2429;
  assign n2431 = ~n2425 & ~n2428;
  assign n2432 = a238 & b238;
  assign n2433 = ~a238 & ~b238;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = ~n2431 & n2434;
  assign n2436 = n2431 & ~n2434;
  assign s238 = ~n2435 & ~n2436;
  assign n2438 = ~n2432 & ~n2435;
  assign n2439 = a239 & b239;
  assign n2440 = ~a239 & ~b239;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = ~n2438 & n2441;
  assign n2443 = n2438 & ~n2441;
  assign s239 = ~n2442 & ~n2443;
  assign n2445 = ~n2439 & ~n2442;
  assign n2446 = a240 & b240;
  assign n2447 = ~a240 & ~b240;
  assign n2448 = ~n2446 & ~n2447;
  assign n2449 = ~n2445 & n2448;
  assign n2450 = n2445 & ~n2448;
  assign s240 = ~n2449 & ~n2450;
  assign n2452 = ~n2446 & ~n2449;
  assign n2453 = a241 & b241;
  assign n2454 = ~a241 & ~b241;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = ~n2452 & n2455;
  assign n2457 = n2452 & ~n2455;
  assign s241 = ~n2456 & ~n2457;
  assign n2459 = ~n2453 & ~n2456;
  assign n2460 = a242 & b242;
  assign n2461 = ~a242 & ~b242;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = ~n2459 & n2462;
  assign n2464 = n2459 & ~n2462;
  assign s242 = ~n2463 & ~n2464;
  assign n2466 = ~n2460 & ~n2463;
  assign n2467 = a243 & b243;
  assign n2468 = ~a243 & ~b243;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = ~n2466 & n2469;
  assign n2471 = n2466 & ~n2469;
  assign s243 = ~n2470 & ~n2471;
  assign n2473 = ~n2467 & ~n2470;
  assign n2474 = a244 & b244;
  assign n2475 = ~a244 & ~b244;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = ~n2473 & n2476;
  assign n2478 = n2473 & ~n2476;
  assign s244 = ~n2477 & ~n2478;
  assign n2480 = ~n2474 & ~n2477;
  assign n2481 = a245 & b245;
  assign n2482 = ~a245 & ~b245;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = ~n2480 & n2483;
  assign n2485 = n2480 & ~n2483;
  assign s245 = ~n2484 & ~n2485;
  assign n2487 = ~n2481 & ~n2484;
  assign n2488 = a246 & b246;
  assign n2489 = ~a246 & ~b246;
  assign n2490 = ~n2488 & ~n2489;
  assign n2491 = ~n2487 & n2490;
  assign n2492 = n2487 & ~n2490;
  assign s246 = ~n2491 & ~n2492;
  assign n2494 = ~n2488 & ~n2491;
  assign n2495 = a247 & b247;
  assign n2496 = ~a247 & ~b247;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2494 & n2497;
  assign n2499 = n2494 & ~n2497;
  assign s247 = ~n2498 & ~n2499;
  assign n2501 = ~n2495 & ~n2498;
  assign n2502 = a248 & b248;
  assign n2503 = ~a248 & ~b248;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2501 & n2504;
  assign n2506 = n2501 & ~n2504;
  assign s248 = ~n2505 & ~n2506;
  assign n2508 = ~n2502 & ~n2505;
  assign n2509 = a249 & b249;
  assign n2510 = ~a249 & ~b249;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = ~n2508 & n2511;
  assign n2513 = n2508 & ~n2511;
  assign s249 = ~n2512 & ~n2513;
  assign n2515 = ~n2509 & ~n2512;
  assign n2516 = a250 & b250;
  assign n2517 = ~a250 & ~b250;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2515 & n2518;
  assign n2520 = n2515 & ~n2518;
  assign s250 = ~n2519 & ~n2520;
  assign n2522 = ~n2516 & ~n2519;
  assign n2523 = a251 & b251;
  assign n2524 = ~a251 & ~b251;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = ~n2522 & n2525;
  assign n2527 = n2522 & ~n2525;
  assign s251 = ~n2526 & ~n2527;
  assign n2529 = ~n2523 & ~n2526;
  assign n2530 = a252 & b252;
  assign n2531 = ~a252 & ~b252;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = ~n2529 & n2532;
  assign n2534 = n2529 & ~n2532;
  assign s252 = ~n2533 & ~n2534;
  assign n2536 = ~n2530 & ~n2533;
  assign n2537 = a253 & b253;
  assign n2538 = ~a253 & ~b253;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = ~n2536 & n2539;
  assign n2541 = n2536 & ~n2539;
  assign s253 = ~n2540 & ~n2541;
  assign n2543 = ~n2537 & ~n2540;
  assign n2544 = a254 & b254;
  assign n2545 = ~a254 & ~b254;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = ~n2543 & n2546;
  assign n2548 = n2543 & ~n2546;
  assign s254 = ~n2547 & ~n2548;
  assign n2550 = ~n2544 & ~n2547;
  assign n2551 = a255 & b255;
  assign n2552 = ~a255 & ~b255;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~n2550 & n2553;
  assign n2555 = n2550 & ~n2553;
  assign s255 = ~n2554 & ~n2555;
  assign s256 = n2551 | n2554;
endmodule


