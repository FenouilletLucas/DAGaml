// Benchmark "vda" written by ABC on Tue May 16 16:07:53 2017

module vda ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q,
    r, s, t, u, v, w, x, y, z, a0, a1, b0, b1, c0, c1, d0, d1, e0, f0, g0,
    h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0,
    z0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q;
  output r, s, t, u, v, w, x, y, z, a0, a1, b0, b1, c0, c1, d0, d1, e0, f0,
    g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0,
    y0, z0;
  wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n170, n171, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n198,
    n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n213, n214, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n231, n233, n234, n235, n239, n240, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n438, n439, n440, n441, n442, n444, n445,
    n446, n447, n448, n449, n450, n452, n453, n454, n455, n456, n457, n458,
    n460, n461, n462, n463, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n476, n477, n478, n479, n481, n482, n483, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n496, n497, n498, n499, n500, n501,
    n502, n503, n505, n506, n507, n509, n510, n511, n512, n514, n516, n517,
    n519, n520, n521, n522, n523, n524;
  assign n57 = ~l & p;
  assign n58 = n & n57;
  assign n59 = ~o & n58;
  assign n60 = ~m & ~q;
  assign n61 = ~f & n60;
  assign n62 = n59 & n61;
  assign n63 = f & n60;
  assign n64 = n59 & n63;
  assign n65 = ~n62 & ~n64;
  assign n66 = n & ~o;
  assign n67 = ~l & ~p;
  assign n68 = n60 & n67;
  assign n69 = n66 & n68;
  assign n70 = n65 & ~n69;
  assign n71 = m & ~q;
  assign n72 = n67 & n71;
  assign n73 = ~n & o;
  assign n74 = o & n58;
  assign n75 = ~m & q;
  assign n76 = g & n75;
  assign n77 = n74 & n76;
  assign n78 = g & n73;
  assign n79 = n72 & n78;
  assign n80 = ~n77 & ~n79;
  assign n81 = l & p;
  assign n82 = n75 & n81;
  assign n83 = n78 & n82;
  assign n84 = ~n & ~o;
  assign n85 = n57 & n84;
  assign n86 = n60 & n85;
  assign n87 = ~l & n73;
  assign z = n60 & n87;
  assign n89 = ~n86 & ~z;
  assign n90 = l & ~p;
  assign n91 = n66 & n90;
  assign n92 = n71 & n91;
  assign n93 = n72 & n84;
  assign n94 = ~n92 & ~n93;
  assign n95 = n57 & n73;
  assign n96 = m & q;
  assign n97 = n95 & n96;
  assign n98 = n94 & ~n97;
  assign n99 = n & o;
  assign n100 = ~p & n60;
  assign n101 = n99 & n100;
  assign n102 = ~l & n60;
  assign n103 = n99 & n102;
  assign n104 = n73 & n90;
  assign n105 = n71 & n104;
  assign n106 = n101 & n103;
  assign n107 = ~n105 & ~n106;
  assign n108 = n81 & n84;
  assign n109 = n96 & n108;
  assign n110 = n59 & n75;
  assign n111 = i & n110;
  assign n112 = ~n109 & ~n111;
  assign n113 = n107 & n112;
  assign n114 = n98 & n113;
  assign n115 = n81 & n96;
  assign n116 = n66 & n115;
  assign n117 = n75 & n84;
  assign n118 = n57 & n117;
  assign n119 = ~b & f;
  assign n120 = n118 & n119;
  assign n121 = ~n116 & ~n120;
  assign n122 = n71 & n95;
  assign n123 = ~g & n96;
  assign n124 = n59 & n123;
  assign n125 = ~g & n122;
  assign n126 = ~n124 & ~n125;
  assign n127 = n75 & n104;
  assign n128 = n126 & ~n127;
  assign n129 = n121 & n128;
  assign n130 = n114 & n129;
  assign n131 = e & h;
  assign n132 = ~i & n71;
  assign n133 = n74 & n132;
  assign n134 = ~f & j;
  assign n135 = n133 & n134;
  assign n136 = n131 & n135;
  assign n137 = ~c & j;
  assign n138 = n133 & n137;
  assign n139 = n131 & n138;
  assign n140 = b & j;
  assign n141 = n133 & n140;
  assign n142 = n131 & n141;
  assign n143 = ~n139 & ~n142;
  assign n144 = ~n136 & n143;
  assign n145 = n60 & n81;
  assign n146 = n84 & n145;
  assign n147 = n144 & ~n146;
  assign n148 = a & n60;
  assign n149 = e & n104;
  assign n150 = n148 & n149;
  assign n151 = e & ~n120;
  assign n152 = n118 & n151;
  assign n153 = ~n150 & ~n152;
  assign n154 = n67 & n75;
  assign n155 = n73 & n154;
  assign n156 = n153 & ~n155;
  assign n157 = n73 & n145;
  assign n158 = c & n67;
  assign n159 = n117 & n158;
  assign n160 = ~n157 & ~n159;
  assign n161 = n99 & n154;
  assign n162 = ~g & n73;
  assign n163 = n82 & n162;
  assign n164 = ~n161 & ~n163;
  assign n165 = n160 & n164;
  assign n166 = n156 & n165;
  assign n167 = n147 & n166;
  assign n168 = n130 & n167;
  assign t = ~n89 | ~n168;
  assign n170 = ~n83 & ~t;
  assign n171 = n80 & n170;
  assign r = ~n70 | ~n171;
  assign n173 = h & n99;
  assign n174 = n72 & n173;
  assign n175 = ~b & c;
  assign n176 = f & n175;
  assign n177 = h & n176;
  assign n178 = n133 & n177;
  assign n179 = ~l & ~n178;
  assign n180 = ~n174 & n179;
  assign n181 = n99 & n180;
  assign n182 = n132 & n181;
  assign n183 = ~n131 & n182;
  assign n184 = ~e & ~f;
  assign n185 = n104 & n184;
  assign n186 = n148 & n185;
  assign n187 = n99 & ~n174;
  assign n188 = n72 & n187;
  assign n189 = n99 & n145;
  assign n190 = ~n188 & ~n189;
  assign n191 = ~n186 & n190;
  assign n192 = ~n183 & n191;
  assign n193 = n60 & n84;
  assign n194 = n67 & n193;
  assign n195 = p & n184;
  assign n196 = n117 & n195;
  assign a1 = n81 & n117;
  assign n198 = ~n196 & ~a1;
  assign n199 = ~n194 & n198;
  assign s = ~n192 | ~n199;
  assign n201 = n96 & n104;
  assign n202 = n82 & n99;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~o & n67;
  assign n205 = n96 & n204;
  assign n206 = n & n205;
  assign n207 = n & n75;
  assign n208 = n90 & n207;
  assign n209 = ~o & n208;
  assign n210 = ~n206 & ~n209;
  assign n211 = n71 & n85;
  assign c0 = n66 & n154;
  assign n213 = ~n211 & ~c0;
  assign n214 = n210 & n213;
  assign u = ~n203 | ~n214;
  assign n216 = d & ~i;
  assign n217 = n110 & n216;
  assign n218 = g & k;
  assign n219 = n122 & n218;
  assign n220 = g & i;
  assign n221 = n122 & n220;
  assign n222 = c & g;
  assign n223 = n122 & n222;
  assign n224 = ~n221 & ~n223;
  assign n225 = ~n219 & n224;
  assign n226 = ~n217 & n225;
  assign n227 = ~d & ~i;
  assign n228 = n110 & n227;
  assign n229 = ~k & n75;
  assign b0 = n95 & n229;
  assign n231 = ~c0 & ~b0;
  assign a0 = ~n80 | ~n231;
  assign n233 = ~u & ~a0;
  assign n234 = ~n83 & n233;
  assign n235 = ~n228 & n234;
  assign y = ~n226 | ~n235;
  assign v = n69 | y;
  assign b1 = j & n174;
  assign n239 = n90 & n193;
  assign n240 = n74 & n96;
  assign c1 = n239 | n240;
  assign n242 = ~n105 & ~n157;
  assign n243 = n85 & n96;
  assign n244 = n242 & ~n243;
  assign n245 = ~n178 & n244;
  assign n246 = n60 & n91;
  assign n247 = n245 & ~n246;
  assign n248 = n71 & n90;
  assign n249 = n99 & n248;
  assign n250 = n192 & ~n249;
  assign n251 = n67 & n73;
  assign n252 = n96 & n251;
  assign n253 = ~n103 & ~n252;
  assign n254 = ~a & n104;
  assign n255 = ~n196 & ~n254;
  assign d1 = n91 & n96;
  assign n257 = ~a1 & ~d1;
  assign n258 = ~n & n71;
  assign n259 = n81 & n258;
  assign n260 = l & n71;
  assign n261 = n84 & n260;
  assign n262 = n84 & n90;
  assign n263 = n96 & n262;
  assign n264 = k & n75;
  assign n265 = n95 & n264;
  assign z0 = n90 & n117;
  assign n267 = p & n71;
  assign n268 = n66 & n267;
  assign n269 = ~n83 & ~z0;
  assign n270 = ~n120 & n269;
  assign n271 = ~n163 & n270;
  assign n272 = ~n127 & n271;
  assign n273 = ~n92 & n272;
  assign n274 = ~n109 & n273;
  assign n275 = ~n265 & n274;
  assign n276 = ~n263 & n275;
  assign n277 = ~n261 & n276;
  assign n278 = ~n259 & n277;
  assign n279 = ~n239 & n278;
  assign n280 = n147 & n279;
  assign n281 = n257 & n280;
  assign n282 = n203 & n281;
  assign n283 = n255 & n282;
  assign n284 = n253 & n283;
  assign n285 = n250 & n284;
  assign n286 = n247 & n285;
  assign d0 = n268 | ~n286;
  assign n288 = ~g & q;
  assign n289 = n74 & n288;
  assign n290 = n72 & n162;
  assign n291 = g & n58;
  assign n292 = n96 & n291;
  assign n293 = ~n174 & ~n289;
  assign n294 = ~n292 & n293;
  assign n295 = ~n290 & n294;
  assign n296 = ~f & ~j;
  assign n297 = m & n296;
  assign n298 = n74 & n297;
  assign n299 = n131 & n298;
  assign n300 = ~c & ~j;
  assign n301 = m & n300;
  assign n302 = n74 & n301;
  assign n303 = n131 & n302;
  assign n304 = b & ~j;
  assign n305 = m & n304;
  assign n306 = n74 & n305;
  assign n307 = n131 & n306;
  assign n308 = ~c & g;
  assign n309 = ~k & n308;
  assign n310 = n132 & n309;
  assign n311 = n95 & n310;
  assign n312 = ~n307 & ~n311;
  assign n313 = ~n303 & n312;
  assign n314 = ~n299 & n313;
  assign n315 = n66 & n145;
  assign n316 = n314 & ~n315;
  assign n317 = i & n71;
  assign n318 = n74 & n317;
  assign n319 = ~n101 & ~n318;
  assign n320 = n66 & n72;
  assign n321 = n319 & ~n320;
  assign n322 = ~n211 & ~n228;
  assign n323 = ~n62 & ~n163;
  assign n324 = ~n109 & n323;
  assign n325 = ~n178 & n324;
  assign n326 = ~n265 & n325;
  assign n327 = ~n261 & n326;
  assign n328 = ~n259 & n327;
  assign n329 = ~n208 & n328;
  assign n330 = ~n205 & n329;
  assign n331 = n126 & n330;
  assign n332 = n80 & n331;
  assign n333 = n98 & n332;
  assign n334 = n322 & n333;
  assign n335 = n257 & n334;
  assign n336 = n203 & n335;
  assign n337 = n321 & n336;
  assign n338 = n316 & n337;
  assign e0 = ~n295 | ~n338;
  assign n340 = ~e & f;
  assign n341 = l & n340;
  assign n342 = n73 & n341;
  assign n343 = n148 & n342;
  assign n344 = b & ~e;
  assign n345 = f & n344;
  assign n346 = n118 & n345;
  assign n347 = ~n343 & ~n346;
  assign n348 = n59 & n71;
  assign n349 = ~n239 & ~n348;
  assign n350 = ~n83 & n164;
  assign n351 = n66 & n82;
  assign n352 = ~n97 & ~n111;
  assign n353 = ~n116 & n352;
  assign n354 = ~n206 & n353;
  assign n355 = ~n351 & n354;
  assign n356 = n226 & n355;
  assign n357 = n350 & n356;
  assign n358 = n70 & n357;
  assign n359 = n257 & n358;
  assign n360 = n314 & n359;
  assign n361 = n231 & n360;
  assign n362 = n253 & n361;
  assign n363 = n349 & n362;
  assign n364 = n347 & n363;
  assign n365 = n321 & n364;
  assign n366 = n247 & n365;
  assign f0 = ~n295 | ~n366;
  assign n368 = m & n73;
  assign n369 = n81 & n368;
  assign n370 = ~n263 & ~n351;
  assign n371 = ~n369 & n370;
  assign n372 = ~n201 & n226;
  assign n373 = ~z & n372;
  assign n374 = ~n62 & ~a1;
  assign n375 = ~n228 & n374;
  assign n376 = ~n259 & n375;
  assign n377 = ~n208 & n376;
  assign n378 = ~n318 & n377;
  assign n379 = n112 & n378;
  assign n380 = n129 & n379;
  assign n381 = n156 & n380;
  assign n382 = n244 & n381;
  assign n383 = n255 & n382;
  assign n384 = n349 & n383;
  assign n385 = n373 & n384;
  assign n386 = n316 & n385;
  assign n387 = n250 & n386;
  assign n388 = n295 & n387;
  assign g0 = ~n371 | ~n388;
  assign n390 = ~b1 & ~z0;
  assign n391 = ~c & ~i;
  assign n392 = n289 & n391;
  assign n393 = p & z;
  assign n394 = ~c0 & ~c1;
  assign n395 = ~d1 & n394;
  assign n396 = ~n155 & n395;
  assign n397 = ~n86 & n396;
  assign n398 = ~n146 & n397;
  assign n399 = ~n161 & n398;
  assign n400 = ~n92 & n399;
  assign n401 = ~n105 & n400;
  assign n402 = ~n211 & n401;
  assign n403 = ~n265 & n402;
  assign n404 = ~n205 & n403;
  assign n405 = n128 & n404;
  assign n406 = n65 & n405;
  assign n407 = n160 & n406;
  assign n408 = n372 & n407;
  assign n409 = n319 & n408;
  assign n410 = n390 & n409;
  assign n411 = n253 & n410;
  assign n412 = n347 & n411;
  assign n413 = n316 & n412;
  assign n414 = n371 & n413;
  assign n415 = ~n393 & n414;
  assign h0 = n392 | ~n415;
  assign n417 = ~c & ~m;
  assign n418 = n84 & n417;
  assign n419 = n67 & n418;
  assign n420 = ~n64 & ~n69;
  assign n421 = ~n161 & n420;
  assign n422 = ~n194 & n421;
  assign n423 = ~n209 & n422;
  assign n424 = ~n261 & n423;
  assign n425 = ~n103 & n424;
  assign n426 = n126 & n425;
  assign n427 = n121 & n426;
  assign n428 = n94 & n427;
  assign n429 = n322 & n428;
  assign n430 = n147 & n429;
  assign n431 = n89 & n430;
  assign n432 = n347 & n431;
  assign n433 = n321 & n432;
  assign n434 = n247 & n433;
  assign n435 = n371 & n434;
  assign i0 = n419 | ~n435;
  assign j0 = n194 | ~n250;
  assign n438 = n130 & n350;
  assign n439 = ~b1 & ~j0;
  assign n440 = ~c1 & n439;
  assign n441 = ~d1 & n440;
  assign n442 = n80 & n441;
  assign k0 = ~n438 | ~n442;
  assign n444 = n70 & ~a0;
  assign n445 = ~n116 & n128;
  assign n446 = n114 & n445;
  assign n447 = n160 & n446;
  assign n448 = n257 & n447;
  assign n449 = n89 & n448;
  assign n450 = n390 & n449;
  assign l0 = ~n444 | ~n450;
  assign n452 = ~n159 & ~c1;
  assign n453 = ~n120 & n452;
  assign n454 = ~n93 & n453;
  assign n455 = n107 & n454;
  assign n456 = n128 & n455;
  assign n457 = n350 & n456;
  assign n458 = n156 & n457;
  assign m0 = ~n89 | ~n458;
  assign n460 = ~n157 & ~c1;
  assign n461 = n257 & n460;
  assign n462 = n390 & n461;
  assign n463 = n438 & n462;
  assign n0 = ~n444 | ~n463;
  assign n465 = n80 & n160;
  assign n466 = ~p & z;
  assign n467 = n153 & ~n466;
  assign n468 = ~b0 & ~j0;
  assign n469 = ~n69 & n468;
  assign n470 = ~n97 & n469;
  assign n471 = n112 & n470;
  assign n472 = n144 & n471;
  assign n473 = n390 & n472;
  assign n474 = n467 & n473;
  assign o0 = ~n465 | ~n474;
  assign n476 = n210 & n322;
  assign n477 = n226 & n476;
  assign n478 = n80 & ~n202;
  assign n479 = n438 & n478;
  assign p0 = ~n477 | ~n479;
  assign n481 = n130 & n147;
  assign n482 = n476 & n481;
  assign n483 = n444 & n482;
  assign q0 = ~n373 | ~n483;
  assign n485 = ~z & ~n97;
  assign n486 = ~n228 & n485;
  assign n487 = n126 & n486;
  assign n488 = n107 & n487;
  assign n489 = n210 & n488;
  assign n490 = n350 & n489;
  assign n491 = n156 & n490;
  assign n492 = n70 & n491;
  assign n493 = n203 & n492;
  assign r0 = ~n231 | ~n493;
  assign s0 = ~n147 | p0;
  assign n496 = ~n69 & ~b0;
  assign n497 = ~n93 & n496;
  assign n498 = ~n127 & n497;
  assign n499 = ~n211 & n498;
  assign n500 = n112 & n499;
  assign n501 = n144 & n500;
  assign n502 = n372 & n501;
  assign n503 = n467 & n502;
  assign t0 = ~n465 | ~n503;
  assign n505 = ~n86 & ~n202;
  assign n506 = n147 & n505;
  assign n507 = n438 & n506;
  assign u0 = ~n465 | ~n507;
  assign n509 = ~n92 & n164;
  assign n510 = n80 & n509;
  assign n511 = n129 & n510;
  assign n512 = n476 & n511;
  assign v0 = ~n373 | ~n512;
  assign n514 = n113 & ~n201;
  assign w0 = ~n156 | ~n514;
  assign n516 = n113 & ~n202;
  assign n517 = n156 & n516;
  assign x0 = ~n477 | ~n517;
  assign n519 = ~n92 & ~c0;
  assign n520 = n121 & n519;
  assign n521 = n164 & n520;
  assign n522 = n113 & n521;
  assign n523 = n65 & n522;
  assign n524 = n467 & n523;
  assign y0 = ~n477 | ~n524;
  assign w = t;
  assign x = t;
endmodule


