// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:38 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_;
  wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n194, n195, n196, n197,
    n198, n199, n200, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
    n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2522,
    n2523, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
    n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3207, n3208, n3209,
    n3210, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3286, n3287, n3288, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3300, n3301, n3302, n3304,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3352, n3353, n3354, n3356, n3357, n3359, n3360,
    n3361, n3362, n3363, n3364, n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3397, n3398, n3399, n3400, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419;
  assign n57 = i_9_ & i_10_;
  assign n58 = ~i_9_ & ~i_10_;
  assign n59 = ~n57 & ~n58;
  assign n60 = ~i_7_ & ~i_8_;
  assign n61 = ~i_6_ & n60;
  assign n62 = i_1_ & ~i_2_;
  assign n63 = ~i_0_ & n62;
  assign n64 = i_3_ & n63;
  assign n65 = ~i_5_ & n64;
  assign n66 = n61 & n65;
  assign n67 = ~n59 & n66;
  assign n68 = ~i_12_ & i_13_;
  assign n69 = ~i_14_ & n68;
  assign n70 = ~i_9_ & i_10_;
  assign n71 = ~i_11_ & n70;
  assign n72 = i_15_ & n71;
  assign n73 = i_9_ & ~i_10_;
  assign n74 = ~i_11_ & n73;
  assign n75 = i_15_ & n74;
  assign n76 = ~n72 & ~n75;
  assign n77 = n69 & ~n76;
  assign n78 = ~i_12_ & ~i_13_;
  assign n79 = i_14_ & n78;
  assign n80 = ~n76 & n79;
  assign n81 = ~n77 & ~n80;
  assign n82 = i_14_ & n68;
  assign n83 = ~i_11_ & ~i_12_;
  assign n84 = ~n82 & n83;
  assign n85 = n59 & ~n84;
  assign n86 = ~i_14_ & n78;
  assign n87 = ~i_15_ & n71;
  assign n88 = n86 & n87;
  assign n89 = ~n85 & ~n88;
  assign n90 = n81 & n89;
  assign n91 = ~i_11_ & n57;
  assign n92 = i_12_ & n91;
  assign n93 = n90 & ~n92;
  assign n94 = ~i_3_ & i_4_;
  assign n95 = ~i_5_ & n94;
  assign n96 = n63 & n95;
  assign n97 = n60 & n96;
  assign n98 = ~n93 & n97;
  assign n99 = i_5_ & n94;
  assign n100 = n63 & n99;
  assign n101 = ~i_3_ & ~i_4_;
  assign n102 = i_5_ & n101;
  assign n103 = n63 & n102;
  assign n104 = ~n100 & ~n103;
  assign n105 = i_6_ & i_8_;
  assign n106 = ~n104 & n105;
  assign n107 = i_11_ & n73;
  assign n108 = ~n57 & ~n107;
  assign n109 = i_6_ & i_7_;
  assign n110 = ~i_8_ & n109;
  assign n111 = ~i_5_ & n101;
  assign n112 = ~i_0_ & ~i_1_;
  assign n113 = ~i_2_ & n112;
  assign n114 = n111 & n113;
  assign n115 = n110 & n114;
  assign n116 = ~n108 & n115;
  assign n117 = i_0_ & n62;
  assign n118 = ~n102 & n117;
  assign o_6_ = i_3_ & n112;
  assign n120 = ~n118 & ~o_6_;
  assign n121 = ~n116 & n120;
  assign n122 = ~n106 & n121;
  assign n123 = ~n98 & n122;
  assign n124 = ~n67 & n123;
  assign n125 = i_6_ & ~i_8_;
  assign n126 = ~n104 & n125;
  assign n127 = ~i_15_ & n74;
  assign n128 = n86 & n127;
  assign n129 = n59 & n90;
  assign n130 = ~n128 & n129;
  assign n131 = n126 & ~n130;
  assign n132 = i_7_ & n131;
  assign n133 = n124 & ~n132;
  assign n134 = ~i_6_ & ~i_7_;
  assign n135 = i_8_ & n134;
  assign n136 = n63 & n111;
  assign n137 = n135 & n136;
  assign n138 = ~i_7_ & n105;
  assign n139 = n136 & n138;
  assign n140 = ~n137 & ~n139;
  assign n141 = ~i_11_ & n58;
  assign n142 = i_15_ & n141;
  assign n143 = n86 & n142;
  assign n144 = ~n76 & n86;
  assign n145 = ~i_11_ & i_12_;
  assign n146 = n59 & n145;
  assign n147 = ~n68 & ~n79;
  assign n148 = ~n146 & n147;
  assign n149 = i_11_ & n70;
  assign n150 = n108 & ~n149;
  assign n151 = n148 & n150;
  assign n152 = ~n144 & n151;
  assign n153 = i_11_ & n58;
  assign n154 = ~i_12_ & ~n153;
  assign n155 = n152 & n154;
  assign n156 = ~n143 & n155;
  assign n157 = ~n140 & ~n156;
  assign n158 = n96 & n138;
  assign n159 = n96 & n135;
  assign n160 = ~n158 & ~n159;
  assign n161 = ~n58 & n152;
  assign n162 = ~n160 & ~n161;
  assign n163 = ~n157 & ~n162;
  assign n164 = n133 & n163;
  assign o_14_ = i_0_ & ~i_1_;
  assign n166 = n102 & o_14_;
  assign n167 = n79 & n87;
  assign n168 = n72 & n86;
  assign n169 = n69 & n87;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n167 & n170;
  assign n172 = ~i_15_ & n91;
  assign n173 = n68 & n172;
  assign n174 = ~i_14_ & n173;
  assign n175 = i_15_ & n91;
  assign n176 = n86 & n175;
  assign n177 = ~n174 & ~n176;
  assign n178 = n171 & n177;
  assign n179 = n79 & n172;
  assign n180 = n75 & n86;
  assign n181 = n69 & n127;
  assign n182 = ~n180 & ~n181;
  assign n183 = n79 & n127;
  assign n184 = n182 & ~n183;
  assign n185 = ~n179 & n184;
  assign n186 = n178 & n185;
  assign n187 = ~n58 & n186;
  assign n188 = n125 & ~n187;
  assign n189 = ~n109 & ~n188;
  assign n190 = n136 & ~n189;
  assign n191 = ~n166 & ~n190;
  assign n192 = ~n139 & n191;
  assign o_2_ = n164 & ~n192;
  assign n194 = ~i_6_ & i_7_;
  assign n195 = n61 & ~n187;
  assign n196 = ~n194 & ~n195;
  assign n197 = n63 & ~n196;
  assign n198 = ~o_14_ & ~n197;
  assign n199 = n111 & ~n198;
  assign n200 = ~n137 & ~n199;
  assign o_7_ = n164 & ~n200;
  assign o_0_ = o_2_ | o_7_;
  assign n203 = n58 & n97;
  assign n204 = n94 & o_14_;
  assign n205 = n125 & ~n186;
  assign n206 = ~n109 & ~n205;
  assign n207 = n96 & ~n206;
  assign n208 = n61 & ~n186;
  assign n209 = ~n194 & ~n208;
  assign n210 = n96 & ~n209;
  assign n211 = ~n207 & ~n210;
  assign n212 = ~n204 & n211;
  assign n213 = n160 & n212;
  assign n214 = ~n203 & n213;
  assign o_1_ = n164 & ~n214;
  assign n216 = n95 & n113;
  assign n217 = ~i_6_ & n216;
  assign n218 = ~i_8_ & n217;
  assign n219 = i_7_ & n218;
  assign n220 = n82 & n127;
  assign n221 = n115 & n220;
  assign n222 = ~n219 & ~n221;
  assign n223 = i_12_ & ~i_13_;
  assign n224 = ~i_14_ & n223;
  assign n225 = n91 & n224;
  assign n226 = i_15_ & n225;
  assign n227 = ~n220 & ~n226;
  assign n228 = i_15_ & n153;
  assign n229 = n224 & n228;
  assign n230 = n75 & n223;
  assign n231 = ~i_14_ & n230;
  assign n232 = ~n229 & ~n231;
  assign n233 = ~i_15_ & n153;
  assign n234 = n82 & n233;
  assign n235 = i_15_ & n149;
  assign n236 = n224 & n235;
  assign n237 = ~n234 & ~n236;
  assign n238 = n232 & n237;
  assign n239 = n227 & n238;
  assign n240 = ~n222 & ~n239;
  assign n241 = n102 & n113;
  assign n242 = n134 & n241;
  assign n243 = i_8_ & n242;
  assign n244 = n107 & n224;
  assign n245 = i_15_ & n244;
  assign n246 = n243 & n245;
  assign n247 = ~n240 & ~n246;
  assign n248 = i_6_ & ~i_7_;
  assign n249 = n114 & n248;
  assign n250 = ~n220 & ~n245;
  assign n251 = ~i_8_ & ~n250;
  assign n252 = ~i_15_ & n149;
  assign n253 = n82 & n252;
  assign n254 = ~i_15_ & n107;
  assign n255 = n82 & n254;
  assign n256 = i_11_ & n57;
  assign n257 = n224 & n256;
  assign n258 = i_15_ & n257;
  assign n259 = ~n255 & ~n258;
  assign n260 = i_8_ & ~n259;
  assign n261 = ~n236 & ~n260;
  assign n262 = ~n253 & n261;
  assign n263 = ~n251 & n262;
  assign n264 = n249 & ~n263;
  assign n265 = ~i_8_ & n242;
  assign n266 = n72 & n224;
  assign n267 = ~n236 & ~n266;
  assign n268 = n232 & n267;
  assign n269 = n227 & n268;
  assign n270 = n265 & ~n269;
  assign n271 = n99 & n113;
  assign n272 = n109 & n271;
  assign n273 = i_8_ & n272;
  assign n274 = ~i_8_ & n248;
  assign n275 = n114 & n274;
  assign n276 = ~n273 & ~n275;
  assign n277 = n71 & n82;
  assign n278 = ~i_15_ & n277;
  assign n279 = i_14_ & n173;
  assign n280 = ~n278 & ~n279;
  assign n281 = ~n229 & ~n234;
  assign n282 = n275 & ~n281;
  assign n283 = n280 & ~n282;
  assign n284 = ~n276 & ~n283;
  assign n285 = ~n270 & ~n284;
  assign n286 = ~n264 & n285;
  assign n287 = n247 & n286;
  assign n288 = n194 & n271;
  assign n289 = ~n275 & ~n288;
  assign n290 = ~i_15_ & n256;
  assign n291 = n82 & n290;
  assign n292 = ~i_8_ & n288;
  assign n293 = n142 & n224;
  assign n294 = ~i_15_ & n141;
  assign n295 = n82 & n294;
  assign n296 = ~n293 & ~n295;
  assign n297 = ~n231 & ~n255;
  assign n298 = ~n236 & ~n245;
  assign n299 = n281 & n298;
  assign n300 = n297 & n299;
  assign n301 = n296 & n300;
  assign n302 = ~n253 & n301;
  assign n303 = n292 & ~n302;
  assign n304 = ~n291 & ~n303;
  assign n305 = ~n289 & ~n304;
  assign n306 = ~n279 & ~n291;
  assign n307 = n114 & n138;
  assign n308 = i_8_ & n217;
  assign n309 = i_7_ & n308;
  assign n310 = ~n307 & ~n309;
  assign n311 = ~n243 & n310;
  assign n312 = ~n306 & ~n311;
  assign n313 = ~i_8_ & n272;
  assign n314 = ~n265 & ~n313;
  assign n315 = n255 & ~n314;
  assign n316 = ~n288 & ~n313;
  assign n317 = ~n220 & ~n234;
  assign n318 = n313 & ~n317;
  assign n319 = ~n279 & ~n318;
  assign n320 = ~n316 & ~n319;
  assign n321 = ~n315 & ~n320;
  assign n322 = ~n312 & n321;
  assign n323 = ~n258 & ~n266;
  assign n324 = n219 & ~n323;
  assign n325 = n248 & n271;
  assign n326 = ~i_8_ & n325;
  assign n327 = ~n226 & ~n279;
  assign n328 = n326 & ~n327;
  assign n329 = ~n292 & ~n313;
  assign n330 = ~n266 & ~n278;
  assign n331 = ~n329 & ~n330;
  assign n332 = n115 & n278;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n328 & n333;
  assign n335 = ~n324 & n334;
  assign n336 = n322 & n335;
  assign n337 = ~n242 & ~n249;
  assign n338 = ~i_8_ & ~n337;
  assign n339 = ~n288 & ~n338;
  assign n340 = ~n243 & ~n309;
  assign n341 = n339 & n340;
  assign n342 = n258 & ~n341;
  assign n343 = ~n288 & ~n309;
  assign n344 = ~n275 & n343;
  assign n345 = n226 & ~n344;
  assign n346 = n253 & n313;
  assign n347 = n272 & n291;
  assign n348 = n220 & n273;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~n346 & n349;
  assign n351 = ~n345 & n350;
  assign n352 = ~n342 & n351;
  assign n353 = n336 & n352;
  assign n354 = ~n305 & n353;
  assign n355 = n287 & n354;
  assign n356 = ~n243 & ~n272;
  assign n357 = n226 & ~n356;
  assign n358 = i_8_ & n288;
  assign n359 = ~n275 & ~n358;
  assign n360 = n293 & ~n359;
  assign n361 = ~n357 & ~n360;
  assign n362 = n220 & ~n343;
  assign n363 = n361 & ~n362;
  assign n364 = ~n265 & ~n309;
  assign n365 = n234 & ~n364;
  assign n366 = n266 & n275;
  assign n367 = ~n232 & n307;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n365 & n368;
  assign n370 = n245 & ~n310;
  assign n371 = ~n295 & n297;
  assign n372 = n275 & ~n371;
  assign n373 = n243 & ~n267;
  assign n374 = ~n372 & ~n373;
  assign n375 = ~n370 & n374;
  assign n376 = n369 & n375;
  assign n377 = n363 & n376;
  assign n378 = n355 & n377;
  assign n379 = ~i_7_ & n217;
  assign n380 = i_7_ & n217;
  assign n381 = ~n242 & ~n380;
  assign n382 = ~i_8_ & ~n381;
  assign n383 = ~n379 & ~n382;
  assign n384 = ~n253 & ~n278;
  assign n385 = n306 & n384;
  assign n386 = ~n383 & ~n385;
  assign n387 = ~n272 & ~n379;
  assign n388 = ~n236 & ~n258;
  assign n389 = ~n387 & ~n388;
  assign n390 = i_12_ & i_13_;
  assign n391 = i_14_ & n390;
  assign n392 = n233 & n391;
  assign n393 = n290 & n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = n275 & ~n394;
  assign n396 = ~n389 & ~n395;
  assign n397 = ~n386 & n396;
  assign n398 = i_7_ & n105;
  assign n399 = n114 & n398;
  assign n400 = ~n382 & n387;
  assign n401 = ~n399 & n400;
  assign n402 = n293 & ~n401;
  assign n403 = ~n227 & n379;
  assign n404 = ~n115 & ~n379;
  assign n405 = ~n313 & n404;
  assign n406 = n229 & ~n405;
  assign n407 = n266 & n273;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n403 & n408;
  assign n410 = ~n402 & n409;
  assign n411 = ~n207 & n410;
  assign n412 = n223 & n294;
  assign n413 = i_14_ & n412;
  assign n414 = ~n275 & ~n292;
  assign n415 = n413 & ~n414;
  assign n416 = n96 & n274;
  assign n417 = n58 & n416;
  assign n418 = ~n158 & ~n417;
  assign n419 = ~n415 & n418;
  assign n420 = n411 & n419;
  assign n421 = n397 & n420;
  assign n422 = n268 & n296;
  assign n423 = n309 & ~n422;
  assign n424 = n105 & n271;
  assign n425 = ~i_7_ & n424;
  assign n426 = ~n330 & n425;
  assign n427 = ~n249 & ~n288;
  assign n428 = i_8_ & ~n427;
  assign n429 = ~n330 & n428;
  assign n430 = i_8_ & ~n337;
  assign n431 = ~n220 & ~n293;
  assign n432 = n430 & ~n431;
  assign n433 = ~n429 & ~n432;
  assign n434 = ~n426 & n433;
  assign n435 = ~n423 & n434;
  assign n436 = n232 & n384;
  assign n437 = n243 & ~n436;
  assign n438 = ~n295 & ~n437;
  assign n439 = ~n242 & ~n288;
  assign n440 = i_8_ & ~n439;
  assign n441 = ~n273 & ~n307;
  assign n442 = ~n399 & n441;
  assign n443 = ~n440 & n442;
  assign n444 = ~n438 & ~n443;
  assign n445 = n234 & ~n441;
  assign n446 = ~n300 & n358;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n444 & n447;
  assign n449 = n435 & n448;
  assign n450 = i_14_ & n223;
  assign n451 = n172 & n450;
  assign n452 = n127 & n223;
  assign n453 = i_14_ & n452;
  assign n454 = ~n451 & ~n453;
  assign n455 = n309 & ~n454;
  assign n456 = n87 & n223;
  assign n457 = i_14_ & n456;
  assign n458 = ~n392 & ~n412;
  assign n459 = ~n457 & n458;
  assign n460 = n307 & ~n459;
  assign n461 = ~n455 & ~n460;
  assign n462 = ~n340 & n457;
  assign n463 = i_15_ & n107;
  assign n464 = n450 & n463;
  assign n465 = n72 & n450;
  assign n466 = ~n464 & ~n465;
  assign n467 = n358 & ~n466;
  assign n468 = n87 & n390;
  assign n469 = i_14_ & n468;
  assign n470 = n307 & n469;
  assign n471 = ~n467 & ~n470;
  assign n472 = ~i_7_ & n308;
  assign n473 = n223 & n233;
  assign n474 = ~i_14_ & n473;
  assign n475 = ~n234 & ~n474;
  assign n476 = n472 & ~n475;
  assign n477 = n471 & ~n476;
  assign n478 = n229 & n273;
  assign n479 = n226 & n307;
  assign n480 = ~n478 & ~n479;
  assign n481 = n79 & n233;
  assign n482 = ~n234 & ~n481;
  assign n483 = n243 & ~n482;
  assign n484 = n358 & n413;
  assign n485 = ~n483 & ~n484;
  assign n486 = n480 & n485;
  assign n487 = n477 & n486;
  assign n488 = ~n462 & n487;
  assign n489 = n461 & n488;
  assign n490 = n449 & n489;
  assign n491 = n218 & ~n454;
  assign n492 = n294 & n391;
  assign n493 = n358 & n492;
  assign n494 = n79 & n254;
  assign n495 = ~n265 & ~n379;
  assign n496 = n494 & ~n495;
  assign n497 = ~n493 & ~n496;
  assign n498 = ~n491 & n497;
  assign n499 = n490 & n498;
  assign n500 = n421 & n499;
  assign n501 = n378 & n500;
  assign n502 = ~n465 & ~n469;
  assign n503 = n425 & ~n502;
  assign n504 = n142 & n450;
  assign n505 = n256 & n450;
  assign n506 = i_15_ & n505;
  assign n507 = n175 & n450;
  assign n508 = ~n506 & ~n507;
  assign n509 = n228 & n450;
  assign n510 = i_14_ & n230;
  assign n511 = ~n509 & ~n510;
  assign n512 = n508 & n511;
  assign n513 = ~n504 & n512;
  assign n514 = n440 & ~n513;
  assign n515 = n235 & n450;
  assign n516 = n358 & n515;
  assign n517 = ~n492 & ~n504;
  assign n518 = n399 & ~n517;
  assign n519 = ~n516 & ~n518;
  assign n520 = ~n514 & n519;
  assign n521 = ~n503 & n520;
  assign n522 = ~n465 & ~n515;
  assign n523 = n252 & n391;
  assign n524 = ~n469 & ~n523;
  assign n525 = n522 & n524;
  assign n526 = ~n492 & n525;
  assign n527 = n243 & ~n526;
  assign n528 = ~n510 & n517;
  assign n529 = ~n310 & ~n528;
  assign n530 = n430 & n464;
  assign n531 = n472 & n510;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~n529 & n532;
  assign n534 = ~n527 & n533;
  assign n535 = ~n441 & n465;
  assign n536 = ~n308 & ~n535;
  assign n537 = ~n509 & ~n515;
  assign n538 = n466 & n537;
  assign n539 = ~n536 & ~n538;
  assign n540 = n508 & n537;
  assign n541 = n307 & ~n540;
  assign n542 = ~n217 & ~n272;
  assign n543 = n507 & ~n542;
  assign n544 = i_8_ & n543;
  assign n545 = ~n541 & ~n544;
  assign n546 = ~n392 & ~n509;
  assign n547 = n425 & ~n546;
  assign n548 = n273 & n492;
  assign n549 = n273 & n392;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n547 & n550;
  assign n552 = n545 & n551;
  assign n553 = ~n539 & n552;
  assign n554 = n534 & n553;
  assign n555 = n521 & n554;
  assign n556 = i_14_ & n473;
  assign n557 = ~n506 & ~n515;
  assign n558 = n252 & n450;
  assign n559 = ~n451 & ~n510;
  assign n560 = ~n558 & n559;
  assign n561 = n557 & n560;
  assign n562 = ~n464 & n561;
  assign n563 = ~n556 & n562;
  assign n564 = n273 & ~n563;
  assign n565 = ~n424 & ~n472;
  assign n566 = n457 & ~n565;
  assign n567 = n194 & n241;
  assign n568 = i_8_ & n567;
  assign n569 = n71 & n568;
  assign n570 = ~i_15_ & n505;
  assign n571 = n273 & n570;
  assign n572 = ~n569 & ~n571;
  assign n573 = ~n358 & ~n472;
  assign n574 = ~n453 & ~n570;
  assign n575 = ~n556 & n574;
  assign n576 = ~n573 & ~n575;
  assign n577 = n216 & n398;
  assign n578 = ~n465 & ~n504;
  assign n579 = n577 & ~n578;
  assign n580 = n141 & n568;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n576 & n581;
  assign n583 = n572 & n582;
  assign n584 = ~n566 & n583;
  assign n585 = ~n564 & n584;
  assign n586 = ~i_14_ & n456;
  assign n587 = ~n167 & ~n586;
  assign n588 = n425 & ~n587;
  assign n589 = ~n494 & n587;
  assign n590 = n358 & ~n589;
  assign n591 = ~n273 & ~n358;
  assign n592 = n481 & ~n591;
  assign n593 = ~n590 & ~n592;
  assign n594 = ~n588 & n593;
  assign n595 = n79 & n294;
  assign n596 = ~i_14_ & n452;
  assign n597 = ~i_15_ & n225;
  assign n598 = n307 & n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = ~n595 & n599;
  assign n601 = ~n310 & ~n600;
  assign n602 = n224 & n252;
  assign n603 = ~n596 & ~n602;
  assign n604 = n440 & ~n603;
  assign n605 = ~n601 & ~n604;
  assign n606 = ~n309 & ~n358;
  assign n607 = ~i_15_ & n257;
  assign n608 = ~n474 & ~n607;
  assign n609 = ~i_14_ & n412;
  assign n610 = ~i_15_ & n244;
  assign n611 = ~n597 & ~n610;
  assign n612 = ~n609 & n611;
  assign n613 = n608 & n612;
  assign n614 = ~n606 & ~n613;
  assign n615 = ~n595 & ~n609;
  assign n616 = ~n243 & ~n399;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~n474 & ~n586;
  assign n619 = n430 & ~n618;
  assign n620 = ~n617 & ~n619;
  assign n621 = ~n614 & n620;
  assign n622 = n605 & n621;
  assign n623 = n594 & n622;
  assign n624 = ~n309 & ~n399;
  assign n625 = ~n273 & n624;
  assign n626 = n413 & ~n625;
  assign n627 = ~n392 & ~n413;
  assign n628 = n243 & ~n627;
  assign n629 = ~n451 & ~n628;
  assign n630 = ~n425 & ~n430;
  assign n631 = ~n472 & n630;
  assign n632 = ~n629 & ~n631;
  assign n633 = ~n626 & ~n632;
  assign n634 = n223 & n254;
  assign n635 = i_14_ & n634;
  assign n636 = ~n558 & ~n570;
  assign n637 = ~n635 & n636;
  assign n638 = n430 & ~n637;
  assign n639 = n135 & n271;
  assign n640 = n595 & n639;
  assign n641 = ~n638 & ~n640;
  assign n642 = ~n586 & ~n602;
  assign n643 = ~n558 & n642;
  assign n644 = ~n556 & n643;
  assign n645 = n309 & ~n644;
  assign n646 = n641 & ~n645;
  assign n647 = n633 & n646;
  assign n648 = n623 & n647;
  assign n649 = n585 & n648;
  assign n650 = n555 & n649;
  assign n651 = n358 & n451;
  assign n652 = ~n313 & ~n651;
  assign n653 = n561 & n642;
  assign n654 = ~n473 & n653;
  assign n655 = ~n652 & ~n654;
  assign n656 = ~n607 & n636;
  assign n657 = ~n393 & n656;
  assign n658 = n292 & ~n657;
  assign n659 = n272 & n597;
  assign n660 = ~n265 & ~n273;
  assign n661 = n453 & ~n660;
  assign n662 = i_14_ & ~n223;
  assign n663 = n233 & n662;
  assign n664 = ~n457 & ~n663;
  assign n665 = n115 & ~n664;
  assign n666 = n110 & n216;
  assign n667 = n507 & n666;
  assign n668 = ~i_8_ & n567;
  assign n669 = n91 & n668;
  assign n670 = ~n667 & ~n669;
  assign n671 = ~n665 & n670;
  assign n672 = ~n661 & n671;
  assign n673 = ~n659 & n672;
  assign n674 = ~n658 & n673;
  assign n675 = ~n655 & n674;
  assign n676 = n127 & n391;
  assign n677 = ~n635 & ~n676;
  assign n678 = ~n392 & ~n469;
  assign n679 = i_14_ & n252;
  assign n680 = ~n393 & ~n679;
  assign n681 = n678 & n680;
  assign n682 = n677 & n681;
  assign n683 = n358 & ~n682;
  assign n684 = ~n509 & n642;
  assign n685 = ~n635 & n684;
  assign n686 = n273 & ~n685;
  assign n687 = ~n683 & ~n686;
  assign n688 = ~n607 & n637;
  assign n689 = n275 & ~n688;
  assign n690 = ~n504 & ~n609;
  assign n691 = ~n400 & ~n690;
  assign n692 = ~n689 & ~n691;
  assign n693 = n687 & n692;
  assign n694 = ~n243 & ~n249;
  assign n695 = ~n115 & n694;
  assign n696 = ~n292 & n695;
  assign n697 = ~n453 & ~n676;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n218 & ~n380;
  assign n700 = ~n265 & n699;
  assign n701 = n570 & ~n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = ~n307 & n356;
  assign n704 = n610 & ~n703;
  assign n705 = n273 & n474;
  assign n706 = ~n704 & ~n705;
  assign n707 = n254 & n391;
  assign n708 = ~n288 & ~n307;
  assign n709 = n707 & ~n708;
  assign n710 = n313 & n596;
  assign n711 = ~n709 & ~n710;
  assign n712 = n706 & n711;
  assign n713 = n702 & n712;
  assign n714 = n693 & n713;
  assign n715 = n675 & n714;
  assign n716 = ~n607 & n677;
  assign n717 = n294 & n662;
  assign n718 = ~n413 & ~n509;
  assign n719 = n313 & ~n718;
  assign n720 = ~n717 & ~n719;
  assign n721 = ~n596 & n611;
  assign n722 = ~n255 & ~n707;
  assign n723 = n721 & n722;
  assign n724 = n720 & n723;
  assign n725 = n716 & n724;
  assign n726 = n379 & ~n725;
  assign n727 = ~n523 & n678;
  assign n728 = n172 & n391;
  assign n729 = ~n393 & ~n728;
  assign n730 = ~n413 & n729;
  assign n731 = n643 & n730;
  assign n732 = n727 & n731;
  assign n733 = ~n383 & ~n732;
  assign n734 = n125 & n271;
  assign n735 = ~n288 & ~n734;
  assign n736 = n313 & n635;
  assign n737 = ~n457 & ~n736;
  assign n738 = ~n735 & ~n737;
  assign n739 = n309 & n506;
  assign n740 = n167 & n639;
  assign n741 = n61 & n271;
  assign n742 = n179 & n741;
  assign n743 = ~n740 & ~n742;
  assign n744 = ~n739 & n743;
  assign n745 = ~n326 & ~n338;
  assign n746 = n451 & ~n745;
  assign n747 = ~n343 & n728;
  assign n748 = ~n746 & ~n747;
  assign n749 = n744 & n748;
  assign n750 = ~n738 & n749;
  assign n751 = ~n733 & n750;
  assign n752 = ~n726 & n751;
  assign n753 = ~n218 & ~n265;
  assign n754 = n696 & n753;
  assign n755 = n556 & ~n754;
  assign n756 = n254 & n662;
  assign n757 = n243 & n756;
  assign n758 = ~n755 & ~n757;
  assign n759 = ~n223 & n679;
  assign n760 = ~n756 & ~n759;
  assign n761 = ~n596 & n760;
  assign n762 = i_8_ & ~n761;
  assign n763 = ~n607 & ~n762;
  assign n764 = n272 & ~n763;
  assign n765 = n758 & ~n764;
  assign n766 = ~n278 & n524;
  assign n767 = ~i_12_ & n679;
  assign n768 = ~n167 & ~n756;
  assign n769 = ~n767 & n768;
  assign n770 = n766 & n769;
  assign n771 = n309 & ~n770;
  assign n772 = ~n717 & ~n756;
  assign n773 = n219 & ~n772;
  assign n774 = ~n771 & ~n773;
  assign n775 = n313 & ~n574;
  assign n776 = n510 & n666;
  assign n777 = n183 & n741;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n775 & n778;
  assign n780 = ~n451 & ~n635;
  assign n781 = n292 & ~n780;
  assign n782 = n74 & n668;
  assign n783 = ~n781 & ~n782;
  assign n784 = n779 & n783;
  assign n785 = ~n265 & ~n380;
  assign n786 = ~n392 & ~n676;
  assign n787 = n309 & ~n786;
  assign n788 = ~n635 & ~n787;
  assign n789 = ~n785 & ~n788;
  assign n790 = ~n314 & ~n720;
  assign n791 = ~n789 & ~n790;
  assign n792 = n784 & n791;
  assign n793 = n774 & n792;
  assign n794 = n765 & n793;
  assign n795 = n752 & n794;
  assign n796 = n715 & n795;
  assign n797 = n650 & n796;
  assign n798 = n79 & n290;
  assign n799 = ~n602 & ~n798;
  assign n800 = n79 & n252;
  assign n801 = ~n607 & ~n800;
  assign n802 = i_8_ & ~n801;
  assign n803 = n799 & ~n802;
  assign n804 = ~n179 & ~n481;
  assign n805 = ~n586 & n804;
  assign n806 = n721 & n805;
  assign n807 = ~i_8_ & ~n806;
  assign n808 = n803 & ~n807;
  assign n809 = n249 & ~n808;
  assign n810 = n183 & ~n660;
  assign n811 = ~n179 & ~n597;
  assign n812 = n326 & ~n811;
  assign n813 = ~n810 & ~n812;
  assign n814 = ~n167 & ~n800;
  assign n815 = ~n183 & n814;
  assign n816 = ~n481 & n815;
  assign n817 = n313 & ~n816;
  assign n818 = n167 & n273;
  assign n819 = n313 & n494;
  assign n820 = ~n818 & ~n819;
  assign n821 = ~n817 & n820;
  assign n822 = n813 & n821;
  assign n823 = ~n809 & n822;
  assign n824 = ~n219 & ~n292;
  assign n825 = ~n494 & n615;
  assign n826 = ~n800 & n825;
  assign n827 = ~n474 & n826;
  assign n828 = ~n481 & n603;
  assign n829 = n587 & n611;
  assign n830 = n828 & n829;
  assign n831 = n827 & n830;
  assign n832 = ~n292 & n721;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n824 & n833;
  assign n835 = n382 & ~n608;
  assign n836 = n219 & n481;
  assign n837 = ~n179 & ~n798;
  assign n838 = n288 & ~n837;
  assign n839 = n265 & n610;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n836 & n840;
  assign n842 = ~n835 & n841;
  assign n843 = n115 & ~n618;
  assign n844 = n242 & n597;
  assign n845 = ~n843 & ~n844;
  assign n846 = n243 & n607;
  assign n847 = ~n115 & ~n265;
  assign n848 = n596 & ~n847;
  assign n849 = ~n846 & ~n848;
  assign n850 = n845 & n849;
  assign n851 = n842 & n850;
  assign n852 = ~n834 & n851;
  assign n853 = n823 & n852;
  assign n854 = n275 & ~n827;
  assign n855 = i_8_ & n595;
  assign n856 = ~n798 & ~n855;
  assign n857 = n272 & ~n856;
  assign n858 = n167 & ~n695;
  assign n859 = ~n217 & ~n265;
  assign n860 = ~n837 & ~n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = ~n857 & n861;
  assign n863 = ~n854 & n862;
  assign n864 = ~n383 & ~n814;
  assign n865 = ~n288 & n695;
  assign n866 = ~n217 & n865;
  assign n867 = n183 & ~n866;
  assign n868 = n307 & n494;
  assign n869 = ~n481 & ~n868;
  assign n870 = n310 & n495;
  assign n871 = ~n869 & ~n870;
  assign n872 = n179 & ~n703;
  assign n873 = n358 & n595;
  assign n874 = ~n798 & ~n800;
  assign n875 = n243 & ~n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = ~n872 & n876;
  assign n878 = ~n871 & n877;
  assign n879 = ~n867 & n878;
  assign n880 = ~n864 & n879;
  assign n881 = n863 & n880;
  assign n882 = n853 & n881;
  assign n883 = ~n507 & n525;
  assign n884 = n292 & ~n883;
  assign n885 = n382 & n507;
  assign n886 = ~n275 & ~n885;
  assign n887 = n508 & ~n523;
  assign n888 = ~n464 & n887;
  assign n889 = ~n886 & ~n888;
  assign n890 = ~n884 & ~n889;
  assign n891 = n218 & n509;
  assign n892 = ~n292 & ~n891;
  assign n893 = ~n506 & n511;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n734 & n753;
  assign n896 = n464 & ~n895;
  assign n897 = ~n894 & ~n896;
  assign n898 = n60 & n217;
  assign n899 = ~n265 & ~n898;
  assign n900 = n465 & ~n899;
  assign n901 = ~n313 & ~n900;
  assign n902 = ~n465 & ~n676;
  assign n903 = ~n507 & ~n728;
  assign n904 = n902 & n903;
  assign n905 = ~n469 & n904;
  assign n906 = ~n901 & ~n905;
  assign n907 = n897 & ~n906;
  assign n908 = n890 & n907;
  assign n909 = ~n523 & ~n728;
  assign n910 = n307 & ~n909;
  assign n911 = ~n338 & ~n898;
  assign n912 = n515 & ~n911;
  assign n913 = ~n510 & ~n676;
  assign n914 = n265 & ~n913;
  assign n915 = ~n707 & ~n728;
  assign n916 = ~n507 & n915;
  assign n917 = n326 & ~n916;
  assign n918 = ~n914 & ~n917;
  assign n919 = ~n912 & n918;
  assign n920 = ~n910 & n919;
  assign n921 = ~n115 & ~n218;
  assign n922 = n510 & ~n921;
  assign n923 = n265 & n506;
  assign n924 = ~n707 & ~n923;
  assign n925 = ~n314 & ~n924;
  assign n926 = ~n922 & ~n925;
  assign n927 = ~n469 & ~n728;
  assign n928 = n273 & ~n927;
  assign n929 = n309 & n393;
  assign n930 = ~n928 & ~n929;
  assign n931 = n926 & n930;
  assign n932 = n920 & n931;
  assign n933 = ~i_8_ & n523;
  assign n934 = ~n393 & ~n933;
  assign n935 = n272 & ~n934;
  assign n936 = n273 & n676;
  assign n937 = ~n935 & ~n936;
  assign n938 = n472 & n506;
  assign n939 = ~n329 & n392;
  assign n940 = ~n938 & ~n939;
  assign n941 = n937 & n940;
  assign n942 = n115 & ~n502;
  assign n943 = ~n509 & ~n942;
  assign n944 = ~n847 & ~n943;
  assign n945 = n557 & n902;
  assign n946 = n219 & ~n945;
  assign n947 = n243 & ~n729;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~n944 & n948;
  assign n950 = n941 & n949;
  assign n951 = n932 & n950;
  assign n952 = n908 & n951;
  assign n953 = ~n508 & n898;
  assign n954 = n511 & n915;
  assign n955 = n502 & n954;
  assign n956 = n275 & ~n955;
  assign n957 = ~n953 & ~n956;
  assign n958 = n292 & n464;
  assign n959 = ~n414 & ~n517;
  assign n960 = n307 & n393;
  assign n961 = ~n959 & ~n960;
  assign n962 = ~n958 & n961;
  assign n963 = n957 & n962;
  assign n964 = n952 & n963;
  assign n965 = ~n475 & n898;
  assign n966 = n231 & n272;
  assign n967 = ~n76 & n224;
  assign n968 = ~n404 & n967;
  assign n969 = ~n966 & ~n968;
  assign n970 = ~n965 & n969;
  assign n971 = n245 & ~n400;
  assign n972 = i_5_ & n204;
  assign n973 = ~n275 & n753;
  assign n974 = n457 & ~n973;
  assign n975 = ~n972 & ~n974;
  assign n976 = ~n971 & n975;
  assign n977 = n970 & n976;
  assign n978 = n964 & n977;
  assign n979 = n882 & n978;
  assign n980 = n797 & n979;
  assign n981 = n501 & n980;
  assign o_3_ = n164 & ~n981;
  assign n983 = n228 & n390;
  assign n984 = i_14_ & n983;
  assign n985 = n400 & n695;
  assign n986 = ~n292 & n985;
  assign n987 = n984 & ~n986;
  assign n988 = ~n537 & n577;
  assign n989 = n639 & n800;
  assign n990 = n481 & n639;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n988 & n991;
  assign n993 = ~n739 & n992;
  assign n994 = n741 & n798;
  assign n995 = n494 & n741;
  assign n996 = ~n994 & ~n995;
  assign n997 = n506 & n666;
  assign n998 = n464 & n666;
  assign n999 = ~n997 & ~n998;
  assign n1000 = n996 & n999;
  assign n1001 = n993 & n1000;
  assign n1002 = ~n987 & n1001;
  assign n1003 = n142 & n391;
  assign n1004 = ~n275 & n383;
  assign n1005 = n329 & n1004;
  assign n1006 = n1003 & ~n1005;
  assign n1007 = ~i_14_ & n390;
  assign n1008 = n172 & n1007;
  assign n1009 = n307 & n1008;
  assign n1010 = n82 & n235;
  assign n1011 = n82 & n228;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = n218 & ~n1012;
  assign n1014 = n79 & n463;
  assign n1015 = ~n707 & ~n1014;
  assign n1016 = i_15_ & n68;
  assign n1017 = n107 & n1016;
  assign n1018 = i_14_ & n1017;
  assign n1019 = n1015 & ~n1018;
  assign n1020 = n307 & ~n1019;
  assign n1021 = ~n1013 & ~n1020;
  assign n1022 = n265 & ~n729;
  assign n1023 = n107 & n1007;
  assign n1024 = ~i_15_ & n1023;
  assign n1025 = n430 & n1024;
  assign n1026 = ~n1022 & ~n1025;
  assign n1027 = n471 & n1026;
  assign n1028 = n1021 & n1027;
  assign n1029 = ~n1009 & n1028;
  assign n1030 = ~n1006 & n1029;
  assign n1031 = n1002 & n1030;
  assign n1032 = n290 & n1007;
  assign n1033 = ~n340 & n1032;
  assign n1034 = ~n275 & ~n1033;
  assign n1035 = n235 & n391;
  assign n1036 = n252 & n1007;
  assign n1037 = ~n1024 & ~n1036;
  assign n1038 = ~n1008 & n1037;
  assign n1039 = i_15_ & n256;
  assign n1040 = n391 & n1039;
  assign n1041 = ~n1032 & ~n1040;
  assign n1042 = n1038 & n1041;
  assign n1043 = ~n1035 & n1042;
  assign n1044 = ~n1034 & ~n1043;
  assign n1045 = n127 & n1007;
  assign n1046 = n294 & n1007;
  assign n1047 = n233 & n1007;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1045 & n1048;
  assign n1050 = ~i_14_ & n983;
  assign n1051 = n75 & n1007;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n1007 & n1039;
  assign n1054 = n235 & n1007;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1052 & n1055;
  assign n1057 = n1049 & n1056;
  assign n1058 = n272 & ~n1057;
  assign n1059 = ~n1044 & ~n1058;
  assign n1060 = n142 & n1007;
  assign n1061 = ~n401 & n1060;
  assign n1062 = n391 & n463;
  assign n1063 = ~n338 & n699;
  assign n1064 = n316 & n1063;
  assign n1065 = ~n326 & n1064;
  assign n1066 = n1062 & ~n1065;
  assign n1067 = i_14_ & ~n390;
  assign n1068 = n142 & n1067;
  assign n1069 = n228 & n1067;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n492 & n1070;
  assign n1072 = ~n1014 & n1071;
  assign n1073 = n313 & ~n1072;
  assign n1074 = ~n1066 & ~n1073;
  assign n1075 = ~n1061 & n1074;
  assign n1076 = n1059 & n1075;
  assign n1077 = ~n404 & ~n1052;
  assign n1078 = n82 & n175;
  assign n1079 = n79 & n175;
  assign n1080 = ~n728 & ~n1079;
  assign n1081 = ~n1008 & n1080;
  assign n1082 = ~n1078 & n1081;
  assign n1083 = n309 & ~n1082;
  assign n1084 = ~n1077 & ~n1083;
  assign n1085 = ~n699 & n1054;
  assign n1086 = n72 & n390;
  assign n1087 = ~i_14_ & n1086;
  assign n1088 = ~n523 & ~n707;
  assign n1089 = ~n1087 & n1088;
  assign n1090 = n273 & ~n1089;
  assign n1091 = ~n1085 & ~n1090;
  assign n1092 = n326 & n984;
  assign n1093 = n107 & n668;
  assign n1094 = n256 & n668;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n1092 & n1095;
  assign n1097 = n1091 & n1096;
  assign n1098 = n1084 & n1097;
  assign n1099 = ~i_14_ & n468;
  assign n1100 = ~n1047 & ~n1099;
  assign n1101 = n1037 & n1100;
  assign n1102 = ~n358 & ~n1047;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n606 & n1103;
  assign n1105 = n79 & n142;
  assign n1106 = ~n1046 & ~n1105;
  assign n1107 = n79 & n235;
  assign n1108 = ~n1036 & ~n1107;
  assign n1109 = n243 & ~n1108;
  assign n1110 = n1106 & ~n1109;
  assign n1111 = ~n309 & n616;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n79 & n228;
  assign n1114 = ~n1047 & ~n1113;
  assign n1115 = n425 & ~n1114;
  assign n1116 = ~n1112 & ~n1115;
  assign n1117 = ~n1104 & n1116;
  assign n1118 = n249 & ~n1106;
  assign n1119 = n358 & n1045;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = n786 & ~n1086;
  assign n1122 = ~n695 & ~n1121;
  assign n1123 = n79 & n1039;
  assign n1124 = ~n242 & ~n307;
  assign n1125 = n1123 & ~n1124;
  assign n1126 = n75 & n391;
  assign n1127 = n273 & n1126;
  assign n1128 = ~n1125 & ~n1127;
  assign n1129 = ~n1122 & n1128;
  assign n1130 = n1120 & n1129;
  assign n1131 = n1117 & n1130;
  assign n1132 = n1098 & n1131;
  assign n1133 = n555 & n1132;
  assign n1134 = n1076 & n1133;
  assign n1135 = n1031 & n1134;
  assign n1136 = n964 & n1135;
  assign n1137 = n75 & n79;
  assign n1138 = ~n676 & ~n1137;
  assign n1139 = n175 & n1007;
  assign n1140 = ~n1087 & ~n1139;
  assign n1141 = ~n393 & ~n1123;
  assign n1142 = ~n1053 & n1141;
  assign n1143 = ~n1014 & ~n1079;
  assign n1144 = n915 & n1143;
  assign n1145 = n1142 & n1144;
  assign n1146 = n1140 & n1145;
  assign n1147 = n1138 & n1146;
  assign n1148 = n379 & ~n1147;
  assign n1149 = ~n696 & n1126;
  assign n1150 = n338 & ~n1143;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1148 & n1151;
  assign n1153 = ~n313 & n383;
  assign n1154 = i_14_ & n1086;
  assign n1155 = ~n1035 & ~n1154;
  assign n1156 = ~n1153 & ~n1155;
  assign n1157 = i_15_ & n1023;
  assign n1158 = ~n1032 & ~n1157;
  assign n1159 = ~n1099 & n1158;
  assign n1160 = n1038 & n1159;
  assign n1161 = ~n400 & ~n1160;
  assign n1162 = ~n1156 & ~n1161;
  assign n1163 = n1152 & n1162;
  assign n1164 = i_15_ & n277;
  assign n1165 = n72 & n79;
  assign n1166 = ~n469 & ~n1165;
  assign n1167 = ~n1164 & n1166;
  assign n1168 = n175 & n391;
  assign n1169 = ~n1126 & ~n1168;
  assign n1170 = n141 & n1016;
  assign n1171 = i_14_ & n1170;
  assign n1172 = ~n1105 & ~n1171;
  assign n1173 = n1019 & n1172;
  assign n1174 = n1169 & n1173;
  assign n1175 = n1167 & n1174;
  assign n1176 = n358 & ~n1175;
  assign n1177 = n325 & n984;
  assign n1178 = i_8_ & n1177;
  assign n1179 = n606 & ~n1178;
  assign n1180 = ~n523 & ~n1107;
  assign n1181 = ~n1010 & n1180;
  assign n1182 = ~n984 & ~n1040;
  assign n1183 = ~n392 & ~n1113;
  assign n1184 = ~n1011 & n1183;
  assign n1185 = n1182 & n1184;
  assign n1186 = n1181 & n1185;
  assign n1187 = ~n1179 & ~n1186;
  assign n1188 = n153 & n568;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1176 & n1189;
  assign n1191 = n74 & n1016;
  assign n1192 = i_14_ & n1191;
  assign n1193 = n1138 & ~n1192;
  assign n1194 = n358 & ~n1193;
  assign n1195 = n149 & n568;
  assign n1196 = n243 & ~n1015;
  assign n1197 = n243 & n1018;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = ~n1040 & ~n1168;
  assign n1200 = ~n1062 & n1199;
  assign n1201 = n1198 & n1200;
  assign n1202 = n430 & ~n1201;
  assign n1203 = ~n1195 & ~n1202;
  assign n1204 = ~n1194 & n1203;
  assign n1205 = n1190 & n1204;
  assign n1206 = n105 & n114;
  assign n1207 = n340 & n591;
  assign n1208 = ~n1206 & n1207;
  assign n1209 = n1070 & ~n1154;
  assign n1210 = ~n1168 & n1209;
  assign n1211 = n273 & ~n1210;
  assign n1212 = ~n493 & ~n1211;
  assign n1213 = ~n1003 & n1212;
  assign n1214 = ~n1208 & ~n1213;
  assign n1215 = n273 & n1040;
  assign n1216 = i_8_ & ~n387;
  assign n1217 = n1062 & n1216;
  assign n1218 = ~n1215 & ~n1217;
  assign n1219 = n425 & n1062;
  assign n1220 = n309 & ~n1019;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = n1218 & n1221;
  assign n1223 = ~n1154 & n1169;
  assign n1224 = ~n1164 & ~n1165;
  assign n1225 = ~n468 & ~n1036;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1223 & n1226;
  assign n1228 = n1193 & n1227;
  assign n1229 = n309 & ~n1228;
  assign n1230 = ~n243 & ~n273;
  assign n1231 = n310 & n1230;
  assign n1232 = n1035 & ~n1231;
  assign n1233 = ~n1229 & ~n1232;
  assign n1234 = n1222 & n1233;
  assign n1235 = ~n1214 & n1234;
  assign n1236 = n1205 & n1235;
  assign n1237 = n1126 & ~n1153;
  assign n1238 = ~i_8_ & n1168;
  assign n1239 = ~n427 & n1238;
  assign n1240 = ~n313 & ~n1239;
  assign n1241 = n75 & n1067;
  assign n1242 = n1199 & ~n1241;
  assign n1243 = ~n1240 & ~n1242;
  assign n1244 = n82 & n1039;
  assign n1245 = ~n1078 & ~n1244;
  assign n1246 = n898 & ~n1245;
  assign n1247 = n1141 & ~n1244;
  assign n1248 = n275 & ~n1247;
  assign n1249 = n292 & ~n1193;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n1246 & n1250;
  assign n1252 = ~n1243 & n1251;
  assign n1253 = ~n1237 & n1252;
  assign n1254 = ~n464 & ~n1018;
  assign n1255 = ~n1014 & ~n1123;
  assign n1256 = ~n1241 & n1255;
  assign n1257 = n1254 & n1256;
  assign n1258 = n273 & ~n1257;
  assign n1259 = ~n506 & ~n1244;
  assign n1260 = ~i_8_ & n1123;
  assign n1261 = n1259 & ~n1260;
  assign n1262 = n272 & ~n1261;
  assign n1263 = n235 & n1067;
  assign n1264 = n272 & n1263;
  assign n1265 = ~n1262 & ~n1264;
  assign n1266 = ~n1258 & n1265;
  assign n1267 = ~n1078 & n1080;
  assign n1268 = n1247 & n1267;
  assign n1269 = n1155 & n1268;
  assign n1270 = ~n1046 & n1269;
  assign n1271 = n288 & ~n1270;
  assign n1272 = n1266 & ~n1271;
  assign n1273 = n1253 & n1272;
  assign n1274 = n1236 & n1273;
  assign n1275 = n1163 & n1274;
  assign n1276 = ~n1045 & ~n1137;
  assign n1277 = n265 & ~n1276;
  assign n1278 = n696 & n699;
  assign n1279 = n1045 & ~n1278;
  assign n1280 = n428 & n1032;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~n1277 & n1281;
  assign n1283 = n309 & n1123;
  assign n1284 = ~n243 & ~n288;
  assign n1285 = n292 & ~n1101;
  assign n1286 = ~n1008 & ~n1285;
  assign n1287 = ~n1284 & ~n1286;
  assign n1288 = ~n400 & n1165;
  assign n1289 = n307 & ~n1108;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1287 & n1290;
  assign n1292 = ~n1283 & n1291;
  assign n1293 = n1282 & n1292;
  assign n1294 = ~n1014 & ~n1024;
  assign n1295 = n326 & ~n1294;
  assign n1296 = ~n1004 & n1107;
  assign n1297 = ~n703 & n1079;
  assign n1298 = ~n1113 & ~n1165;
  assign n1299 = n1100 & n1298;
  assign n1300 = ~n1137 & n1299;
  assign n1301 = ~n695 & ~n1300;
  assign n1302 = n1106 & n1114;
  assign n1303 = ~n383 & ~n1302;
  assign n1304 = ~n1301 & ~n1303;
  assign n1305 = ~n1297 & n1304;
  assign n1306 = ~n1296 & n1305;
  assign n1307 = ~n1295 & n1306;
  assign n1308 = n1293 & n1307;
  assign n1309 = n1041 & ~n1165;
  assign n1310 = ~n1105 & ~n1113;
  assign n1311 = ~n1107 & n1310;
  assign n1312 = n1309 & n1311;
  assign n1313 = n1019 & n1312;
  assign n1314 = n292 & ~n1313;
  assign n1315 = n1019 & n1268;
  assign n1316 = ~n1137 & n1315;
  assign n1317 = n219 & ~n1316;
  assign n1318 = n517 & n1199;
  assign n1319 = ~n1171 & n1318;
  assign n1320 = n727 & n1319;
  assign n1321 = ~n1317 & n1320;
  assign n1322 = ~n383 & ~n1321;
  assign n1323 = n472 & n1045;
  assign n1324 = ~n1024 & ~n1244;
  assign n1325 = n309 & ~n1324;
  assign n1326 = ~n1323 & ~n1325;
  assign n1327 = ~n1322 & n1326;
  assign n1328 = ~n1314 & n1327;
  assign n1329 = n1308 & n1328;
  assign n1330 = n1275 & n1329;
  assign n1331 = ~n1050 & ~n1157;
  assign n1332 = ~n1054 & n1331;
  assign n1333 = n358 & ~n1332;
  assign n1334 = n1052 & ~n1192;
  assign n1335 = ~n1171 & n1334;
  assign n1336 = n243 & ~n1335;
  assign n1337 = ~n624 & n1171;
  assign n1338 = ~n1078 & ~n1164;
  assign n1339 = ~n1230 & ~n1338;
  assign n1340 = ~n1337 & ~n1339;
  assign n1341 = ~n1336 & n1340;
  assign n1342 = ~n1333 & n1341;
  assign n1343 = ~n606 & n1087;
  assign n1344 = ~n1010 & ~n1244;
  assign n1345 = n430 & ~n1344;
  assign n1346 = ~n1343 & ~n1345;
  assign n1347 = ~n311 & n1060;
  assign n1348 = n1346 & ~n1347;
  assign n1349 = ~n1011 & ~n1050;
  assign n1350 = n425 & ~n1349;
  assign n1351 = ~n307 & ~n472;
  assign n1352 = ~n1011 & ~n1192;
  assign n1353 = n1338 & n1352;
  assign n1354 = ~n1351 & ~n1353;
  assign n1355 = ~n1350 & ~n1354;
  assign n1356 = ~n1010 & ~n1018;
  assign n1357 = n472 & ~n1356;
  assign n1358 = n1355 & ~n1357;
  assign n1359 = n1348 & n1358;
  assign n1360 = n1342 & n1359;
  assign n1361 = ~n1060 & n1332;
  assign n1362 = n292 & ~n1361;
  assign n1363 = ~n326 & ~n898;
  assign n1364 = ~n275 & n1363;
  assign n1365 = n1018 & ~n1364;
  assign n1366 = ~n1362 & ~n1365;
  assign n1367 = ~n358 & ~n380;
  assign n1368 = n1053 & ~n1367;
  assign n1369 = n382 & ~n1334;
  assign n1370 = ~n1054 & ~n1244;
  assign n1371 = n265 & ~n1370;
  assign n1372 = n1140 & ~n1371;
  assign n1373 = ~n265 & ~n292;
  assign n1374 = ~n219 & n1373;
  assign n1375 = ~n1372 & ~n1374;
  assign n1376 = ~n1369 & ~n1375;
  assign n1377 = ~n1368 & n1376;
  assign n1378 = ~n309 & n359;
  assign n1379 = n1139 & ~n1378;
  assign n1380 = n1377 & ~n1379;
  assign n1381 = n1366 & n1380;
  assign n1382 = n313 & n1087;
  assign n1383 = ~n1164 & ~n1382;
  assign n1384 = ~n115 & ~n898;
  assign n1385 = n1373 & n1384;
  assign n1386 = ~n219 & n1385;
  assign n1387 = ~n313 & n1386;
  assign n1388 = ~n1383 & ~n1387;
  assign n1389 = n326 & n1157;
  assign n1390 = n115 & n1011;
  assign n1391 = n243 & n1157;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~n1389 & n1392;
  assign n1394 = ~n265 & n414;
  assign n1395 = n1010 & ~n1394;
  assign n1396 = n1393 & ~n1395;
  assign n1397 = ~n1011 & ~n1053;
  assign n1398 = ~n242 & ~n292;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = n1192 & ~n1384;
  assign n1401 = ~n1018 & ~n1078;
  assign n1402 = ~n314 & ~n1401;
  assign n1403 = ~n1400 & ~n1402;
  assign n1404 = ~n1399 & n1403;
  assign n1405 = n472 & n1244;
  assign n1406 = ~i_8_ & n1050;
  assign n1407 = n1055 & ~n1171;
  assign n1408 = ~n1406 & n1407;
  assign n1409 = n249 & ~n1408;
  assign n1410 = ~n1405 & ~n1409;
  assign n1411 = n1404 & n1410;
  assign n1412 = n1396 & n1411;
  assign n1413 = ~n1388 & n1412;
  assign n1414 = n1381 & n1413;
  assign n1415 = n1360 & n1414;
  assign n1416 = ~n703 & n1139;
  assign n1417 = ~n243 & ~n472;
  assign n1418 = n1054 & ~n1417;
  assign n1419 = ~n359 & n1060;
  assign n1420 = n292 & n1171;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~n1418 & n1421;
  assign n1423 = ~n1416 & n1422;
  assign n1424 = ~n310 & ~n1331;
  assign n1425 = ~n1051 & ~n1424;
  assign n1426 = ~n249 & n343;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1157 & n1353;
  assign n1429 = n275 & ~n1428;
  assign n1430 = ~n1427 & ~n1429;
  assign n1431 = n1423 & n1430;
  assign n1432 = n1415 & n1431;
  assign n1433 = n1330 & n1432;
  assign n1434 = n1136 & n1433;
  assign o_4_ = n164 & ~n1434;
  assign n1436 = n355 & n1415;
  assign n1437 = n952 & n1436;
  assign n1438 = ~i_14_ & n1191;
  assign n1439 = n69 & n235;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = n380 & ~n1440;
  assign n1442 = n69 & n256;
  assign n1443 = i_15_ & n1442;
  assign n1444 = ~n439 & n1443;
  assign n1445 = n69 & n72;
  assign n1446 = n69 & n228;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n387 & ~n1447;
  assign n1449 = ~i_14_ & n1017;
  assign n1450 = n249 & n1449;
  assign n1451 = ~n1448 & ~n1450;
  assign n1452 = ~n1444 & n1451;
  assign n1453 = ~n1441 & n1452;
  assign n1454 = i_8_ & ~n1453;
  assign n1455 = ~i_14_ & ~n68;
  assign n1456 = n142 & n1455;
  assign n1457 = n399 & n1456;
  assign n1458 = n358 & n1438;
  assign n1459 = ~n1018 & ~n1439;
  assign n1460 = ~n441 & ~n1459;
  assign n1461 = ~n1458 & ~n1460;
  assign n1462 = ~n1457 & n1461;
  assign n1463 = ~n1454 & n1462;
  assign n1464 = n69 & n175;
  assign n1465 = ~i_14_ & n1170;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1017 & n1466;
  assign n1468 = ~n1439 & n1467;
  assign n1469 = n243 & ~n1468;
  assign n1470 = ~n624 & n1465;
  assign n1471 = ~n606 & n1446;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n273 & n1351;
  assign n1474 = n1443 & ~n1473;
  assign n1475 = ~n1192 & n1344;
  assign n1476 = n1466 & n1475;
  assign n1477 = n273 & ~n1476;
  assign n1478 = ~n1351 & n1464;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1474 & n1479;
  assign n1481 = n1472 & n1480;
  assign n1482 = ~n1469 & n1481;
  assign n1483 = n1463 & n1482;
  assign n1484 = ~n183 & ~n1051;
  assign n1485 = ~n481 & ~n1050;
  assign n1486 = n232 & n1485;
  assign n1487 = n1484 & n1486;
  assign n1488 = ~n236 & ~n1054;
  assign n1489 = ~n800 & n1488;
  assign n1490 = ~n494 & n1489;
  assign n1491 = n1487 & n1490;
  assign n1492 = n898 & ~n1491;
  assign n1493 = ~n1078 & n1370;
  assign n1494 = n837 & n1493;
  assign n1495 = n380 & ~n1494;
  assign n1496 = n379 & n474;
  assign n1497 = n86 & n1039;
  assign n1498 = i_8_ & n143;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = n272 & ~n1499;
  assign n1501 = ~n1496 & ~n1500;
  assign n1502 = ~n1495 & n1501;
  assign n1503 = n69 & n252;
  assign n1504 = ~n700 & n1503;
  assign n1505 = ~n245 & ~n1157;
  assign n1506 = n454 & n1505;
  assign n1507 = ~n699 & ~n1506;
  assign n1508 = ~n1504 & ~n1507;
  assign n1509 = n898 & ~n1259;
  assign n1510 = n472 & n1503;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = n179 & n265;
  assign n1513 = n1511 & ~n1512;
  assign n1514 = n1508 & n1513;
  assign n1515 = n69 & n294;
  assign n1516 = ~n393 & ~n1515;
  assign n1517 = n459 & n1516;
  assign n1518 = n249 & ~n1517;
  assign n1519 = ~n313 & ~n379;
  assign n1520 = ~n226 & ~n1139;
  assign n1521 = ~n258 & ~n1053;
  assign n1522 = n1520 & n1521;
  assign n1523 = n837 & n1522;
  assign n1524 = ~n1519 & ~n1523;
  assign n1525 = ~n1518 & ~n1524;
  assign n1526 = n115 & n183;
  assign n1527 = n1525 & ~n1526;
  assign n1528 = n1514 & n1527;
  assign n1529 = n1502 & n1528;
  assign n1530 = ~n1492 & n1529;
  assign n1531 = n1483 & n1530;
  assign n1532 = n69 & n233;
  assign n1533 = ~n169 & ~n1515;
  assign n1534 = n265 & ~n1533;
  assign n1535 = ~n1532 & ~n1534;
  assign n1536 = ~n1385 & ~n1535;
  assign n1537 = ~i_15_ & n1442;
  assign n1538 = n313 & n1537;
  assign n1539 = ~n1536 & ~n1538;
  assign n1540 = ~n169 & ~n181;
  assign n1541 = n115 & ~n1540;
  assign n1542 = n69 & n254;
  assign n1543 = ~n174 & ~n1542;
  assign n1544 = ~n181 & n1543;
  assign n1545 = ~n753 & ~n1544;
  assign n1546 = ~n1541 & ~n1545;
  assign n1547 = n1539 & n1546;
  assign n1548 = ~n169 & ~n1503;
  assign n1549 = n1543 & n1548;
  assign n1550 = n313 & ~n1549;
  assign n1551 = ~n177 & ~n414;
  assign n1552 = n86 & n235;
  assign n1553 = n86 & n228;
  assign n1554 = ~n1532 & ~n1553;
  assign n1555 = ~n1552 & n1554;
  assign n1556 = ~n180 & ~n1537;
  assign n1557 = n170 & n1556;
  assign n1558 = n1555 & n1557;
  assign n1559 = n219 & ~n1558;
  assign n1560 = ~n1551 & ~n1559;
  assign n1561 = ~n1550 & n1560;
  assign n1562 = n1547 & n1561;
  assign n1563 = n86 & n463;
  assign n1564 = ~n1542 & ~n1563;
  assign n1565 = ~n1503 & ~n1552;
  assign n1566 = ~n1553 & n1565;
  assign n1567 = n1564 & n1566;
  assign n1568 = ~n143 & ~n1515;
  assign n1569 = n1567 & n1568;
  assign n1570 = ~n144 & n1569;
  assign n1571 = n292 & ~n1570;
  assign n1572 = ~n168 & ~n1552;
  assign n1573 = ~n1553 & n1572;
  assign n1574 = ~n1563 & n1573;
  assign n1575 = ~n180 & n1574;
  assign n1576 = n265 & ~n1575;
  assign n1577 = ~n176 & ~n1497;
  assign n1578 = ~n358 & n381;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n292 & ~n307;
  assign n1581 = n307 & n1552;
  assign n1582 = ~n1497 & ~n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584 = ~n1579 & ~n1583;
  assign n1585 = ~n1576 & n1584;
  assign n1586 = ~n911 & n1537;
  assign n1587 = n170 & n182;
  assign n1588 = n1567 & n1587;
  assign n1589 = n275 & ~n1588;
  assign n1590 = ~n1586 & ~n1589;
  assign n1591 = n1585 & n1590;
  assign n1592 = ~n1571 & n1591;
  assign n1593 = n1562 & n1592;
  assign n1594 = ~n266 & ~n1087;
  assign n1595 = ~n167 & n1594;
  assign n1596 = n1489 & n1595;
  assign n1597 = ~n1417 & ~n1596;
  assign n1598 = n183 & n243;
  assign n1599 = ~n220 & n1484;
  assign n1600 = ~n234 & n1485;
  assign n1601 = n1599 & n1600;
  assign n1602 = n309 & ~n1601;
  assign n1603 = ~n1598 & ~n1602;
  assign n1604 = ~n1597 & n1603;
  assign n1605 = ~n494 & n1505;
  assign n1606 = n1487 & n1605;
  assign n1607 = ~n1351 & ~n1606;
  assign n1608 = ~n595 & ~n1060;
  assign n1609 = ~n293 & n1608;
  assign n1610 = n1523 & n1609;
  assign n1611 = n273 & ~n1610;
  assign n1612 = n1599 & n1609;
  assign n1613 = n358 & ~n1612;
  assign n1614 = n249 & n1087;
  assign n1615 = i_8_ & n1614;
  assign n1616 = ~n1613 & ~n1615;
  assign n1617 = ~n1611 & n1616;
  assign n1618 = ~n1607 & n1617;
  assign n1619 = n1604 & n1618;
  assign n1620 = n1593 & n1619;
  assign n1621 = n1531 & n1620;
  assign n1622 = n1437 & n1621;
  assign n1623 = n273 & ~n1548;
  assign n1624 = n243 & ~n1543;
  assign n1625 = n399 & n1515;
  assign n1626 = ~n440 & ~n1625;
  assign n1627 = ~n1568 & ~n1626;
  assign n1628 = ~n1624 & ~n1627;
  assign n1629 = ~n1623 & n1628;
  assign n1630 = ~n170 & ~n606;
  assign n1631 = ~n174 & n1554;
  assign n1632 = ~n143 & n1631;
  assign n1633 = ~n310 & ~n1632;
  assign n1634 = ~n1630 & ~n1633;
  assign n1635 = ~n1515 & ~n1532;
  assign n1636 = n1216 & ~n1635;
  assign n1637 = ~n441 & n1542;
  assign n1638 = ~n168 & n1548;
  assign n1639 = n430 & ~n1638;
  assign n1640 = ~n1637 & ~n1639;
  assign n1641 = ~n1636 & n1640;
  assign n1642 = n1634 & n1641;
  assign n1643 = n1629 & n1642;
  assign n1644 = n358 & ~n1567;
  assign n1645 = n174 & ~n573;
  assign n1646 = n243 & ~n1555;
  assign n1647 = ~n1542 & ~n1552;
  assign n1648 = n309 & ~n1647;
  assign n1649 = ~n1646 & ~n1648;
  assign n1650 = ~n1645 & n1649;
  assign n1651 = ~n1644 & n1650;
  assign n1652 = n1643 & n1651;
  assign n1653 = n695 & n824;
  assign n1654 = n1438 & ~n1653;
  assign n1655 = ~n754 & n1446;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = n1652 & n1656;
  assign n1658 = ~n217 & ~n430;
  assign n1659 = n1563 & ~n1658;
  assign n1660 = n385 & ~n1456;
  assign n1661 = ~n383 & ~n1660;
  assign n1662 = ~n1659 & ~n1661;
  assign n1663 = ~n1063 & n1443;
  assign n1664 = ~n1244 & ~n1497;
  assign n1665 = n275 & ~n1664;
  assign n1666 = ~n1449 & ~n1665;
  assign n1667 = ~n273 & n414;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~n1663 & ~n1668;
  assign n1670 = n243 & n255;
  assign n1671 = n1012 & ~n1192;
  assign n1672 = n358 & ~n1671;
  assign n1673 = ~n1670 & ~n1672;
  assign n1674 = ~n1011 & ~n1171;
  assign n1675 = n273 & ~n1674;
  assign n1676 = n292 & n1442;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n1673 & n1677;
  assign n1679 = n1669 & n1678;
  assign n1680 = n1662 & n1679;
  assign n1681 = ~n180 & ~n1438;
  assign n1682 = n317 & n1577;
  assign n1683 = n1573 & n1682;
  assign n1684 = n1681 & n1683;
  assign n1685 = ~n1449 & n1684;
  assign n1686 = n379 & ~n1685;
  assign n1687 = n1012 & ~n1515;
  assign n1688 = ~n699 & ~n1687;
  assign n1689 = ~n1464 & ~n1688;
  assign n1690 = ~n1064 & ~n1689;
  assign n1691 = ~n1686 & ~n1690;
  assign n1692 = n1245 & ~n1439;
  assign n1693 = n288 & ~n1692;
  assign n1694 = ~n115 & ~n272;
  assign n1695 = n228 & n1455;
  assign n1696 = n176 & n272;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~n1694 & ~n1697;
  assign n1699 = ~n1693 & ~n1698;
  assign n1700 = ~n314 & n1438;
  assign n1701 = n72 & n1455;
  assign n1702 = n273 & n1701;
  assign n1703 = n463 & n1455;
  assign n1704 = n313 & n1703;
  assign n1705 = ~n1702 & ~n1704;
  assign n1706 = ~n1700 & n1705;
  assign n1707 = n1699 & n1706;
  assign n1708 = i_8_ & n1164;
  assign n1709 = ~n1018 & ~n1708;
  assign n1710 = n380 & ~n1709;
  assign n1711 = ~n1449 & ~n1710;
  assign n1712 = ~n265 & n1367;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = n1707 & ~n1713;
  assign n1715 = n273 & n1438;
  assign n1716 = n115 & n1455;
  assign n1717 = ~n76 & n1716;
  assign n1718 = ~n1715 & ~n1717;
  assign n1719 = ~n1449 & ~n1465;
  assign n1720 = ~n1439 & n1719;
  assign n1721 = n313 & ~n1720;
  assign n1722 = ~n292 & ~n309;
  assign n1723 = n1192 & ~n1722;
  assign n1724 = ~n1721 & ~n1723;
  assign n1725 = n1718 & n1724;
  assign n1726 = n1714 & n1725;
  assign n1727 = n1691 & n1726;
  assign n1728 = n1680 & n1727;
  assign n1729 = n181 & ~n311;
  assign n1730 = n176 & n307;
  assign n1731 = n174 & n273;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1729 & n1732;
  assign n1734 = n310 & ~n440;
  assign n1735 = ~n1556 & ~n1734;
  assign n1736 = ~n181 & ~n1537;
  assign n1737 = n1216 & ~n1736;
  assign n1738 = n472 & n1542;
  assign n1739 = ~n1737 & ~n1738;
  assign n1740 = ~n1735 & n1739;
  assign n1741 = n1733 & n1740;
  assign n1742 = ~n1004 & n1439;
  assign n1743 = n383 & n427;
  assign n1744 = n1465 & ~n1743;
  assign n1745 = ~n1742 & ~n1744;
  assign n1746 = ~n180 & n1488;
  assign n1747 = ~n231 & ~n1051;
  assign n1748 = i_8_ & n1703;
  assign n1749 = ~n1552 & ~n1748;
  assign n1750 = n1747 & n1749;
  assign n1751 = n1746 & n1750;
  assign n1752 = n272 & ~n1751;
  assign n1753 = ~n1443 & ~n1456;
  assign n1754 = ~n168 & ~n1445;
  assign n1755 = n1753 & n1754;
  assign n1756 = ~n181 & ~n1515;
  assign n1757 = n69 & n153;
  assign n1758 = ~n1011 & ~n1757;
  assign n1759 = n1756 & n1758;
  assign n1760 = n1755 & n1759;
  assign n1761 = n1475 & n1760;
  assign n1762 = n313 & ~n1761;
  assign n1763 = ~n1752 & ~n1762;
  assign n1764 = n1745 & n1763;
  assign n1765 = n1741 & n1764;
  assign n1766 = n1728 & n1765;
  assign n1767 = ~n358 & n1153;
  assign n1768 = n1171 & ~n1767;
  assign n1769 = n700 & n865;
  assign n1770 = n1445 & ~n1769;
  assign n1771 = ~n1768 & ~n1770;
  assign n1772 = n449 & n1771;
  assign n1773 = n1766 & n1772;
  assign n1774 = n1657 & n1773;
  assign n1775 = ~n507 & ~n1078;
  assign n1776 = n1595 & n1775;
  assign n1777 = n898 & ~n1776;
  assign n1778 = ~n218 & ~n242;
  assign n1779 = ~n380 & n1778;
  assign n1780 = n457 & ~n1779;
  assign n1781 = n167 & ~n847;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = n169 & n379;
  assign n1784 = ~n179 & n1520;
  assign n1785 = n430 & ~n1784;
  assign n1786 = ~n167 & ~n469;
  assign n1787 = n249 & ~n1786;
  assign n1788 = ~n1785 & ~n1787;
  assign n1789 = ~n1783 & n1788;
  assign n1790 = n1782 & n1789;
  assign n1791 = ~n1777 & n1790;
  assign n1792 = ~n255 & ~n494;
  assign n1793 = ~n1157 & n1792;
  assign n1794 = n275 & ~n1793;
  assign n1795 = ~n231 & n1484;
  assign n1796 = ~n717 & ~n1456;
  assign n1797 = n578 & n1796;
  assign n1798 = n1795 & n1797;
  assign n1799 = n1353 & n1798;
  assign n1800 = ~n474 & ~n1532;
  assign n1801 = n1594 & n1800;
  assign n1802 = n954 & n1801;
  assign n1803 = n1799 & n1802;
  assign n1804 = n275 & ~n1803;
  assign n1805 = ~n1794 & ~n1804;
  assign n1806 = n219 & ~n815;
  assign n1807 = n338 & n800;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = n181 & n358;
  assign n1810 = ~n504 & ~n1171;
  assign n1811 = n292 & ~n1810;
  assign n1812 = ~n1809 & ~n1811;
  assign n1813 = n482 & ~n798;
  assign n1814 = n242 & ~n1813;
  assign n1815 = n1812 & ~n1814;
  assign n1816 = n1808 & n1815;
  assign n1817 = n288 & ~n1709;
  assign n1818 = n292 & ~n1540;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = n358 & n1532;
  assign n1821 = ~n958 & ~n1820;
  assign n1822 = ~n467 & n1821;
  assign n1823 = n1819 & n1822;
  assign n1824 = ~n413 & ~n492;
  assign n1825 = n288 & ~n1824;
  assign n1826 = n292 & ~n1599;
  assign n1827 = n265 & ~n1605;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1825 & n1828;
  assign n1830 = n1823 & n1829;
  assign n1831 = n1816 & n1830;
  assign n1832 = n1805 & n1831;
  assign n1833 = n1791 & n1832;
  assign n1834 = n853 & n1833;
  assign n1835 = n1774 & n1834;
  assign n1836 = n797 & n1835;
  assign n1837 = n1622 & n1836;
  assign o_5_ = n164 & ~n1837;
  assign n1839 = ~n383 & n1503;
  assign n1840 = ~n143 & n1635;
  assign n1841 = n275 & ~n1840;
  assign n1842 = ~n1818 & ~n1841;
  assign n1843 = ~n1839 & n1842;
  assign n1844 = n1593 & n1843;
  assign n1845 = n253 & n358;
  assign n1846 = ~n309 & ~n1845;
  assign n1847 = ~n384 & ~n1846;
  assign n1848 = n1483 & ~n1847;
  assign n1849 = n1844 & n1848;
  assign n1850 = ~n383 & ~n1505;
  assign n1851 = ~n1087 & n1522;
  assign n1852 = n1052 & n1851;
  assign n1853 = n268 & n1852;
  assign n1854 = n379 & ~n1853;
  assign n1855 = n295 & ~n1153;
  assign n1856 = ~n1854 & ~n1855;
  assign n1857 = ~n210 & n1856;
  assign n1858 = ~n1850 & n1857;
  assign n1859 = n61 & n96;
  assign n1860 = n58 & n1859;
  assign n1861 = n217 & n255;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = n1039 & n1455;
  assign n1864 = i_8_ & n1456;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = n272 & ~n1865;
  assign n1867 = ~n159 & ~n1866;
  assign n1868 = ~n253 & ~n255;
  assign n1869 = n273 & ~n1868;
  assign n1870 = ~n1783 & ~n1869;
  assign n1871 = ~n1817 & n1870;
  assign n1872 = n1867 & n1871;
  assign n1873 = n1862 & n1872;
  assign n1874 = n309 & n1503;
  assign n1875 = n307 & n1515;
  assign n1876 = ~n1820 & ~n1875;
  assign n1877 = ~n1874 & n1876;
  assign n1878 = ~i_5_ & n204;
  assign n1879 = n1877 & ~n1878;
  assign n1880 = ~n694 & n1087;
  assign n1881 = ~n479 & ~n1880;
  assign n1882 = ~n699 & ~n1493;
  assign n1883 = ~n115 & ~n243;
  assign n1884 = n234 & ~n1883;
  assign n1885 = ~n1882 & ~n1884;
  assign n1886 = n1881 & n1885;
  assign n1887 = ~n1809 & n1886;
  assign n1888 = n1879 & n1887;
  assign n1889 = n1873 & n1888;
  assign n1890 = n1858 & n1889;
  assign n1891 = n378 & n1890;
  assign n1892 = n1774 & n1891;
  assign n1893 = n1849 & n1892;
  assign n1894 = n1432 & n1893;
  assign o_8_ = n164 & ~n1894;
  assign n1896 = n1117 & n1877;
  assign n1897 = n128 & n273;
  assign n1898 = ~n180 & ~n596;
  assign n1899 = ~i_14_ & n254;
  assign n1900 = i_12_ & n1899;
  assign n1901 = ~n1563 & ~n1900;
  assign n1902 = n1898 & n1901;
  assign n1903 = n472 & ~n1902;
  assign n1904 = n86 & n290;
  assign n1905 = n1216 & n1904;
  assign n1906 = ~n1903 & ~n1905;
  assign n1907 = ~n1897 & n1906;
  assign n1908 = ~n607 & ~n1032;
  assign n1909 = ~n1497 & n1908;
  assign n1910 = ~n176 & ~n1008;
  assign n1911 = ~n597 & n1910;
  assign n1912 = n1909 & n1911;
  assign n1913 = n273 & ~n1912;
  assign n1914 = ~n1008 & ~n1904;
  assign n1915 = n307 & ~n1914;
  assign n1916 = ~n1809 & ~n1915;
  assign n1917 = ~n1913 & n1916;
  assign n1918 = ~n128 & ~n1045;
  assign n1919 = ~n573 & ~n1918;
  assign n1920 = n1917 & ~n1919;
  assign n1921 = n1907 & n1920;
  assign n1922 = n1741 & n1921;
  assign n1923 = n78 & n1899;
  assign n1924 = ~n311 & n1923;
  assign n1925 = n1922 & ~n1924;
  assign n1926 = n1896 & n1925;
  assign n1927 = ~n439 & n1904;
  assign n1928 = ~n1118 & ~n1927;
  assign n1929 = ~n602 & ~n1036;
  assign n1930 = ~n1552 & n1929;
  assign n1931 = ~n586 & ~n1099;
  assign n1932 = ~n168 & n1931;
  assign n1933 = n1930 & n1932;
  assign n1934 = ~n387 & ~n1933;
  assign n1935 = n1928 & ~n1934;
  assign n1936 = i_8_ & ~n1935;
  assign n1937 = n358 & n1923;
  assign n1938 = n86 & n172;
  assign n1939 = n472 & n1938;
  assign n1940 = ~n1937 & ~n1939;
  assign n1941 = n309 & ~n814;
  assign n1942 = ~n800 & ~n1046;
  assign n1943 = n358 & ~n1942;
  assign n1944 = n86 & n252;
  assign n1945 = n273 & n1944;
  assign n1946 = ~n1943 & ~n1945;
  assign n1947 = ~n1941 & n1946;
  assign n1948 = n1940 & n1947;
  assign n1949 = n86 & n294;
  assign n1950 = ~n1208 & n1949;
  assign n1951 = n1948 & ~n1950;
  assign n1952 = ~n1936 & n1951;
  assign n1953 = n86 & n233;
  assign n1954 = ~n88 & ~n1953;
  assign n1955 = ~n606 & ~n1954;
  assign n1956 = ~n273 & ~n1955;
  assign n1957 = ~n609 & ~n1046;
  assign n1958 = ~n143 & n1957;
  assign n1959 = ~n1047 & ~n1553;
  assign n1960 = n1958 & n1959;
  assign n1961 = n1954 & n1960;
  assign n1962 = ~n705 & n1961;
  assign n1963 = ~n1956 & ~n1962;
  assign n1964 = ~n430 & n606;
  assign n1965 = n1944 & ~n1964;
  assign n1966 = n1901 & ~n1938;
  assign n1967 = ~n307 & n1230;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n1965 & ~n1968;
  assign n1970 = ~n1963 & n1969;
  assign n1971 = n1952 & n1970;
  assign n1972 = n1652 & n1971;
  assign n1973 = n1926 & n1972;
  assign n1974 = n272 & ~n1311;
  assign n1975 = ~n381 & n1032;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~n128 & n1954;
  assign n1978 = ~n696 & ~n1977;
  assign n1979 = ~n699 & n1938;
  assign n1980 = ~n313 & n699;
  assign n1981 = n128 & ~n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1983 = ~n1978 & n1982;
  assign n1984 = ~n1045 & n1898;
  assign n1985 = ~n494 & n1984;
  assign n1986 = n273 & ~n1985;
  assign n1987 = n472 & ~n1909;
  assign n1988 = n481 & ~n1883;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1986 & n1989;
  assign n1991 = n1983 & n1990;
  assign n1992 = n1976 & n1991;
  assign n1993 = n623 & n1992;
  assign n1994 = ~n399 & n1153;
  assign n1995 = n143 & ~n1994;
  assign n1996 = ~n383 & ~n825;
  assign n1997 = n307 & n609;
  assign n1998 = ~n595 & ~n1938;
  assign n1999 = n313 & ~n1998;
  assign n2000 = ~n1997 & ~n1999;
  assign n2001 = ~n542 & n1137;
  assign n2002 = n273 & n800;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = n243 & ~n1255;
  assign n2005 = n115 & n144;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = n2003 & n2006;
  assign n2008 = n2000 & n2007;
  assign n2009 = ~n338 & ~n358;
  assign n2010 = n1938 & ~n2009;
  assign n2011 = n2008 & ~n2010;
  assign n2012 = ~n1996 & n2011;
  assign n2013 = ~n1995 & n2012;
  assign n2014 = ~n1944 & ~n1949;
  assign n2015 = ~n1005 & ~n2014;
  assign n2016 = ~n405 & n1553;
  assign n2017 = ~n340 & n494;
  assign n2018 = n1143 & n1298;
  assign n2019 = ~n1107 & n2018;
  assign n2020 = n309 & ~n2019;
  assign n2021 = ~n2017 & ~n2020;
  assign n2022 = ~n2016 & n2021;
  assign n2023 = n1572 & n1898;
  assign n2024 = ~n610 & n2023;
  assign n2025 = n898 & ~n2024;
  assign n2026 = n2022 & ~n2025;
  assign n2027 = ~n2015 & n2026;
  assign n2028 = n2013 & n2027;
  assign n2029 = n1993 & n2028;
  assign n2030 = n1973 & n2029;
  assign n2031 = ~n1515 & n1957;
  assign n2032 = ~n181 & n1984;
  assign n2033 = ~n1047 & n1800;
  assign n2034 = n1901 & n1909;
  assign n2035 = n2033 & n2034;
  assign n2036 = n1933 & n2035;
  assign n2037 = n2032 & n2036;
  assign n2038 = n2031 & n2037;
  assign n2039 = n313 & ~n2038;
  assign n2040 = n898 & ~n1909;
  assign n2041 = n329 & n899;
  assign n2042 = n1904 & ~n2041;
  assign n2043 = ~n2040 & ~n2042;
  assign n2044 = ~n1153 & ~n1954;
  assign n2045 = n338 & ~n1038;
  assign n2046 = n1037 & ~n1563;
  assign n2047 = ~n1515 & n2046;
  assign n2048 = ~n699 & ~n2047;
  assign n2049 = n1106 & ~n1904;
  assign n2050 = n275 & ~n2049;
  assign n2051 = ~n1519 & ~n1911;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = ~n2048 & n2052;
  assign n2054 = ~n2045 & n2053;
  assign n2055 = ~n2044 & n2054;
  assign n2056 = n2043 & n2055;
  assign n2057 = ~n2039 & n2056;
  assign n2058 = ~n272 & n1743;
  assign n2059 = ~n1255 & ~n2058;
  assign n2060 = ~n288 & n1004;
  assign n2061 = n1079 & ~n2060;
  assign n2062 = ~n2059 & ~n2061;
  assign n2063 = ~n1537 & n1908;
  assign n2064 = ~n1046 & ~n1938;
  assign n2065 = n2063 & n2064;
  assign n2066 = n292 & ~n2065;
  assign n2067 = n400 & n414;
  assign n2068 = n1923 & ~n2067;
  assign n2069 = ~n80 & n1311;
  assign n2070 = n288 & ~n2069;
  assign n2071 = ~n2068 & ~n2070;
  assign n2072 = ~n2066 & n2071;
  assign n2073 = n2062 & n2072;
  assign n2074 = n2057 & n2073;
  assign n2075 = n1308 & n2074;
  assign n2076 = ~n602 & n1931;
  assign n2077 = ~n700 & ~n2076;
  assign n2078 = ~i_8_ & n128;
  assign n2079 = n242 & n2078;
  assign n2080 = n380 & ~n1914;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = ~n2077 & n2081;
  assign n2083 = n275 & ~n1909;
  assign n2084 = ~n1783 & ~n2083;
  assign n2085 = ~n1496 & n2084;
  assign n2086 = n2082 & n2085;
  assign n2087 = n1844 & n2086;
  assign n2088 = n2075 & n2087;
  assign n2089 = n882 & n2088;
  assign n2090 = n2030 & n2089;
  assign o_9_ = n164 & ~n2090;
  assign n2092 = ~n278 & n1166;
  assign n2093 = n1784 & n1911;
  assign n2094 = ~n465 & ~n1164;
  assign n2095 = ~n174 & n2094;
  assign n2096 = n2093 & n2095;
  assign n2097 = n2092 & n2096;
  assign n2098 = n273 & ~n2097;
  assign n2099 = n1166 & n2094;
  assign n2100 = ~n278 & n1595;
  assign n2101 = n1932 & n2100;
  assign n2102 = n2099 & n2101;
  assign n2103 = ~n169 & n2102;
  assign n2104 = n313 & ~n2103;
  assign n2105 = ~n2098 & ~n2104;
  assign n2106 = n1796 & n2031;
  assign n2107 = ~n1241 & n2106;
  assign n2108 = n313 & ~n2107;
  assign n2109 = ~n279 & n1080;
  assign n2110 = n273 & ~n2109;
  assign n2111 = ~n1464 & ~n1938;
  assign n2112 = i_8_ & ~n1775;
  assign n2113 = n2111 & ~n2112;
  assign n2114 = n272 & ~n2113;
  assign n2115 = ~n2110 & ~n2114;
  assign n2116 = ~n2108 & n2115;
  assign n2117 = n272 & n1068;
  assign n2118 = n273 & n295;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~n451 & ~n1168;
  assign n2121 = n273 & ~n2120;
  assign n2122 = n127 & n662;
  assign n2123 = ~n1923 & ~n2122;
  assign n2124 = n313 & ~n2123;
  assign n2125 = ~n2121 & ~n2124;
  assign n2126 = ~n548 & n2125;
  assign n2127 = n107 & n391;
  assign n2128 = ~n635 & ~n2127;
  assign n2129 = ~n1014 & ~n1018;
  assign n2130 = n68 & n254;
  assign n2131 = ~n464 & ~n1449;
  assign n2132 = ~n2130 & n2131;
  assign n2133 = n2129 & n2132;
  assign n2134 = n2128 & n2133;
  assign n2135 = n313 & ~n2134;
  assign n2136 = n2126 & ~n2135;
  assign n2137 = n2119 & n2136;
  assign n2138 = n2116 & n2137;
  assign n2139 = ~n1695 & n2033;
  assign n2140 = ~i_8_ & ~n2139;
  assign n2141 = i_8_ & ~n1800;
  assign n2142 = ~n229 & ~n1050;
  assign n2143 = n1959 & n2142;
  assign n2144 = i_8_ & ~n2143;
  assign n2145 = ~n2141 & ~n2144;
  assign n2146 = ~n1069 & n2145;
  assign n2147 = ~n663 & n2146;
  assign n2148 = ~n2140 & n2147;
  assign n2149 = n272 & ~n2148;
  assign n2150 = n2138 & ~n2149;
  assign n2151 = n2105 & n2150;
  assign n2152 = ~n453 & ~n1126;
  assign n2153 = ~n1438 & n2152;
  assign n2154 = ~i_8_ & ~n2153;
  assign n2155 = ~n556 & ~n984;
  assign n2156 = ~n1446 & ~n1953;
  assign n2157 = n2155 & n2156;
  assign n2158 = ~n2154 & n2157;
  assign n2159 = ~n2078 & n2158;
  assign n2160 = ~n1465 & ~n1949;
  assign n2161 = ~n635 & ~n1449;
  assign n2162 = ~n1923 & n2161;
  assign n2163 = ~n1062 & n2162;
  assign n2164 = n2160 & n2163;
  assign n2165 = i_8_ & ~n2164;
  assign n2166 = n2159 & ~n2165;
  assign n2167 = n272 & ~n2166;
  assign n2168 = n273 & ~n1595;
  assign n2169 = n1605 & n1901;
  assign n2170 = n313 & ~n2169;
  assign n2171 = ~n2168 & ~n2170;
  assign n2172 = ~n2167 & n2171;
  assign n2173 = n2151 & n2172;
  assign n2174 = ~n640 & ~n777;
  assign n2175 = n991 & n2174;
  assign n2176 = n743 & n996;
  assign n2177 = n2175 & n2176;
  assign n2178 = ~n78 & n1899;
  assign n2179 = n2031 & ~n2178;
  assign n2180 = ~n183 & n2179;
  assign n2181 = n273 & ~n2180;
  assign n2182 = ~n764 & ~n2181;
  assign n2183 = ~n1032 & ~n1045;
  assign n2184 = n1929 & n2183;
  assign n2185 = ~n181 & n2184;
  assign n2186 = n272 & ~n2185;
  assign n2187 = n313 & n800;
  assign n2188 = n273 & n1537;
  assign n2189 = n272 & n1503;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = ~n2187 & n2190;
  assign n2192 = ~n2186 & n2191;
  assign n2193 = n350 & n937;
  assign n2194 = n2192 & n2193;
  assign n2195 = n1266 & ~n1752;
  assign n2196 = ~n710 & ~n1866;
  assign n2197 = ~n1538 & n2196;
  assign n2198 = ~n857 & n2197;
  assign n2199 = n2195 & n2198;
  assign n2200 = n2194 & n2199;
  assign n2201 = n2182 & n2200;
  assign n2202 = n273 & ~n2153;
  assign n2203 = n2201 & ~n2202;
  assign n2204 = n2177 & n2203;
  assign n2205 = n273 & ~n1932;
  assign n2206 = n1911 & n2109;
  assign n2207 = n1784 & n2206;
  assign n2208 = n1775 & n2207;
  assign n2209 = n313 & ~n2208;
  assign n2210 = ~n558 & ~n1439;
  assign n2211 = ~n1035 & n2210;
  assign n2212 = ~n1443 & ~n1904;
  assign n2213 = n2211 & n2212;
  assign n2214 = n273 & ~n2213;
  assign n2215 = ~n1944 & n2211;
  assign n2216 = n313 & ~n2215;
  assign n2217 = ~n2214 & ~n2216;
  assign n2218 = ~n570 & ~n1040;
  assign n2219 = ~n169 & n2218;
  assign n2220 = n273 & ~n2219;
  assign n2221 = n174 & n313;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = n2217 & n2222;
  assign n2224 = ~n2209 & n2223;
  assign n2225 = ~n457 & ~n1445;
  assign n2226 = ~n88 & ~n1154;
  assign n2227 = n2225 & n2226;
  assign n2228 = ~n1238 & n2227;
  assign n2229 = n272 & ~n2228;
  assign n2230 = n313 & ~n2212;
  assign n2231 = n313 & n451;
  assign n2232 = n313 & ~n2218;
  assign n2233 = ~n1945 & ~n2232;
  assign n2234 = ~n2231 & n2233;
  assign n2235 = ~n2230 & n2234;
  assign n2236 = ~n2229 & n2235;
  assign n2237 = n2224 & n2236;
  assign n2238 = ~n2205 & n2237;
  assign n2239 = ~n413 & ~n1003;
  assign n2240 = n272 & ~n2239;
  assign n2241 = n313 & ~n2160;
  assign n2242 = ~n1897 & ~n2241;
  assign n2243 = ~n2240 & n2242;
  assign n2244 = n2238 & n2243;
  assign n2245 = n2204 & n2244;
  assign n2246 = n2173 & n2245;
  assign o_10_ = n164 & ~n2246;
  assign n2248 = ~n474 & ~n509;
  assign n2249 = ~n1011 & n2248;
  assign n2250 = n1554 & n2142;
  assign n2251 = n2249 & n2250;
  assign n2252 = ~n663 & n2251;
  assign n2253 = n115 & ~n2252;
  assign n2254 = ~n277 & ~n456;
  assign n2255 = ~n169 & ~n1701;
  assign n2256 = n2254 & n2255;
  assign n2257 = n115 & ~n2256;
  assign n2258 = ~n942 & ~n2257;
  assign n2259 = ~n518 & ~n1457;
  assign n2260 = n2258 & n2259;
  assign n2261 = ~n2253 & n2260;
  assign n2262 = n2160 & n2239;
  assign n2263 = n1172 & n2262;
  assign n2264 = n2031 & n2263;
  assign n2265 = ~n595 & n2264;
  assign n2266 = ~n295 & n2265;
  assign n2267 = n399 & ~n2266;
  assign n2268 = ~n1445 & n1918;
  assign n2269 = n2226 & n2268;
  assign n2270 = n1299 & n2157;
  assign n2271 = n2269 & n2270;
  assign n2272 = ~n167 & n2271;
  assign n2273 = n115 & ~n2272;
  assign n2274 = n182 & n1138;
  assign n2275 = ~n231 & n1599;
  assign n2276 = ~n596 & n2275;
  assign n2277 = ~n510 & ~n1192;
  assign n2278 = n2153 & n2277;
  assign n2279 = n2276 & n2278;
  assign n2280 = n2274 & n2279;
  assign n2281 = n115 & ~n2280;
  assign n2282 = ~n2273 & ~n2281;
  assign n2283 = ~n2267 & n2282;
  assign o_11_ = ~n2261 | ~n2283;
  assign n2285 = ~n556 & ~n1446;
  assign n2286 = ~n1542 & n2169;
  assign n2287 = n2285 & n2286;
  assign n2288 = i_8_ & ~n2287;
  assign n2289 = n1184 & ~n1532;
  assign n2290 = n482 & n2248;
  assign n2291 = n2143 & n2290;
  assign n2292 = ~n464 & n1019;
  assign n2293 = ~n255 & n2292;
  assign n2294 = ~i_8_ & ~n2293;
  assign n2295 = n2291 & ~n2294;
  assign n2296 = n2289 & n2295;
  assign n2297 = ~n2288 & n2296;
  assign n2298 = n379 & ~n2297;
  assign n2299 = ~n767 & n1488;
  assign n2300 = n1180 & n2299;
  assign n2301 = n557 & n1344;
  assign n2302 = ~n1442 & ~n1904;
  assign n2303 = ~n1944 & n2302;
  assign n2304 = n1930 & n2303;
  assign n2305 = n2301 & n2304;
  assign n2306 = n2300 & n2305;
  assign n2307 = n472 & ~n2306;
  assign n2308 = n1511 & ~n2307;
  assign n2309 = n379 & ~n2211;
  assign n2310 = n1489 & n2218;
  assign n2311 = ~n1944 & n2310;
  assign n2312 = n898 & ~n2311;
  assign n2313 = ~n2309 & ~n2312;
  assign n2314 = n2308 & n2313;
  assign n2315 = n722 & ~n1014;
  assign n2316 = n2162 & n2315;
  assign n2317 = n1106 & n1796;
  assign n2318 = ~n609 & n2317;
  assign n2319 = ~n1062 & n1254;
  assign n2320 = n2318 & n2319;
  assign n2321 = n2032 & n2320;
  assign n2322 = n2316 & n2321;
  assign n2323 = n1533 & n2322;
  assign n2324 = n472 & ~n2323;
  assign n2325 = n2314 & ~n2324;
  assign n2326 = ~n2298 & n2325;
  assign n2327 = ~n451 & ~n1464;
  assign n2328 = ~n295 & n2327;
  assign n2329 = n1224 & n1533;
  assign n2330 = n2328 & n2329;
  assign n2331 = ~n1010 & ~n1107;
  assign n2332 = n1106 & n2331;
  assign n2333 = ~n1099 & n1572;
  assign n2334 = n2332 & n2333;
  assign n2335 = n2330 & n2334;
  assign n2336 = n2225 & n2285;
  assign n2337 = n2335 & n2336;
  assign n2338 = ~n1503 & n1929;
  assign n2339 = ~n253 & n2338;
  assign n2340 = ~n515 & n2339;
  assign n2341 = n1776 & n2340;
  assign n2342 = n2337 & n2341;
  assign n2343 = ~n492 & n1998;
  assign n2344 = n1909 & n2343;
  assign n2345 = n766 & n2344;
  assign n2346 = ~n181 & ~n609;
  assign n2347 = ~n1904 & n2346;
  assign n2348 = ~n465 & ~n1456;
  assign n2349 = ~n586 & n2348;
  assign n2350 = n2347 & n2349;
  assign n2351 = n2345 & n2350;
  assign n2352 = ~n220 & n1138;
  assign n2353 = n1984 & n2352;
  assign n2354 = n2163 & n2353;
  assign n2355 = n2351 & n2354;
  assign n2356 = n2342 & n2355;
  assign n2357 = n898 & ~n2356;
  assign n2358 = ~n291 & ~n798;
  assign n2359 = n1521 & n2358;
  assign n2360 = ~n393 & n2359;
  assign n2361 = ~n1123 & n2360;
  assign n2362 = ~n1442 & n2361;
  assign n2363 = n898 & ~n2362;
  assign n2364 = n1909 & n2360;
  assign n2365 = ~n1123 & n2364;
  assign n2366 = n472 & ~n2365;
  assign n2367 = n898 & ~n2286;
  assign n2368 = n1795 & n2277;
  assign n2369 = n379 & ~n2368;
  assign n2370 = n379 & n2112;
  assign n2371 = n472 & ~n2352;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n2369 & n2372;
  assign n2374 = ~n2367 & n2373;
  assign n2375 = ~n2366 & n2374;
  assign n2376 = ~n2363 & n2375;
  assign n2377 = ~n2357 & n2376;
  assign n2378 = ~n1938 & n2327;
  assign n2379 = ~n174 & n2218;
  assign n2380 = n2207 & n2379;
  assign n2381 = n2378 & n2380;
  assign n2382 = n472 & ~n2381;
  assign n2383 = n1080 & n2093;
  assign n2384 = ~n173 & n2383;
  assign n2385 = n898 & ~n2384;
  assign n2386 = ~n2382 & ~n2385;
  assign n2387 = ~n450 & ~n1016;
  assign n2388 = n71 & ~n2387;
  assign n2389 = n1166 & ~n2388;
  assign n2390 = n2101 & n2389;
  assign n2391 = n472 & ~n2390;
  assign n2392 = n1223 & n1810;
  assign n2393 = ~n1438 & n1954;
  assign n2394 = ~n984 & n2393;
  assign n2395 = n2262 & n2394;
  assign n2396 = n2392 & n2395;
  assign n2397 = ~n128 & ~n453;
  assign n2398 = n2396 & n2397;
  assign n2399 = n379 & ~n2398;
  assign n2400 = ~n2391 & ~n2399;
  assign n2401 = n2386 & n2400;
  assign n2402 = n2377 & n2401;
  assign o_12_ = ~n2326 | ~n2402;
  assign n2404 = ~n244 & n1564;
  assign n2405 = ~n1456 & n2404;
  assign n2406 = ~n570 & ~n1443;
  assign n2407 = ~n596 & ~n1137;
  assign n2408 = ~n181 & n2407;
  assign n2409 = n2406 & n2408;
  assign n2410 = n2405 & n2409;
  assign n2411 = ~n1062 & ~n1923;
  assign n2412 = n678 & n2270;
  assign n2413 = n2264 & n2412;
  assign n2414 = ~n167 & n2413;
  assign n2415 = n280 & n2414;
  assign n2416 = ~n179 & ~n1024;
  assign n2417 = ~n1904 & n2416;
  assign n2418 = ~n504 & n2417;
  assign n2419 = n2415 & n2418;
  assign n2420 = n2411 & n2419;
  assign n2421 = n2410 & n2420;
  assign n2422 = ~i_8_ & ~n2421;
  assign n2423 = ~i_8_ & ~n2161;
  assign n2424 = ~n635 & ~n1563;
  assign n2425 = ~n1024 & n2424;
  assign n2426 = ~n1062 & ~n1449;
  assign n2427 = ~n245 & n2426;
  assign n2428 = n2425 & n2427;
  assign n2429 = ~n390 & n1899;
  assign n2430 = n2428 & ~n2429;
  assign n2431 = i_8_ & ~n2430;
  assign n2432 = ~n464 & ~n2431;
  assign n2433 = ~n2423 & n2432;
  assign n2434 = ~n607 & ~n1537;
  assign n2435 = i_8_ & n2434;
  assign n2436 = ~n759 & ~n1107;
  assign n2437 = n1488 & n2436;
  assign n2438 = ~i_8_ & ~n1040;
  assign n2439 = ~n1010 & ~n1552;
  assign n2440 = n2438 & n2439;
  assign n2441 = n2437 & n2440;
  assign n2442 = ~n2435 & ~n2441;
  assign n2443 = ~n515 & n2215;
  assign n2444 = ~n2442 & n2443;
  assign n2445 = n1184 & n2157;
  assign n2446 = i_8_ & ~n2445;
  assign n2447 = ~i_8_ & n1011;
  assign n2448 = n2250 & ~n2447;
  assign n2449 = n2290 & n2448;
  assign n2450 = ~n2446 & n2449;
  assign n2451 = n2444 & n2450;
  assign n2452 = n2433 & n2451;
  assign n2453 = ~n143 & n517;
  assign n2454 = n2346 & n2453;
  assign n2455 = n2262 & n2454;
  assign n2456 = ~n1171 & n1609;
  assign n2457 = ~n1047 & n2456;
  assign n2458 = n2455 & n2457;
  assign n2459 = n2335 & n2458;
  assign n2460 = n1746 & n2459;
  assign n2461 = i_8_ & ~n2460;
  assign n2462 = ~n1157 & n2338;
  assign n2463 = n2129 & n2269;
  assign n2464 = ~n456 & ~n1938;
  assign n2465 = n2152 & n2464;
  assign n2466 = n2463 & n2465;
  assign n2467 = n2462 & n2466;
  assign n2468 = ~n2461 & n2467;
  assign n2469 = n1520 & n2327;
  assign n2470 = ~i_8_ & ~n2469;
  assign n2471 = n1082 & ~n2470;
  assign n2472 = ~n179 & ~n279;
  assign n2473 = n1520 & n2472;
  assign n2474 = n2212 & n2218;
  assign n2475 = n2473 & n2474;
  assign n2476 = i_8_ & ~n2475;
  assign n2477 = ~n176 & ~n1168;
  assign n2478 = ~n507 & ~n597;
  assign n2479 = ~n174 & n2478;
  assign n2480 = n2477 & n2479;
  assign n2481 = ~n2476 & n2480;
  assign n2482 = n2471 & n2481;
  assign n2483 = n2468 & n2482;
  assign n2484 = n2452 & n2483;
  assign n2485 = ~n2422 & n2484;
  assign n2486 = n380 & ~n2485;
  assign n2487 = n72 & n223;
  assign n2488 = ~n1087 & ~n2487;
  assign n2489 = n380 & ~n2488;
  assign n2490 = n170 & ~n1164;
  assign n2491 = n219 & ~n2490;
  assign n2492 = ~n2489 & ~n2491;
  assign n2493 = n774 & n2492;
  assign n2494 = ~n1032 & n1142;
  assign n2495 = n2358 & n2494;
  assign n2496 = ~n82 & ~n86;
  assign n2497 = ~n223 & n2496;
  assign n2498 = n1039 & ~n2497;
  assign n2499 = n2495 & ~n2498;
  assign n2500 = n219 & ~n2499;
  assign n2501 = n913 & n2275;
  assign n2502 = ~n1191 & n2501;
  assign n2503 = ~n180 & n2502;
  assign n2504 = n219 & ~n2503;
  assign n2505 = ~n230 & ~n596;
  assign n2506 = ~n1191 & n1484;
  assign n2507 = n2352 & n2506;
  assign n2508 = n2505 & n2507;
  assign n2509 = n309 & ~n2508;
  assign n2510 = ~n739 & ~n2509;
  assign n2511 = ~n2504 & n2510;
  assign n2512 = ~n2500 & n2511;
  assign n2513 = ~n1863 & n2358;
  assign n2514 = n1247 & n2513;
  assign n2515 = ~n1032 & n2514;
  assign n2516 = n309 & ~n2515;
  assign n2517 = n219 & ~n2434;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = n2512 & n2518;
  assign n2520 = n2493 & n2519;
  assign o_13_ = n2486 | ~n2520;
  assign n2522 = ~i_2_ & o_14_;
  assign n2523 = ~i_0_ & i_2_;
  assign o_15_ = n2522 | n2523;
  assign n2525 = ~n1054 & ~n1515;
  assign n2526 = n2268 & n2515;
  assign n2527 = n2525 & n2526;
  assign n2528 = n2111 & n2527;
  assign n2529 = n309 & ~n2528;
  assign n2530 = n1138 & n2271;
  assign n2531 = ~n1011 & n2530;
  assign n2532 = n243 & ~n2531;
  assign n2533 = n1619 & ~n2532;
  assign n2534 = ~n2529 & n2533;
  assign n2535 = n2092 & n2318;
  assign n2536 = n2207 & n2535;
  assign n2537 = n2365 & n2536;
  assign n2538 = n1183 & n2352;
  assign n2539 = i_13_ & n679;
  assign n2540 = ~n1107 & ~n2539;
  assign n2541 = n1548 & n1959;
  assign n2542 = ~n1040 & n2541;
  assign n2543 = n2540 & n2542;
  assign n2544 = n2538 & n2543;
  assign n2545 = n2215 & n2396;
  assign n2546 = n2544 & n2545;
  assign n2547 = n2537 & n2546;
  assign n2548 = n472 & ~n2547;
  assign n2549 = ~n1170 & n2530;
  assign n2550 = ~n167 & n2549;
  assign n2551 = n307 & ~n2550;
  assign n2552 = ~n2548 & ~n2551;
  assign n2553 = ~n176 & n2473;
  assign n2554 = n1082 & n2553;
  assign n2555 = ~n606 & ~n2554;
  assign n2556 = n273 & ~n2300;
  assign n2557 = n243 & ~n2153;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = n273 & ~n2315;
  assign n2560 = n358 & ~n2378;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = ~n2110 & n2561;
  assign n2563 = n2558 & n2562;
  assign n2564 = ~n2555 & n2563;
  assign n2565 = ~n740 & n993;
  assign n2566 = n1360 & n2565;
  assign n2567 = n2564 & n2566;
  assign n2568 = n2552 & n2567;
  assign n2569 = n2534 & n2568;
  assign n2570 = n307 & ~n1775;
  assign n2571 = n1080 & ~n1139;
  assign n2572 = n2472 & n2571;
  assign n2573 = n2153 & n2572;
  assign n2574 = ~n2130 & n2573;
  assign n2575 = n307 & ~n2574;
  assign n2576 = n243 & ~n1793;
  assign n2577 = ~n1020 & ~n2576;
  assign n2578 = ~n2575 & n2577;
  assign n2579 = ~n2570 & n2578;
  assign n2580 = n273 & ~n2162;
  assign n2581 = ~n472 & ~n2580;
  assign n2582 = ~n2316 & ~n2581;
  assign n2583 = n309 & ~n1793;
  assign n2584 = ~n635 & n2426;
  assign n2585 = n358 & ~n2584;
  assign n2586 = ~n2583 & ~n2585;
  assign n2587 = ~n1196 & n2586;
  assign n2588 = ~n2582 & n2587;
  assign n2589 = n1930 & n2437;
  assign n2590 = n307 & ~n2589;
  assign n2591 = n2588 & ~n2590;
  assign n2592 = ~n291 & n1605;
  assign n2593 = ~n983 & n2592;
  assign n2594 = n2353 & n2593;
  assign n2595 = n1141 & n1795;
  assign n2596 = n1595 & n2595;
  assign n2597 = n2092 & n2596;
  assign n2598 = n2594 & n2597;
  assign n2599 = n273 & ~n2598;
  assign n2600 = ~n570 & n2212;
  assign n2601 = n2428 & n2600;
  assign n2602 = n309 & ~n2601;
  assign n2603 = ~n1154 & ~n1465;
  assign n2604 = n2225 & n2603;
  assign n2605 = n2211 & n2604;
  assign n2606 = n358 & ~n2605;
  assign n2607 = ~n2602 & ~n2606;
  assign n2608 = ~n2599 & n2607;
  assign n2609 = n2591 & n2608;
  assign n2610 = n2579 & n2609;
  assign n2611 = n1236 & n2610;
  assign n2612 = n1973 & n2611;
  assign n2613 = ~n257 & n2495;
  assign n2614 = ~n1497 & n2613;
  assign n2615 = n243 & ~n2614;
  assign n2616 = n472 & ~n1259;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = n243 & ~n2208;
  assign n2619 = ~n244 & n2425;
  assign n2620 = n243 & ~n2619;
  assign n2621 = ~n1624 & ~n2620;
  assign n2622 = ~n2618 & n2621;
  assign n2623 = n358 & ~n2515;
  assign n2624 = n307 & ~n2365;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = ~n2202 & n2625;
  assign n2627 = n2622 & n2626;
  assign n2628 = n2617 & n2627;
  assign n2629 = n490 & n1848;
  assign n2630 = n2628 & n2629;
  assign n2631 = n2612 & n2630;
  assign n2632 = n650 & n2631;
  assign n2633 = n2569 & n2632;
  assign o_16_ = n164 & ~n2633;
  assign n2635 = n380 & ~n2433;
  assign n2636 = n273 & ~n2361;
  assign n2637 = ~n1262 & ~n2636;
  assign n2638 = n313 & ~n2364;
  assign n2639 = ~n1538 & ~n2638;
  assign n2640 = n2637 & n2639;
  assign n2641 = n2518 & n2640;
  assign n2642 = ~n1537 & n2614;
  assign n2643 = n265 & ~n2642;
  assign n2644 = n242 & n1443;
  assign n2645 = ~n505 & ~n1904;
  assign n2646 = ~n1040 & n2645;
  assign n2647 = ~n1244 & n2646;
  assign n2648 = n243 & ~n2647;
  assign n2649 = ~n2644 & ~n2648;
  assign n2650 = ~n1094 & n2649;
  assign n2651 = ~n2643 & n2650;
  assign n2652 = n313 & n1443;
  assign n2653 = n2043 & ~n2652;
  assign n2654 = ~n1537 & n2359;
  assign n2655 = n275 & ~n2654;
  assign n2656 = ~n1040 & n2406;
  assign n2657 = n292 & ~n2656;
  assign n2658 = n219 & ~n2600;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = ~n2655 & n2659;
  assign n2661 = i_8_ & n2218;
  assign n2662 = n249 & ~n2474;
  assign n2663 = ~n2661 & n2662;
  assign n2664 = n307 & ~n1259;
  assign n2665 = ~n2083 & ~n2664;
  assign n2666 = ~n2663 & n2665;
  assign n2667 = n2660 & n2666;
  assign n2668 = n2653 & n2667;
  assign n2669 = ~n2363 & n2668;
  assign n2670 = n2651 & n2669;
  assign n2671 = n2641 & n2670;
  assign n2672 = ~n2635 & n2671;
  assign n2673 = n2131 & n2411;
  assign n2674 = n243 & ~n2673;
  assign n2675 = n2315 & n2411;
  assign n2676 = ~n635 & n2169;
  assign n2677 = n2675 & n2676;
  assign n2678 = i_8_ & ~n2677;
  assign n2679 = ~n245 & n1564;
  assign n2680 = ~n634 & n2679;
  assign n2681 = ~i_8_ & ~n2680;
  assign n2682 = ~n1017 & ~n2681;
  assign n2683 = ~n464 & n2682;
  assign n2684 = ~n2678 & n2683;
  assign n2685 = n249 & ~n2684;
  assign n2686 = ~n2674 & ~n2685;
  assign n2687 = n1254 & n1793;
  assign n2688 = n2679 & n2687;
  assign n2689 = n265 & ~n2688;
  assign n2690 = ~n1093 & ~n2689;
  assign n2691 = ~n839 & n2690;
  assign n2692 = ~n571 & n2691;
  assign n2693 = ~n899 & ~n2161;
  assign n2694 = ~n1794 & ~n2693;
  assign n2695 = ~n1197 & n2694;
  assign n2696 = ~n2620 & n2695;
  assign n2697 = ~n707 & n1294;
  assign n2698 = n338 & ~n2697;
  assign n2699 = ~n2170 & ~n2698;
  assign n2700 = ~n2135 & n2699;
  assign n2701 = n2696 & n2700;
  assign n2702 = ~n1391 & ~n1937;
  assign n2703 = n2701 & n2702;
  assign n2704 = n2692 & n2703;
  assign n2705 = n288 & ~n2292;
  assign n2706 = ~i_8_ & n1923;
  assign n2707 = ~n1023 & ~n2706;
  assign n2708 = n2404 & n2707;
  assign n2709 = n1792 & n2708;
  assign n2710 = n288 & ~n2709;
  assign n2711 = n273 & ~n2286;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = ~n2705 & n2712;
  assign n2714 = n1222 & n2588;
  assign n2715 = n2713 & n2714;
  assign n2716 = ~n973 & ~n2411;
  assign n2717 = n430 & n1542;
  assign n2718 = n472 & ~n1254;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2716 & n2719;
  assign n2721 = n1019 & n2169;
  assign n2722 = ~n2130 & n2721;
  assign n2723 = n219 & ~n2722;
  assign n2724 = n2319 & n2697;
  assign n2725 = ~n1157 & n2724;
  assign n2726 = n326 & ~n2725;
  assign n2727 = ~n2723 & ~n2726;
  assign n2728 = n2720 & n2727;
  assign n2729 = n2715 & n2728;
  assign n2730 = n2704 & n2729;
  assign n2731 = n2686 & n2730;
  assign n2732 = n2672 & n2731;
  assign n2733 = ~n2154 & n2352;
  assign n2734 = ~n596 & n2733;
  assign n2735 = n249 & ~n2734;
  assign n2736 = n2579 & ~n2735;
  assign n2737 = ~n182 & n275;
  assign n2738 = ~n225 & n2368;
  assign n2739 = n307 & ~n2738;
  assign n2740 = ~n2737 & ~n2739;
  assign n2741 = ~n2079 & n2740;
  assign n2742 = n2736 & n2741;
  assign n2743 = n2628 & n2742;
  assign n2744 = n2063 & n2514;
  assign n2745 = ~n506 & n2744;
  assign n2746 = n292 & ~n2745;
  assign n2747 = n2561 & ~n2746;
  assign n2748 = n1254 & n2353;
  assign n2749 = n2368 & n2748;
  assign n2750 = n273 & ~n2749;
  assign n2751 = ~n1194 & ~n2750;
  assign n2752 = n2747 & n2751;
  assign n2753 = n181 & n292;
  assign n2754 = n358 & n510;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = n1747 & n2208;
  assign n2757 = n2032 & n2756;
  assign n2758 = n313 & ~n2757;
  assign n2759 = n2755 & ~n2758;
  assign n2760 = n2752 & n2759;
  assign n2761 = n508 & ~n676;
  assign n2762 = ~n180 & ~n220;
  assign n2763 = n2293 & n2762;
  assign n2764 = n2761 & n2763;
  assign n2765 = n898 & ~n2764;
  assign n2766 = ~n742 & n2125;
  assign n2767 = ~n2765 & n2766;
  assign n2768 = n177 & ~n225;
  assign n2769 = ~n1008 & n2768;
  assign n2770 = n292 & ~n2769;
  assign n2771 = n1681 & n2397;
  assign n2772 = n2505 & n2771;
  assign n2773 = n292 & ~n2772;
  assign n2774 = n358 & ~n2152;
  assign n2775 = ~n1826 & ~n2774;
  assign n2776 = n358 & ~n2474;
  assign n2777 = n2775 & ~n2776;
  assign n2778 = ~n2773 & n2777;
  assign n2779 = ~n2770 & n2778;
  assign n2780 = n218 & ~n2408;
  assign n2781 = n217 & n453;
  assign n2782 = ~n1458 & ~n2781;
  assign n2783 = ~n2780 & n2782;
  assign n2784 = n273 & ~n1784;
  assign n2785 = n472 & ~n1605;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = n265 & ~n1259;
  assign n2788 = n2786 & ~n2787;
  assign n2789 = n2783 & n2788;
  assign n2790 = ~n359 & n506;
  assign n2791 = ~n995 & ~n2790;
  assign n2792 = ~n998 & ~n2221;
  assign n2793 = n292 & ~n2426;
  assign n2794 = n2792 & ~n2793;
  assign n2795 = n2791 & n2794;
  assign n2796 = ~n606 & n607;
  assign n2797 = n2795 & ~n2796;
  assign n2798 = n2789 & n2797;
  assign n2799 = n2779 & n2798;
  assign n2800 = n2767 & n2799;
  assign n2801 = n1126 & ~n1722;
  assign n2802 = n275 & ~n2368;
  assign n2803 = ~n2801 & ~n2802;
  assign n2804 = ~n1474 & n2803;
  assign n2805 = ~n1279 & n2804;
  assign n2806 = ~n2281 & n2805;
  assign n2807 = n358 & ~n2276;
  assign n2808 = n128 & ~n695;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = n1438 & ~n1519;
  assign n2811 = n570 & ~n899;
  assign n2812 = ~n753 & n1040;
  assign n2813 = ~n2811 & ~n2812;
  assign n2814 = ~n2810 & n2813;
  assign n2815 = n1982 & n2814;
  assign n2816 = n784 & n2815;
  assign n2817 = n2809 & n2816;
  assign n2818 = n2806 & n2817;
  assign n2819 = n2800 & n2818;
  assign n2820 = n2760 & n2819;
  assign n2821 = n2743 & n2820;
  assign n2822 = n174 & n307;
  assign n2823 = n2378 & n2553;
  assign n2824 = n2479 & n2823;
  assign n2825 = n275 & ~n2824;
  assign n2826 = n2111 & n2120;
  assign n2827 = n430 & ~n2826;
  assign n2828 = ~n2825 & ~n2827;
  assign n2829 = ~n2822 & n2828;
  assign n2830 = n380 & ~n2482;
  assign n2831 = n2115 & ~n2830;
  assign n2832 = n2829 & n2831;
  assign n2833 = n2768 & n2826;
  assign n2834 = n1775 & n2833;
  assign n2835 = n265 & ~n2834;
  assign n2836 = ~n669 & ~n2835;
  assign n2837 = ~i_8_ & ~n903;
  assign n2838 = ~n451 & ~n2837;
  assign n2839 = n325 & ~n2838;
  assign n2840 = ~n328 & ~n812;
  assign n2841 = ~n2839 & n2840;
  assign n2842 = ~n2570 & n2841;
  assign n2843 = ~n2618 & n2842;
  assign n2844 = n275 & n1078;
  assign n2845 = ~n2231 & ~n2844;
  assign n2846 = n338 & ~n1081;
  assign n2847 = n265 & n1139;
  assign n2848 = n174 & n243;
  assign n2849 = n379 & n1168;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2847 & n2850;
  assign n2852 = ~n2846 & n2851;
  assign n2853 = n2845 & n2852;
  assign n2854 = n358 & n1168;
  assign n2855 = n292 & ~n2111;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = ~n508 & n666;
  assign n2858 = n2856 & ~n2857;
  assign n2859 = ~n994 & n2858;
  assign n2860 = n1775 & n2572;
  assign n2861 = n292 & ~n2860;
  assign n2862 = n2859 & ~n2861;
  assign n2863 = n2853 & n2862;
  assign n2864 = n2843 & n2863;
  assign n2865 = n2836 & n2864;
  assign n2866 = n2479 & n2554;
  assign n2867 = n358 & ~n2866;
  assign n2868 = n307 & ~n2206;
  assign n2869 = n382 & ~n2472;
  assign n2870 = ~n309 & ~n898;
  assign n2871 = ~n2327 & ~n2870;
  assign n2872 = ~n2869 & ~n2871;
  assign n2873 = ~n2868 & n2872;
  assign n2874 = ~n2867 & n2873;
  assign n2875 = n2386 & n2874;
  assign n2876 = n2865 & n2875;
  assign n2877 = n2832 & n2876;
  assign n2878 = n2152 & n2508;
  assign n2879 = n243 & ~n2878;
  assign n2880 = n182 & ~n452;
  assign n2881 = n1276 & n2502;
  assign n2882 = n2880 & n2881;
  assign n2883 = n265 & ~n2882;
  assign n2884 = ~n2879 & ~n2883;
  assign n2885 = n1922 & n2375;
  assign n2886 = n2884 & n2885;
  assign n2887 = n1253 & n2512;
  assign n2888 = n2886 & n2887;
  assign n2889 = n2877 & n2888;
  assign n2890 = n2821 & n2889;
  assign n2891 = n2732 & n2890;
  assign o_17_ = n164 & ~n2891;
  assign n2893 = ~n115 & n1779;
  assign n2894 = n1445 & ~n2893;
  assign n2895 = ~n277 & ~n2487;
  assign n2896 = i_8_ & ~n2895;
  assign n2897 = n170 & ~n2896;
  assign n2898 = n2228 & n2897;
  assign n2899 = ~n278 & n2898;
  assign n2900 = ~n586 & n2899;
  assign n2901 = n249 & ~n2900;
  assign n2902 = ~n278 & n1931;
  assign n2903 = ~n700 & ~n2902;
  assign n2904 = ~n695 & n1099;
  assign n2905 = n309 & ~n1167;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~n2903 & n2906;
  assign n2908 = ~n2901 & n2907;
  assign n2909 = ~n2894 & n2908;
  assign n2910 = ~n2121 & ~n2229;
  assign n2911 = n358 & ~n2227;
  assign n2912 = ~n88 & n2120;
  assign n2913 = n2225 & n2912;
  assign n2914 = n292 & ~n2913;
  assign n2915 = ~n2911 & ~n2914;
  assign n2916 = n325 & n457;
  assign n2917 = ~n588 & ~n2916;
  assign n2918 = ~n426 & ~n503;
  assign n2919 = n2917 & n2918;
  assign n2920 = ~n2770 & n2919;
  assign n2921 = n2915 & n2920;
  assign n2922 = ~n989 & ~n2370;
  assign n2923 = n469 & ~n1778;
  assign n2924 = ~n651 & ~n2923;
  assign n2925 = n358 & ~n2111;
  assign n2926 = n292 & n1154;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = ~n366 & n2927;
  assign n2929 = n2924 & n2928;
  assign n2930 = n2922 & n2929;
  assign n2931 = ~n1979 & n2492;
  assign n2932 = n358 & ~n1931;
  assign n2933 = n167 & n380;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = n2931 & n2934;
  assign n2936 = n2930 & n2935;
  assign n2937 = n2921 & n2936;
  assign n2938 = ~n911 & ~n2094;
  assign n2939 = ~n2168 & ~n2938;
  assign n2940 = ~n2205 & n2258;
  assign n2941 = n2939 & n2940;
  assign n2942 = n168 & n898;
  assign n2943 = ~n522 & n577;
  assign n2944 = ~n1614 & ~n2943;
  assign n2945 = ~n2942 & n2944;
  assign n2946 = n744 & n2945;
  assign n2947 = n859 & n1883;
  assign n2948 = ~n2226 & ~n2947;
  assign n2949 = ~n1630 & ~n2948;
  assign n2950 = n2946 & n2949;
  assign n2951 = n2941 & n2950;
  assign n2952 = n1791 & n2951;
  assign n2953 = n2937 & n2952;
  assign n2954 = n2910 & n2953;
  assign n2955 = n2909 & n2954;
  assign n2956 = n2224 & ~n2391;
  assign n2957 = n358 & ~n2100;
  assign n2958 = ~n277 & n587;
  assign n2959 = ~n168 & ~n468;
  assign n2960 = n2488 & n2959;
  assign n2961 = n2958 & n2960;
  assign n2962 = n292 & ~n2961;
  assign n2963 = ~n2957 & ~n2962;
  assign n2964 = n169 & n292;
  assign n2965 = n358 & ~n2099;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = n2963 & n2966;
  assign n2968 = n2956 & n2967;
  assign n2969 = n2955 & n2968;
  assign n2970 = ~n754 & n1165;
  assign n2971 = n242 & ~n2255;
  assign n2972 = ~n465 & n2958;
  assign n2973 = n243 & ~n2972;
  assign n2974 = ~n569 & ~n2973;
  assign n2975 = ~n2971 & n2974;
  assign n2976 = ~n2970 & n2975;
  assign n2977 = n2105 & n2976;
  assign n2978 = n2671 & n2977;
  assign n2979 = n2969 & n2978;
  assign n2980 = ~n515 & ~n767;
  assign n2981 = n1181 & n2980;
  assign n2982 = ~i_8_ & ~n2981;
  assign n2983 = n2215 & ~n2982;
  assign n2984 = n288 & ~n2983;
  assign n2985 = n358 & ~n2745;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = n309 & ~n2299;
  assign n2988 = n380 & ~n2338;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = ~n2500 & n2989;
  assign n2991 = ~n2366 & n2990;
  assign n2992 = n898 & ~n2340;
  assign n2993 = n265 & n1035;
  assign n2994 = n1181 & ~n1552;
  assign n2995 = ~n2870 & ~n2994;
  assign n2996 = ~n2993 & ~n2995;
  assign n2997 = ~n2776 & n2996;
  assign n2998 = ~n2992 & n2997;
  assign n2999 = n2233 & n2998;
  assign n3000 = n2314 & n2999;
  assign n3001 = n2991 & n3000;
  assign n3002 = n380 & ~n2444;
  assign n3003 = ~n515 & ~n1010;
  assign n3004 = n1909 & n3003;
  assign n3005 = i_8_ & ~n3004;
  assign n3006 = n1930 & ~n3005;
  assign n3007 = n272 & ~n3006;
  assign n3008 = n2191 & ~n3007;
  assign n3009 = n1488 & ~n2539;
  assign n3010 = ~n1263 & n3009;
  assign n3011 = n313 & ~n3010;
  assign n3012 = ~n2556 & ~n3011;
  assign n3013 = n3008 & n3012;
  assign n3014 = n358 & n1010;
  assign n3015 = n1488 & n1929;
  assign n3016 = n1565 & n3015;
  assign n3017 = n288 & ~n3016;
  assign n3018 = ~n515 & n2436;
  assign n3019 = n358 & ~n3018;
  assign n3020 = ~n3017 & ~n3019;
  assign n3021 = ~n3014 & n3020;
  assign n3022 = ~n2746 & n3021;
  assign n3023 = n3013 & n3022;
  assign n3024 = ~n3002 & n3023;
  assign n3025 = n3001 & n3024;
  assign n3026 = n2986 & n3025;
  assign n3027 = n149 & ~n2387;
  assign n3028 = ~n767 & ~n1035;
  assign n3029 = ~n3027 & n3028;
  assign n3030 = n3016 & n3029;
  assign n3031 = n2642 & n3030;
  assign n3032 = n243 & ~n3031;
  assign n3033 = ~n1195 & ~n3032;
  assign n3034 = n1259 & n2210;
  assign n3035 = n2439 & n3034;
  assign n3036 = n2310 & n3035;
  assign n3037 = n2340 & n3036;
  assign n3038 = n265 & ~n3037;
  assign n3039 = n1180 & ~n1944;
  assign n3040 = n242 & ~n3039;
  assign n3041 = ~n3038 & ~n3040;
  assign n3042 = n3033 & n3041;
  assign n3043 = n1141 & n2212;
  assign n3044 = ~n1503 & n3043;
  assign n3045 = n3004 & n3044;
  assign n3046 = n307 & ~n3045;
  assign n3047 = n1929 & n3003;
  assign n3048 = n2540 & n3047;
  assign n3049 = ~n506 & n1565;
  assign n3050 = n1247 & n3049;
  assign n3051 = n3048 & n3050;
  assign n3052 = n1489 & n3051;
  assign n3053 = ~i_8_ & ~n3052;
  assign n3054 = n2215 & ~n3053;
  assign n3055 = n2654 & n3054;
  assign n3056 = n249 & ~n3055;
  assign n3057 = ~n2590 & ~n3056;
  assign n3058 = ~n3046 & n3057;
  assign n3059 = n3042 & n3058;
  assign n3060 = n3026 & n3059;
  assign n3061 = n2979 & n3060;
  assign n3062 = n2877 & n3061;
  assign o_18_ = n164 & ~n3062;
  assign n3064 = n265 & ~n1114;
  assign n3065 = ~n1532 & ~n3064;
  assign n3066 = n338 & ~n3065;
  assign n3067 = n1002 & ~n3066;
  assign n3068 = ~n1047 & n2450;
  assign n3069 = n380 & ~n3068;
  assign n3070 = ~n695 & n1047;
  assign n3071 = n2285 & ~n2706;
  assign n3072 = n272 & ~n3071;
  assign n3073 = ~n3070 & ~n3072;
  assign n3074 = ~n2253 & n3073;
  assign n3075 = n275 & ~n2249;
  assign n3076 = ~n392 & ~n3075;
  assign n3077 = ~n337 & ~n3076;
  assign n3078 = ~n985 & n1953;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = n3074 & n3079;
  assign n3081 = ~n3069 & n3080;
  assign n3082 = n3067 & n3081;
  assign n3083 = ~n2149 & ~n2298;
  assign n3084 = n695 & n753;
  assign n3085 = n1446 & ~n3084;
  assign n3086 = ~n696 & n1113;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n308 & ~n2218;
  assign n3089 = ~n309 & ~n3088;
  assign n3090 = ~n2474 & ~n3089;
  assign n3091 = n358 & ~n2155;
  assign n3092 = n288 & ~n2156;
  assign n3093 = n292 & ~n2584;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = ~n3091 & n3094;
  assign n3096 = n273 & ~n2293;
  assign n3097 = n3095 & ~n3096;
  assign n3098 = ~n547 & ~n1177;
  assign n3099 = ~n1350 & n3098;
  assign n3100 = ~n1115 & n3099;
  assign n3101 = ~n2367 & n3100;
  assign n3102 = n3097 & n3101;
  assign n3103 = ~n3090 & n3102;
  assign n3104 = n3087 & n3103;
  assign n3105 = n3083 & n3104;
  assign n3106 = n358 & ~n2289;
  assign n3107 = ~n1011 & ~n1532;
  assign n3108 = ~n392 & n3107;
  assign n3109 = ~i_8_ & ~n3108;
  assign n3110 = n2291 & ~n3109;
  assign n3111 = n288 & ~n3110;
  assign n3112 = ~n3106 & ~n3111;
  assign n3113 = ~i_8_ & n224;
  assign n3114 = ~i_15_ & ~n3113;
  assign n3115 = n153 & ~n3114;
  assign n3116 = ~n2497 & n3115;
  assign n3117 = n1600 & ~n3116;
  assign n3118 = ~n2141 & n3117;
  assign n3119 = n242 & ~n3118;
  assign n3120 = ~n1188 & ~n3119;
  assign n3121 = n2217 & n3120;
  assign n3122 = n219 & ~n1183;
  assign n3123 = n482 & n2251;
  assign n3124 = n307 & ~n3123;
  assign n3125 = n281 & n1485;
  assign n3126 = ~n1553 & n3125;
  assign n3127 = n275 & ~n3126;
  assign n3128 = ~n3124 & ~n3127;
  assign n3129 = n758 & n3128;
  assign n3130 = ~n3122 & n3129;
  assign n3131 = n3121 & n3130;
  assign n3132 = n3112 & n3131;
  assign n3133 = n3105 & n3132;
  assign n3134 = n3082 & n3133;
  assign n3135 = n3060 & n3134;
  assign n3136 = n2732 & n3135;
  assign o_19_ = n164 & ~n3136;
  assign n3138 = n2651 & n2884;
  assign n3139 = n3042 & n3138;
  assign n3140 = n2239 & n2826;
  assign n3141 = n2453 & n3140;
  assign n3142 = n1793 & ~n1949;
  assign n3143 = n3141 & n3142;
  assign n3144 = ~n1170 & n1918;
  assign n3145 = n296 & n1756;
  assign n3146 = ~n1060 & n3145;
  assign n3147 = n3144 & n3146;
  assign n3148 = n1106 & n3147;
  assign n3149 = n3143 & n3148;
  assign n3150 = n2412 & n3149;
  assign n3151 = n243 & ~n3150;
  assign n3152 = n1198 & ~n2079;
  assign n3153 = ~n782 & ~n2847;
  assign n3154 = ~n580 & n3153;
  assign n3155 = ~n2674 & n3154;
  assign n3156 = n3152 & n3155;
  assign n3157 = ~n180 & n615;
  assign n3158 = n243 & ~n3157;
  assign n3159 = n2227 & ~n2423;
  assign n3160 = n242 & ~n3159;
  assign n3161 = ~n3158 & ~n3160;
  assign n3162 = n3156 & n3161;
  assign n3163 = n2836 & n3162;
  assign n3164 = n2975 & n3163;
  assign n3165 = n2691 & n3164;
  assign n3166 = n2622 & n3165;
  assign n3167 = ~n3151 & n3166;
  assign n3168 = n1144 & n2349;
  assign n3169 = ~n1008 & n2411;
  assign n3170 = ~n1035 & ~n1532;
  assign n3171 = ~n1126 & ~n1164;
  assign n3172 = ~n717 & n3171;
  assign n3173 = n3170 & n3172;
  assign n3174 = n3169 & n3173;
  assign n3175 = n2419 & n3174;
  assign n3176 = n3168 & n3175;
  assign n3177 = n265 & ~n3176;
  assign n3178 = n3120 & ~n3177;
  assign n3179 = n3167 & n3178;
  assign n3180 = n3139 & n3179;
  assign n3181 = ~n180 & ~n295;
  assign n3182 = ~n181 & n3181;
  assign n3183 = n2453 & n3182;
  assign n3184 = n1910 & n3183;
  assign n3185 = n1609 & n3184;
  assign n3186 = n307 & ~n3185;
  assign n3187 = ~n1024 & n1143;
  assign n3188 = n3169 & n3187;
  assign n3189 = n275 & ~n3188;
  assign n3190 = ~n3186 & ~n3189;
  assign n3191 = ~n2901 & n3190;
  assign n3192 = n2829 & n3191;
  assign n3193 = ~n1615 & n2666;
  assign n3194 = n2686 & n3193;
  assign n3195 = n3192 & n3194;
  assign n3196 = n1918 & n2414;
  assign n3197 = n249 & ~n3196;
  assign n3198 = n1805 & n3128;
  assign n3199 = ~n3197 & n3198;
  assign n3200 = n2742 & n3199;
  assign n3201 = n3058 & n3200;
  assign n3202 = ~o_11_ & n3201;
  assign n3203 = n3195 & n3202;
  assign n3204 = n3180 & n3203;
  assign o_20_ = n164 & ~n3204;
  assign o_21_ = n164 & ~n3180;
  assign n3207 = ~n998 & n2177;
  assign n3208 = ~n579 & ~n988;
  assign n3209 = ~n2857 & n3208;
  assign n3210 = ~n776 & n3209;
  assign o_22_ = ~n3207 | ~n3210;
  assign n3212 = n103 & n274;
  assign n3213 = n60 & n136;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = n60 & n100;
  assign n3216 = ~n97 & ~n3215;
  assign n3217 = n3214 & n3216;
  assign n3218 = n179 & ~n3217;
  assign n3219 = ~n1127 & ~n3218;
  assign n3220 = ~n2205 & n2236;
  assign n3221 = n3219 & n3220;
  assign n3222 = ~n177 & ~n3217;
  assign n3223 = n2224 & ~n3222;
  assign n3224 = i_4_ & n64;
  assign n3225 = i_5_ & n3224;
  assign n3226 = n134 & n3225;
  assign n3227 = n2456 & n3181;
  assign n3228 = ~n128 & n690;
  assign n3229 = n170 & n1931;
  assign n3230 = n3228 & n3229;
  assign n3231 = n2163 & n3230;
  assign n3232 = n3227 & n3231;
  assign n3233 = n358 & ~n3232;
  assign n3234 = n273 & n453;
  assign n3235 = ~n1249 & ~n3234;
  assign n3236 = n292 & ~n1608;
  assign n3237 = ~n1458 & ~n3236;
  assign n3238 = ~n1119 & n3237;
  assign n3239 = n3235 & n3238;
  assign n3240 = ~n1715 & n2856;
  assign n3241 = n3239 & n3240;
  assign n3242 = n1812 & n3241;
  assign n3243 = ~n3233 & n3242;
  assign n3244 = ~n492 & n1568;
  assign n3245 = n1106 & n3244;
  assign n3246 = n2262 & n3245;
  assign n3247 = n288 & ~n3246;
  assign n3248 = n3095 & ~n3247;
  assign n3249 = n2243 & n2915;
  assign n3250 = n3248 & n3249;
  assign n3251 = n2779 & n3250;
  assign n3252 = n3243 & n3251;
  assign n3253 = n296 & ~n1126;
  assign n3254 = n2656 & n3253;
  assign n3255 = ~n1045 & ~n1904;
  assign n3256 = ~n609 & n3255;
  assign n3257 = n2155 & n3256;
  assign n3258 = n3254 & n3257;
  assign n3259 = n2860 & n3258;
  assign n3260 = n292 & ~n3259;
  assign n3261 = n2986 & ~n3260;
  assign n3262 = n3252 & n3261;
  assign n3263 = n2201 & n3022;
  assign n3264 = n3262 & n3263;
  assign n3265 = n559 & n678;
  assign n3266 = ~n1011 & n3265;
  assign n3267 = i_8_ & ~n3266;
  assign n3268 = n1015 & n1298;
  assign n3269 = ~n3267 & n3268;
  assign n3270 = n288 & ~n3269;
  assign n3271 = n2963 & ~n3270;
  assign n3272 = ~n2807 & ~n2867;
  assign n3273 = ~n1194 & n2927;
  assign n3274 = n1823 & n3273;
  assign n3275 = ~n2710 & n3274;
  assign n3276 = ~n3111 & n3275;
  assign n3277 = n3272 & n3276;
  assign n3278 = n3271 & n3277;
  assign n3279 = n2151 & n3278;
  assign n3280 = n3264 & n3279;
  assign n3281 = n2172 & n3280;
  assign n3282 = ~n3226 & n3281;
  assign n3283 = n3223 & n3282;
  assign n3284 = n3221 & n3283;
  assign o_23_ = n164 & ~n3284;
  assign n3286 = ~n140 & n1949;
  assign n3287 = ~i_6_ & n3215;
  assign n3288 = ~n186 & n3287;
  assign o_24_ = n3286 | n3288;
  assign n3290 = n313 & n1900;
  assign n3291 = n273 & ~n1931;
  assign n3292 = ~n1127 & ~n3291;
  assign n3293 = ~n3290 & n3292;
  assign n3294 = n820 & n3293;
  assign n3295 = ~n2167 & n3294;
  assign n3296 = n1705 & n2237;
  assign n3297 = n3280 & n3296;
  assign n3298 = n3295 & n3297;
  assign o_25_ = n164 & ~n3298;
  assign n3300 = n2841 & n3100;
  assign n3301 = ~n1219 & ~n2726;
  assign n3302 = n2919 & n3301;
  assign o_26_ = ~n3300 | ~n3302;
  assign n3304 = n109 & n117;
  assign o_27_ = n164 & n3304;
  assign n3306 = ~i_3_ & o_14_;
  assign n3307 = ~i_7_ & n3306;
  assign n3308 = n58 & n135;
  assign n3309 = n65 & n3308;
  assign n3310 = ~n3307 & ~n3309;
  assign n3311 = n66 & n70;
  assign n3312 = ~n134 & n3224;
  assign n3313 = ~i_5_ & n3312;
  assign n3314 = ~n3311 & ~n3313;
  assign n3315 = ~n126 & ~n3287;
  assign n3316 = ~n3213 & n3315;
  assign n3317 = ~n97 & n3316;
  assign n3318 = ~n171 & ~n3317;
  assign n3319 = n3314 & ~n3318;
  assign n3320 = n3310 & n3319;
  assign o_28_ = n164 & ~n3320;
  assign n3322 = n109 & n1878;
  assign n3323 = ~n416 & n3316;
  assign n3324 = n183 & ~n3323;
  assign n3325 = ~n3322 & ~n3324;
  assign n3326 = ~n182 & ~n3317;
  assign n3327 = n3325 & ~n3326;
  assign n3328 = n66 & n73;
  assign n3329 = n194 & n3306;
  assign n3330 = ~n134 & n3225;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = ~n3328 & n3331;
  assign n3333 = n183 & n1859;
  assign n3334 = i_5_ & n109;
  assign n3335 = i_4_ & ~n3334;
  assign n3336 = n3306 & ~n3335;
  assign n3337 = n109 & n3336;
  assign n3338 = ~n3333 & ~n3337;
  assign n3339 = ~n3309 & n3338;
  assign n3340 = n3332 & n3339;
  assign n3341 = n3327 & n3340;
  assign o_29_ = n164 & ~n3341;
  assign n3343 = ~n109 & n3306;
  assign n3344 = ~n96 & ~n136;
  assign n3345 = i_7_ & ~n3344;
  assign n3346 = ~n3336 & ~n3345;
  assign n3347 = ~n3343 & n3346;
  assign n3348 = ~n3318 & ~n3333;
  assign n3349 = n3347 & n3348;
  assign n3350 = n3327 & n3349;
  assign o_30_ = n164 & ~n3350;
  assign n3352 = n59 & n66;
  assign n3353 = n58 & ~n3214;
  assign n3354 = ~n3309 & ~n3353;
  assign o_31_ = n3352 | ~n3354;
  assign n3356 = n109 & n3224;
  assign n3357 = ~n3345 & ~n3356;
  assign o_32_ = n3226 | ~n3357;
  assign n3359 = n144 & ~n3317;
  assign n3360 = ~i_6_ & n3306;
  assign n3361 = n176 & ~n3217;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = ~n3359 & n3362;
  assign n3364 = ~n203 & n3363;
  assign o_33_ = n164 & ~n3364;
  assign n3366 = n2223 & n2713;
  assign n3367 = n2640 & n3366;
  assign n3368 = n1609 & n1756;
  assign n3369 = n1958 & n3368;
  assign n3370 = n273 & ~n3369;
  assign n3371 = ~n3017 & ~n3370;
  assign n3372 = n292 & ~n1298;
  assign n3373 = n58 & n94;
  assign n3374 = n63 & n3373;
  assign n3375 = n274 & n3374;
  assign n3376 = ~n3372 & ~n3375;
  assign n3377 = i_6_ & n3307;
  assign n3378 = ~n2926 & ~n3377;
  assign n3379 = n3376 & n3378;
  assign n3380 = n3338 & n3379;
  assign n3381 = n3371 & n3380;
  assign n3382 = n358 & ~n2981;
  assign n3383 = n167 & ~n3317;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n3325 & n3384;
  assign n3386 = n3381 & n3385;
  assign n3387 = n3272 & n3386;
  assign n3388 = n2967 & n3387;
  assign n3389 = n3367 & n3388;
  assign n3390 = n3013 & n3112;
  assign n3391 = n3221 & n3390;
  assign n3392 = n3262 & n3391;
  assign n3393 = n3389 & n3392;
  assign n3394 = n2760 & n3393;
  assign n3395 = n2173 & n3394;
  assign o_34_ = n164 & ~n3395;
  assign n3397 = ~n1540 & ~n3317;
  assign n3398 = n174 & ~n3217;
  assign n3399 = ~n3397 & ~n3398;
  assign n3400 = ~n1860 & n3399;
  assign o_35_ = n164 & ~n3400;
  assign n3402 = ~n66 & ~n3309;
  assign n3403 = i_4_ & ~n3402;
  assign n3404 = ~n1127 & ~n3403;
  assign n3405 = n100 & n110;
  assign n3406 = n3404 & ~n3405;
  assign n3407 = ~n186 & n3215;
  assign n3408 = n212 & ~n3407;
  assign n3409 = n2238 & n3408;
  assign n3410 = n3282 & n3409;
  assign n3411 = n3406 & n3410;
  assign o_36_ = n164 & ~n3411;
  assign n3413 = ~i_4_ & ~n3402;
  assign n3414 = ~n187 & n3212;
  assign n3415 = n103 & n110;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~n3413 & n3416;
  assign n3418 = ~n199 & n3417;
  assign n3419 = n191 & n3418;
  assign o_37_ = n164 & ~n3419;
  assign o_38_ = n194 & n3224;
  assign o_39_ = n248 & n3224;
endmodule


