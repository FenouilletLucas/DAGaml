// Benchmark "i5" written by ABC on Tue May 16 16:07:50 2017

module i5 ( 
    \V64(3) , \V28(13) , \V52(11) , \V52(10) , \V64(5) , \V28(15) ,
    \V109(3) , \V64(6) , \V28(14) , \V109(2) , \V132(1) , \V64(7) ,
    \V132(0) , \V64(9) , \V28(11) , \V115(3) , \V28(10) , \V115(2) ,
    \V88(1) , \V109(1) , \V16(1) , \V88(2) , \V121(3) , \V16(2) , \V88(3) ,
    \V121(2) , \V16(3) , \V64(13) , \V115(1) , \V88(5) , \V16(5) ,
    \V88(6) , \V16(6) , \V64(15) , \V88(7) , \V16(7) , \V64(14) ,
    \V121(1) , \V88(9) , \V16(9) , \V100(3) , \V100(2) , \V64(11) ,
    \V100(5) , \V64(10) , \V4(0) , \V100(1) , \V4(1) , \V118(3) ,
    \V118(2) , \V52(1) , \V52(2) , \V124(3) , \V52(3) , \V124(2) ,
    \V128(3) , \V100(7) , \V76(13) , \V128(2) , \V100(6) , \V118(1) ,
    \V52(5) , \V100(9) , \V76(15) , \V52(6) , \V76(14) , \V52(7) ,
    \V100(11) , \V124(1) , \V100(10) , \V52(9) , \V128(1) , \V103(3) ,
    \V100(13) , \V76(11) , \V128(0) , \V103(2) , \V76(10) , \V100(15) ,
    \V76(1) , \V100(14) , \V76(2) , \V76(3) , \V103(1) , \V76(5) ,
    \V76(6) , \V76(7) , \V76(9) , \V40(13) , \V88(13) , \V40(15) ,
    \V28(1) , \V40(14) , \V88(15) , \V28(2) , \V88(14) , \V28(3) ,
    \V16(13) , \V40(11) , \V28(5) , \V40(10) , \V16(15) , \V88(11) ,
    \V106(3) , \V28(6) , \V16(14) , \V88(10) , \V106(2) , \V28(7) ,
    \V40(1) , \V2(0) , \V133(0) , \V28(9) , \V40(2) , \V112(3) , \V16(11) ,
    \V2(1) , \V40(3) , \V112(2) , \V16(10) , \V106(1) , \V40(5) , \V40(6) ,
    \V40(7) , \V112(1) , \V52(13) , \V40(9) , \V52(15) , \V132(3) ,
    \V52(14) , \V64(1) , \V132(2) , \V64(2) ,
    \V167(4) , \V167(1) , \V167(0) , \V183(3) , \V183(2) , \V183(5) ,
    \V183(4) , \V167(7) , \V151(11) , \V167(6) , \V151(10) , \V199(11) ,
    \V167(9) , \V183(1) , \V151(13) , \V199(10) , \V167(8) , \V183(0) ,
    \V151(12) , \V199(13) , \V151(15) , \V199(12) , \V151(14) , \V199(15) ,
    \V199(14) , \V183(7) , \V183(6) , \V183(9) , \V183(8) , \V135(1) ,
    \V135(0) , \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) ,
    \V151(0) , \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V183(11) ,
    \V183(10) , \V183(13) , \V183(12) , \V167(11) , \V199(3) , \V183(15) ,
    \V167(10) , \V199(2) , \V183(14) , \V167(13) , \V199(5) , \V167(12) ,
    \V199(4) , \V167(15) , \V167(14) , \V199(1) , \V199(0) , \V199(7) ,
    \V199(6) , \V199(9) , \V199(8) , \V167(3) , \V167(2) , \V167(5)   );
  input  \V64(3) , \V28(13) , \V52(11) , \V52(10) , \V64(5) , \V28(15) ,
    \V109(3) , \V64(6) , \V28(14) , \V109(2) , \V132(1) , \V64(7) ,
    \V132(0) , \V64(9) , \V28(11) , \V115(3) , \V28(10) , \V115(2) ,
    \V88(1) , \V109(1) , \V16(1) , \V88(2) , \V121(3) , \V16(2) , \V88(3) ,
    \V121(2) , \V16(3) , \V64(13) , \V115(1) , \V88(5) , \V16(5) ,
    \V88(6) , \V16(6) , \V64(15) , \V88(7) , \V16(7) , \V64(14) ,
    \V121(1) , \V88(9) , \V16(9) , \V100(3) , \V100(2) , \V64(11) ,
    \V100(5) , \V64(10) , \V4(0) , \V100(1) , \V4(1) , \V118(3) ,
    \V118(2) , \V52(1) , \V52(2) , \V124(3) , \V52(3) , \V124(2) ,
    \V128(3) , \V100(7) , \V76(13) , \V128(2) , \V100(6) , \V118(1) ,
    \V52(5) , \V100(9) , \V76(15) , \V52(6) , \V76(14) , \V52(7) ,
    \V100(11) , \V124(1) , \V100(10) , \V52(9) , \V128(1) , \V103(3) ,
    \V100(13) , \V76(11) , \V128(0) , \V103(2) , \V76(10) , \V100(15) ,
    \V76(1) , \V100(14) , \V76(2) , \V76(3) , \V103(1) , \V76(5) ,
    \V76(6) , \V76(7) , \V76(9) , \V40(13) , \V88(13) , \V40(15) ,
    \V28(1) , \V40(14) , \V88(15) , \V28(2) , \V88(14) , \V28(3) ,
    \V16(13) , \V40(11) , \V28(5) , \V40(10) , \V16(15) , \V88(11) ,
    \V106(3) , \V28(6) , \V16(14) , \V88(10) , \V106(2) , \V28(7) ,
    \V40(1) , \V2(0) , \V133(0) , \V28(9) , \V40(2) , \V112(3) , \V16(11) ,
    \V2(1) , \V40(3) , \V112(2) , \V16(10) , \V106(1) , \V40(5) , \V40(6) ,
    \V40(7) , \V112(1) , \V52(13) , \V40(9) , \V52(15) , \V132(3) ,
    \V52(14) , \V64(1) , \V132(2) , \V64(2) ;
  output \V167(4) , \V167(1) , \V167(0) , \V183(3) , \V183(2) , \V183(5) ,
    \V183(4) , \V167(7) , \V151(11) , \V167(6) , \V151(10) , \V199(11) ,
    \V167(9) , \V183(1) , \V151(13) , \V199(10) , \V167(8) , \V183(0) ,
    \V151(12) , \V199(13) , \V151(15) , \V199(12) , \V151(14) , \V199(15) ,
    \V199(14) , \V183(7) , \V183(6) , \V183(9) , \V183(8) , \V135(1) ,
    \V135(0) , \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) ,
    \V151(0) , \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V183(11) ,
    \V183(10) , \V183(13) , \V183(12) , \V167(11) , \V199(3) , \V183(15) ,
    \V167(10) , \V199(2) , \V183(14) , \V167(13) , \V199(5) , \V167(12) ,
    \V199(4) , \V167(15) , \V167(14) , \V199(1) , \V199(0) , \V199(7) ,
    \V199(6) , \V199(9) , \V199(8) , \V167(3) , \V167(2) , \V167(5) ;
  wire n200, n202, n204, n206, n208, n210, n212, n214, n216, n218, n220,
    n222, n224, n226, n228, n230, n232, n234, n236, n238, n240, n242, n244,
    n246, n248, n250, n252, n254, n256, n258, n260, n262, n264, n266, n268,
    n270, n272, n274, n276, n278, n280, n282, n284, n286, n288, n290, n292,
    n294, n296, n298, n300, n302, n304, n306, n308, n310, n312, n314, n316,
    n318, n320, n322, n324, n326, n328, n330;
  assign n200 = \V133(0)  & \V132(3) ;
  assign \V199(0)  = \V128(3)  | n200;
  assign n202 = \V132(2)  & \V199(0) ;
  assign \V183(0)  = \V128(2)  | n202;
  assign n204 = \V112(3)  & \V183(0) ;
  assign \V167(12)  = \V109(3)  | n204;
  assign n206 = \V112(2)  & \V167(12) ;
  assign \V167(8)  = \V109(2)  | n206;
  assign n208 = \V112(1)  & \V167(8) ;
  assign \V167(4)  = \V109(1)  | n208;
  assign n210 = \V52(3)  & \V167(4) ;
  assign \V167(3)  = \V40(3)  | n210;
  assign n212 = \V52(2)  & \V167(3) ;
  assign \V167(2)  = \V40(2)  | n212;
  assign n214 = \V52(1)  & \V167(2) ;
  assign \V167(1)  = \V40(1)  | n214;
  assign n216 = \V132(1)  & \V183(0) ;
  assign \V167(0)  = \V128(1)  | n216;
  assign n218 = \V118(3)  & \V199(0) ;
  assign \V183(12)  = \V115(3)  | n218;
  assign n220 = \V118(2)  & \V183(12) ;
  assign \V183(8)  = \V115(2)  | n220;
  assign n222 = \V118(1)  & \V183(8) ;
  assign \V183(4)  = \V115(1)  | n222;
  assign n224 = \V76(3)  & \V183(4) ;
  assign \V183(3)  = \V64(3)  | n224;
  assign n226 = \V76(2)  & \V183(3) ;
  assign \V183(2)  = \V64(2)  | n226;
  assign n228 = \V76(7)  & \V183(8) ;
  assign \V183(7)  = \V64(7)  | n228;
  assign n230 = \V76(6)  & \V183(7) ;
  assign \V183(6)  = \V64(6)  | n230;
  assign n232 = \V76(5)  & \V183(6) ;
  assign \V183(5)  = \V64(5)  | n232;
  assign n234 = \V52(7)  & \V167(8) ;
  assign \V167(7)  = \V40(7)  | n234;
  assign n236 = \V106(3)  & \V167(0) ;
  assign \V151(12)  = \V103(3)  | n236;
  assign n238 = \V28(11)  & \V151(12) ;
  assign \V151(11)  = \V16(11)  | n238;
  assign n240 = \V52(6)  & \V167(7) ;
  assign \V167(6)  = \V40(6)  | n240;
  assign n242 = \V28(10)  & \V151(11) ;
  assign \V151(10)  = \V16(10)  | n242;
  assign n244 = \V124(3)  & \V133(0) ;
  assign \V199(12)  = \V121(3)  | n244;
  assign n246 = \V100(11)  & \V199(12) ;
  assign \V199(11)  = \V88(11)  | n246;
  assign n248 = \V52(11)  & \V167(12) ;
  assign \V167(11)  = \V40(11)  | n248;
  assign n250 = \V52(10)  & \V167(11) ;
  assign \V167(10)  = \V40(10)  | n250;
  assign n252 = \V52(9)  & \V167(10) ;
  assign \V167(9)  = \V40(9)  | n252;
  assign n254 = \V76(1)  & \V183(2) ;
  assign \V183(1)  = \V64(1)  | n254;
  assign n256 = \V28(15)  & \V167(0) ;
  assign \V151(15)  = \V16(15)  | n256;
  assign n258 = \V28(14)  & \V151(15) ;
  assign \V151(14)  = \V16(14)  | n258;
  assign n260 = \V28(13)  & \V151(14) ;
  assign \V151(13)  = \V16(13)  | n260;
  assign n262 = \V100(10)  & \V199(11) ;
  assign \V199(10)  = \V88(10)  | n262;
  assign n264 = \V100(15)  & \V133(0) ;
  assign \V199(15)  = \V88(15)  | n264;
  assign n266 = \V100(14)  & \V199(15) ;
  assign \V199(14)  = \V88(14)  | n266;
  assign n268 = \V100(13)  & \V199(14) ;
  assign \V199(13)  = \V88(13)  | n268;
  assign n270 = \V76(11)  & \V183(12) ;
  assign \V183(11)  = \V64(11)  | n270;
  assign n272 = \V76(10)  & \V183(11) ;
  assign \V183(10)  = \V64(10)  | n272;
  assign n274 = \V76(9)  & \V183(10) ;
  assign \V183(9)  = \V64(9)  | n274;
  assign n276 = \V132(0)  & \V167(0) ;
  assign \V151(0)  = \V128(0)  | n276;
  assign n278 = \V4(1)  & \V151(0) ;
  assign \V135(1)  = \V2(1)  | n278;
  assign n280 = \V4(0)  & \V135(1) ;
  assign \V135(0)  = \V2(0)  | n280;
  assign n282 = \V106(2)  & \V151(12) ;
  assign \V151(8)  = \V103(2)  | n282;
  assign n284 = \V106(1)  & \V151(8) ;
  assign \V151(4)  = \V103(1)  | n284;
  assign n286 = \V28(3)  & \V151(4) ;
  assign \V151(3)  = \V16(3)  | n286;
  assign n288 = \V28(2)  & \V151(3) ;
  assign \V151(2)  = \V16(2)  | n288;
  assign n290 = \V28(7)  & \V151(8) ;
  assign \V151(7)  = \V16(7)  | n290;
  assign n292 = \V28(6)  & \V151(7) ;
  assign \V151(6)  = \V16(6)  | n292;
  assign n294 = \V28(5)  & \V151(6) ;
  assign \V151(5)  = \V16(5)  | n294;
  assign n296 = \V28(1)  & \V151(2) ;
  assign \V151(1)  = \V16(1)  | n296;
  assign n298 = \V28(9)  & \V151(10) ;
  assign \V151(9)  = \V16(9)  | n298;
  assign n300 = \V76(15)  & \V199(0) ;
  assign \V183(15)  = \V64(15)  | n300;
  assign n302 = \V76(14)  & \V183(15) ;
  assign \V183(14)  = \V64(14)  | n302;
  assign n304 = \V76(13)  & \V183(14) ;
  assign \V183(13)  = \V64(13)  | n304;
  assign n306 = \V124(2)  & \V199(12) ;
  assign \V199(8)  = \V121(2)  | n306;
  assign n308 = \V124(1)  & \V199(8) ;
  assign \V199(4)  = \V121(1)  | n308;
  assign n310 = \V100(3)  & \V199(4) ;
  assign \V199(3)  = \V88(3)  | n310;
  assign n312 = \V100(2)  & \V199(3) ;
  assign \V199(2)  = \V88(2)  | n312;
  assign n314 = \V52(15)  & \V183(0) ;
  assign \V167(15)  = \V40(15)  | n314;
  assign n316 = \V52(14)  & \V167(15) ;
  assign \V167(14)  = \V40(14)  | n316;
  assign n318 = \V52(13)  & \V167(14) ;
  assign \V167(13)  = \V40(13)  | n318;
  assign n320 = \V100(7)  & \V199(8) ;
  assign \V199(7)  = \V88(7)  | n320;
  assign n322 = \V100(6)  & \V199(7) ;
  assign \V199(6)  = \V88(6)  | n322;
  assign n324 = \V100(5)  & \V199(6) ;
  assign \V199(5)  = \V88(5)  | n324;
  assign n326 = \V100(1)  & \V199(2) ;
  assign \V199(1)  = \V88(1)  | n326;
  assign n328 = \V100(9)  & \V199(10) ;
  assign \V199(9)  = \V88(9)  | n328;
  assign n330 = \V52(5)  & \V167(6) ;
  assign \V167(5)  = \V40(5)  | n330;
endmodule


