// Benchmark "f51m" written by ABC on Tue May 16 16:07:49 2017

module f51m ( 
    \1 , 2, 3, 4, 5, 6, 7, 8,
    44, 45, 46, 47, 48, 49, 50, 51  );
  input  \1 , 2, 3, 4, 5, 6, 7, 8;
  output 44, 45, 46, 47, 48, 49, 50, 51;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n247, n248, n249,
    n250, n251, n253, n254;
  assign n17 = ~\1  & ~2;
  assign n18 = 3 & n17;
  assign n19 = ~5 & n18;
  assign n20 = ~6 & n19;
  assign n21 = ~8 & n20;
  assign n22 = \1  & 2;
  assign n23 = 3 & n22;
  assign n24 = 6 & n23;
  assign n25 = 7 & n24;
  assign n26 = 8 & n25;
  assign n27 = ~\1  & 2;
  assign n28 = ~3 & n27;
  assign n29 = 5 & n28;
  assign n30 = 6 & n29;
  assign n31 = 8 & n30;
  assign n32 = ~7 & n20;
  assign n33 = 7 & n30;
  assign n34 = \1  & ~3;
  assign n35 = ~4 & n34;
  assign n36 = ~7 & n35;
  assign n37 = ~8 & n36;
  assign n38 = ~\1  & 3;
  assign n39 = ~4 & n38;
  assign n40 = ~5 & n39;
  assign n41 = ~8 & n40;
  assign n42 = \1  & 3;
  assign n43 = 4 & n42;
  assign n44 = 7 & n43;
  assign n45 = 8 & n44;
  assign n46 = \1  & ~2;
  assign n47 = ~3 & n46;
  assign n48 = ~6 & n47;
  assign n49 = ~7 & n48;
  assign n50 = ~7 & n40;
  assign n51 = ~\1  & ~3;
  assign n52 = 4 & n51;
  assign n53 = 5 & n52;
  assign n54 = 7 & n53;
  assign n55 = ~6 & n40;
  assign n56 = 6 & n53;
  assign n57 = ~6 & n35;
  assign n58 = 6 & n43;
  assign n59 = ~5 & n35;
  assign n60 = ~5 & n47;
  assign n61 = 5 & n43;
  assign n62 = 5 & n23;
  assign n63 = ~4 & n47;
  assign n64 = ~4 & n18;
  assign n65 = 4 & n28;
  assign n66 = 4 & n23;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~n64 & n67;
  assign n69 = ~n63 & n68;
  assign n70 = ~n62 & n69;
  assign n71 = ~n61 & n70;
  assign n72 = ~n60 & n71;
  assign n73 = ~n59 & n72;
  assign n74 = ~n58 & n73;
  assign n75 = ~n57 & n74;
  assign n76 = ~n56 & n75;
  assign n77 = ~n55 & n76;
  assign n78 = ~n54 & n77;
  assign n79 = ~n50 & n78;
  assign n80 = ~n49 & n79;
  assign n81 = ~n45 & n80;
  assign n82 = ~n41 & n81;
  assign n83 = ~n37 & n82;
  assign n84 = ~n33 & n83;
  assign n85 = ~n32 & n84;
  assign n86 = ~n31 & n85;
  assign n87 = ~n26 & n86;
  assign 44 = n21 | ~n87;
  assign n89 = 2 & 3;
  assign n90 = ~5 & n89;
  assign n91 = ~6 & n90;
  assign n92 = 7 & n91;
  assign n93 = 8 & n92;
  assign n94 = ~2 & 3;
  assign n95 = ~4 & n94;
  assign n96 = 6 & n95;
  assign n97 = 7 & n96;
  assign n98 = 8 & n97;
  assign n99 = 2 & ~3;
  assign n100 = ~4 & n99;
  assign n101 = ~7 & n100;
  assign n102 = ~8 & n101;
  assign n103 = ~2 & 4;
  assign n104 = ~5 & n103;
  assign n105 = ~6 & n104;
  assign n106 = ~8 & n105;
  assign n107 = ~2 & ~4;
  assign n108 = 5 & n107;
  assign n109 = 6 & n108;
  assign n110 = 8 & n109;
  assign n111 = ~7 & n105;
  assign n112 = ~2 & ~3;
  assign n113 = 4 & n112;
  assign n114 = ~6 & n113;
  assign n115 = ~7 & n114;
  assign n116 = 7 & n109;
  assign n117 = 2 & ~4;
  assign n118 = ~5 & n117;
  assign n119 = ~8 & n118;
  assign n120 = ~7 & n118;
  assign n121 = 2 & 4;
  assign n122 = 5 & n121;
  assign n123 = 7 & n122;
  assign n124 = ~6 & n100;
  assign n125 = 6 & n122;
  assign n126 = 4 & n89;
  assign n127 = 6 & n126;
  assign n128 = ~5 & n100;
  assign n129 = ~5 & n113;
  assign n130 = 5 & n95;
  assign n131 = 5 & n126;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~n129 & n132;
  assign n134 = ~n128 & n133;
  assign n135 = ~n127 & n134;
  assign n136 = ~n125 & n135;
  assign n137 = ~n124 & n136;
  assign n138 = ~n123 & n137;
  assign n139 = ~n120 & n138;
  assign n140 = ~n119 & n139;
  assign n141 = ~n116 & n140;
  assign n142 = ~n115 & n141;
  assign n143 = ~n111 & n142;
  assign n144 = ~n110 & n143;
  assign n145 = ~n106 & n144;
  assign n146 = ~n102 & n145;
  assign n147 = ~n98 & n146;
  assign 45 = n93 | ~n147;
  assign n149 = ~3 & ~4;
  assign n150 = 5 & n149;
  assign n151 = ~7 & n150;
  assign n152 = ~8 & n151;
  assign n153 = 3 & ~4;
  assign n154 = 6 & n153;
  assign n155 = ~7 & n154;
  assign n156 = 8 & n155;
  assign n157 = ~3 & ~5;
  assign n158 = 6 & n157;
  assign n159 = 7 & n158;
  assign n160 = 8 & n159;
  assign n161 = ~3 & 4;
  assign n162 = ~5 & n161;
  assign n163 = 7 & n162;
  assign n164 = 8 & n163;
  assign n165 = 3 & ~5;
  assign n166 = ~6 & n165;
  assign n167 = ~8 & n166;
  assign n168 = ~5 & n153;
  assign n169 = ~8 & n168;
  assign n170 = ~7 & n166;
  assign n171 = ~3 & 5;
  assign n172 = ~6 & n171;
  assign n173 = ~7 & n172;
  assign n174 = 3 & 5;
  assign n175 = 6 & n174;
  assign n176 = 7 & n175;
  assign n177 = 3 & 4;
  assign n178 = 5 & n177;
  assign n179 = 7 & n178;
  assign n180 = ~6 & n168;
  assign n181 = ~6 & n150;
  assign n182 = 6 & n162;
  assign n183 = 6 & n178;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~n181 & n184;
  assign n186 = ~n180 & n185;
  assign n187 = ~n179 & n186;
  assign n188 = ~n176 & n187;
  assign n189 = ~n173 & n188;
  assign n190 = ~n170 & n189;
  assign n191 = ~n169 & n190;
  assign n192 = ~n167 & n191;
  assign n193 = ~n164 & n192;
  assign n194 = ~n160 & n193;
  assign n195 = ~n156 & n194;
  assign 46 = n152 | ~n195;
  assign n197 = ~4 & 6;
  assign n198 = ~7 & n197;
  assign n199 = ~8 & n198;
  assign n200 = 4 & ~5;
  assign n201 = ~6 & n200;
  assign n202 = ~8 & n201;
  assign n203 = ~4 & ~5;
  assign n204 = 6 & n203;
  assign n205 = ~8 & n204;
  assign n206 = 4 & 5;
  assign n207 = ~7 & n206;
  assign n208 = 8 & n207;
  assign n209 = ~4 & ~6;
  assign n210 = 7 & n209;
  assign n211 = 8 & n210;
  assign n212 = 4 & 6;
  assign n213 = 7 & n212;
  assign n214 = 8 & n213;
  assign n215 = ~7 & n204;
  assign n216 = ~4 & 5;
  assign n217 = ~6 & n216;
  assign n218 = 7 & n217;
  assign n219 = 6 & n206;
  assign n220 = 7 & n219;
  assign n221 = 4 & ~6;
  assign n222 = ~7 & n221;
  assign n223 = ~n220 & ~n222;
  assign n224 = ~n218 & n223;
  assign n225 = ~n215 & n224;
  assign n226 = ~n214 & n225;
  assign n227 = ~n211 & n226;
  assign n228 = ~n208 & n227;
  assign n229 = ~n205 & n228;
  assign n230 = ~n202 & n229;
  assign 47 = n199 | ~n230;
  assign n232 = ~5 & 6;
  assign n233 = ~7 & n232;
  assign n234 = 8 & n233;
  assign n235 = 5 & ~7;
  assign n236 = ~8 & n235;
  assign n237 = ~5 & 7;
  assign n238 = ~8 & n237;
  assign n239 = 5 & ~6;
  assign n240 = ~7 & n239;
  assign n241 = 5 & 7;
  assign n242 = 8 & n241;
  assign n243 = ~n240 & ~n242;
  assign n244 = ~n238 & n243;
  assign n245 = ~n236 & n244;
  assign 48 = n234 | ~n245;
  assign n247 = ~6 & ~7;
  assign n248 = 8 & n247;
  assign n249 = 6 & ~8;
  assign n250 = 6 & 7;
  assign n251 = ~n249 & ~n250;
  assign 49 = n248 | ~n251;
  assign n253 = 7 & ~8;
  assign n254 = ~7 & 8;
  assign 50 = n253 | n254;
  assign 51 = ~8;
endmodule


