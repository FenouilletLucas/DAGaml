// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:57 2016

module TOP ( clock, 
    Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, Pi408, Pi407,
    Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, Pi398, Pi397,
    Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, Pi388, Pi387,
    Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, Pi378, Pi377,
    Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, Pi368, Pi367,
    Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, Pi358, Pi357,
    Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, Pi348, Pi347,
    Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, Pi338, Pi337,
    Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, Pi328, Pi327,
    Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, Pi318, Pi317,
    Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, Pi308, Pi307,
    Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, Pi298, Pi297,
    Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, Pi288, Pi287,
    Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, Pi278, Pi277,
    Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, Pi268, Pi267,
    Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, Pi258, Pi257,
    Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, Pi248, Pi247,
    Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, Pi238, Pi237,
    Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, Pi228, Pi227,
    Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, Pi218, Pi217,
    Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, Pi208, Pi207,
    Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, Pi198, Pi197,
    Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, Pi188, Pi187,
    Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, Pi178, Pi177,
    Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, Pi168, Pi167,
    Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, Pi158, Pi157,
    Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, Pi148, Pi147,
    Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, Pi138, Pi137,
    Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, Pi128, Pi127,
    Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, Pi118, Pi117,
    Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, Pi108, Pi107,
    Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, Pi98, Pi97,
    Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, Pi88, Pi87, Pi86, Pi85,
    Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, Pi78, Pi77, Pi76, Pi75, Pi74, Pi73,
    Pi72, Pi71, Pi70, Pi69, Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62, Pi61,
    Pi60, Pi59, Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50, Pi49,
    Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, Pi18, Pi17,
    Pi16, Pi15, PCLK,
    P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1, P__cmxcl_0,
    P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32, P__cmx1ad_31,
    P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27, P__cmx1ad_26,
    P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22, P__cmx1ad_21,
    P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17, P__cmx1ad_16,
    P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12, P__cmx1ad_11,
    P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7, P__cmx1ad_6,
    P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2, P__cmx1ad_1,
    P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33, P__cmx0ad_32,
    P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28, P__cmx0ad_27,
    P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23, P__cmx0ad_22,
    P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18, P__cmx0ad_17,
    P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13, P__cmx0ad_12,
    P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8, P__cmx0ad_7,
    P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3, P__cmx0ad_2,
    P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0, P__cmndst1p0,
    P__cmndst0p0  );
  input  clock;
  input  Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, Pi408,
    Pi407, Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, Pi398,
    Pi397, Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, Pi388,
    Pi387, Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, Pi378,
    Pi377, Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, Pi368,
    Pi367, Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, Pi358,
    Pi357, Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, Pi348,
    Pi347, Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, Pi338,
    Pi337, Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, Pi328,
    Pi327, Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, Pi318,
    Pi317, Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, Pi308,
    Pi307, Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, Pi298,
    Pi297, Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, Pi288,
    Pi287, Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, Pi278,
    Pi277, Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, Pi268,
    Pi267, Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, Pi258,
    Pi257, Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, Pi248,
    Pi247, Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, Pi238,
    Pi237, Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, Pi228,
    Pi227, Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, Pi218,
    Pi217, Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, Pi208,
    Pi207, Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, Pi198,
    Pi197, Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, Pi188,
    Pi187, Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, Pi178,
    Pi177, Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, Pi168,
    Pi167, Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, Pi158,
    Pi157, Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, Pi148,
    Pi147, Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, Pi138,
    Pi137, Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, Pi128,
    Pi127, Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, Pi118,
    Pi117, Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, Pi108,
    Pi107, Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, Pi98,
    Pi97, Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, Pi88, Pi87, Pi86,
    Pi85, Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, Pi78, Pi77, Pi76, Pi75, Pi74,
    Pi73, Pi72, Pi71, Pi70, Pi69, Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62,
    Pi61, Pi60, Pi59, Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50,
    Pi49, Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, Pi18,
    Pi17, Pi16, Pi15, PCLK;
  output P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1,
    P__cmxcl_0, P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32,
    P__cmx1ad_31, P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27,
    P__cmx1ad_26, P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22,
    P__cmx1ad_21, P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17,
    P__cmx1ad_16, P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12,
    P__cmx1ad_11, P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7,
    P__cmx1ad_6, P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2,
    P__cmx1ad_1, P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33,
    P__cmx0ad_32, P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28,
    P__cmx0ad_27, P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23,
    P__cmx0ad_22, P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18,
    P__cmx0ad_17, P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13,
    P__cmx0ad_12, P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8,
    P__cmx0ad_7, P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3,
    P__cmx0ad_2, P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0,
    P__cmndst1p0, P__cmndst0p0;
  reg Ni48, Ni47, Ni46, Ni45, Ni44, Ni43, Ni42, Ni41, Ni40, Ni39, Ni38,
    Ni37, Ni36, Ni35, Ni34, Ni33, Ni32, Ni31, Ni30, n18, Ni14, Ni13, Ni12,
    Ni11, Ni10, Ni9, Ni8, Ni7, Ni6, Ni5, Ni4, Ni3, Ni2;
  wire n568, n569, n570, n571, n574, n575, n576, n577, n578, n579, n580,
    n582, n583, n584, n602, n604, n616, n617, n635, n637, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n700, n701, n703,
    n704, n706, n707, n708, n709, n710, n711, n713, n714, n716, n717, n718,
    n719, n720, n721, n723, n724, n726, n727, n728, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n802, n803, n804, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932_1, n933,
    n934, n935, n936, n937_1, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962_1, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977_1, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992_1, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002_1, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012_1, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027_1, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042_1, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057_1, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072_1, n1073, n1074, n1075, n1076, n1077_1, n1078, n1079, n1080,
    n1081, n1082_1, n1083, n1084, n1085, n1086_1, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
    n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
    n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
    n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
    n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
    n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
    n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
    n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
    n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
    n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
    n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
    n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
    n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
    n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
    n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
    n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
    n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
    n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
    n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
    n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
    n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4995, n4996, n4997, n4998, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
    n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
    n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
    n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
    n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
    n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
    n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
    n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
    n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
    n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
    n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
    n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
    n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
    n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
    n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
    n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
    n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
    n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
    n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
    n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
    n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
    n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
    n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
    n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7949, n7950, n7951, n7952, n7954, n7955, n7956, n7957, n7958,
    n7959, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7981,
    n7982, n7983, n7984, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
    n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
    n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n932, n937, n942_1, n947_1, n952_1, n957_1,
    n962, n967_1, n972_1, n977, n982_1, n987_1, n992, n997_1, n1002,
    n1007_1, n1012, n1017_1, n1022_1, n1027, n1032_1, n1037_1, n1042,
    n1047_1, n1052_1, n1057, n1062_1, n1067_1, n1072, n1077, n1082, n1086,
    n1091_1;
  assign P__cmxig_1 = Ni33 & n18;
  assign P__cmxcl_1 = ~Ni3 & ~Ni2;
  assign n568 = ~Ni13 & ~Ni11;
  assign n569 = ~Ni12 & n568;
  assign n570 = Ni14 & n569;
  assign n571 = P__cmxcl_1 & n570;
  assign P__cmxir_1 = ~P__cmxig_1 & n571;
  assign P__cmxig_0 = ~Ni33 & n18;
  assign n574 = Ni10 & ~P__cmxig_0;
  assign n575 = Pi25 & ~Ni10;
  assign n576 = ~Ni9 & ~n575;
  assign n577 = ~n574 & n576;
  assign n578 = ~Ni8 & ~Ni7;
  assign n579 = ~Ni9 & n578;
  assign n580 = P__cmxcl_1 & n579;
  assign P__cmxir_0 = ~n577 & n580;
  assign n582 = ~Ni12 & ~Ni11;
  assign n583 = Ni14 & Ni13;
  assign n584 = n582 & n583;
  assign P__cmx1ad_9 = P__cmxcl_1 & n584;
  assign P__cmx1ad_31 = Pi255 & P__cmx1ad_9;
  assign P__cmx1ad_30 = Pi254 & P__cmx1ad_9;
  assign P__cmx1ad_29 = Pi253 & P__cmx1ad_9;
  assign P__cmx1ad_28 = Pi252 & P__cmx1ad_9;
  assign P__cmx1ad_27 = Pi251 & P__cmx1ad_9;
  assign P__cmx1ad_26 = Pi250 & P__cmx1ad_9;
  assign P__cmx1ad_25 = Pi249 & P__cmx1ad_9;
  assign P__cmx1ad_24 = Pi248 & P__cmx1ad_9;
  assign P__cmx1ad_23 = Pi247 & P__cmx1ad_9;
  assign P__cmx1ad_22 = Pi246 & P__cmx1ad_9;
  assign P__cmx1ad_21 = Pi245 & P__cmx1ad_9;
  assign P__cmx1ad_20 = Pi244 & P__cmx1ad_9;
  assign P__cmx1ad_19 = Pi243 & P__cmx1ad_9;
  assign P__cmx1ad_18 = Pi242 & P__cmx1ad_9;
  assign P__cmx1ad_17 = Pi241 & P__cmx1ad_9;
  assign P__cmx1ad_16 = Pi240 & P__cmx1ad_9;
  assign n602 = Pi27 & Pi26;
  assign P__cmx1ad_15 = P__cmx1ad_9 & n602;
  assign n604 = ~Pi27 & ~Pi26;
  assign P__cmx1ad_13 = P__cmx1ad_9 & ~n604;
  assign P__cmx1ad_14 = ~n602 & P__cmx1ad_13;
  assign P__cmx1ad_12 = ~Pi27 & P__cmx1ad_9;
  assign P__cmx1ad_7 = Pi239 & P__cmx1ad_9;
  assign P__cmx1ad_6 = Pi238 & P__cmx1ad_9;
  assign P__cmx1ad_5 = Pi237 & P__cmx1ad_9;
  assign P__cmx1ad_4 = Pi236 & P__cmx1ad_9;
  assign P__cmx1ad_3 = Pi235 & P__cmx1ad_9;
  assign P__cmx1ad_2 = Pi234 & P__cmx1ad_9;
  assign P__cmx1ad_1 = Pi233 & P__cmx1ad_9;
  assign P__cmx1ad_0 = Pi232 & P__cmx1ad_9;
  assign n616 = Ni10 & Ni9;
  assign n617 = n578 & n616;
  assign P__cmx0ad_9 = P__cmxcl_1 & n617;
  assign P__cmx0ad_31 = Pi72 & P__cmx0ad_9;
  assign P__cmx0ad_30 = Pi71 & P__cmx0ad_9;
  assign P__cmx0ad_29 = Pi70 & P__cmx0ad_9;
  assign P__cmx0ad_28 = Pi69 & P__cmx0ad_9;
  assign P__cmx0ad_27 = Pi68 & P__cmx0ad_9;
  assign P__cmx0ad_26 = Pi67 & P__cmx0ad_9;
  assign P__cmx0ad_25 = Pi66 & P__cmx0ad_9;
  assign P__cmx0ad_24 = Pi65 & P__cmx0ad_9;
  assign P__cmx0ad_23 = Pi64 & P__cmx0ad_9;
  assign P__cmx0ad_22 = Pi63 & P__cmx0ad_9;
  assign P__cmx0ad_21 = Pi62 & P__cmx0ad_9;
  assign P__cmx0ad_20 = Pi61 & P__cmx0ad_9;
  assign P__cmx0ad_19 = Pi60 & P__cmx0ad_9;
  assign P__cmx0ad_18 = Pi59 & P__cmx0ad_9;
  assign P__cmx0ad_17 = Pi58 & P__cmx0ad_9;
  assign P__cmx0ad_16 = Pi57 & P__cmx0ad_9;
  assign n635 = Pi24 & Pi23;
  assign P__cmx0ad_15 = P__cmx0ad_9 & n635;
  assign n637 = ~Pi24 & ~Pi23;
  assign P__cmx0ad_13 = P__cmx0ad_9 & ~n637;
  assign P__cmx0ad_14 = ~n635 & P__cmx0ad_13;
  assign P__cmx0ad_12 = ~Pi24 & P__cmx0ad_9;
  assign P__cmx0ad_7 = Pi56 & P__cmx0ad_9;
  assign P__cmx0ad_6 = Pi55 & P__cmx0ad_9;
  assign P__cmx0ad_5 = Pi54 & P__cmx0ad_9;
  assign P__cmx0ad_4 = Pi53 & P__cmx0ad_9;
  assign P__cmx0ad_3 = Pi52 & P__cmx0ad_9;
  assign P__cmx0ad_2 = Pi51 & P__cmx0ad_9;
  assign P__cmx0ad_1 = Pi50 & P__cmx0ad_9;
  assign P__cmx0ad_0 = Pi49 & P__cmx0ad_9;
  assign n1091_1 = Ni3 & ~Ni2;
  assign n650 = ~Ni4 & n1091_1;
  assign n651 = Ni5 & n650;
  assign n652 = Ni31 & Ni30;
  assign n653 = ~Ni36 & ~Ni32;
  assign n654 = ~Ni41 & Ni32;
  assign n655 = ~n653 & ~n654;
  assign n656 = n652 & ~n655;
  assign n657 = n651 & n656;
  assign n658 = ~Ni6 & n657;
  assign n659 = Ni31 & ~Ni30;
  assign n660 = Ni6 & ~Ni5;
  assign n661 = n650 & n660;
  assign n662 = n659 & n661;
  assign n663 = n652 & n655;
  assign n664 = Ni4 & n1091_1;
  assign n665 = n660 & n664;
  assign n666 = n663 & n665;
  assign n667 = ~n662 & ~n666;
  assign n668 = ~n658 & n667;
  assign n669 = Ni33 & ~n668;
  assign n670 = Ni12 & ~Ni11;
  assign n671 = ~Ni13 & n670;
  assign n672 = ~Ni14 & ~n604;
  assign n673 = n671 & ~n672;
  assign n674 = ~Pi27 & Ni14;
  assign n675 = P__cmxcl_1 & ~n674;
  assign n676 = n673 & n675;
  assign n677 = ~Pi27 & Pi26;
  assign n678 = Ni14 & ~Ni13;
  assign n679 = ~Ni12 & n678;
  assign n680 = Ni11 & n679;
  assign n681 = n677 & n680;
  assign n682 = P__cmxcl_1 & n681;
  assign n683 = ~n676 & ~n682;
  assign P__cmnxcp_1 = n669 | ~n683;
  assign n685 = ~Pi24 & Ni10;
  assign n686 = ~Ni9 & ~Ni7;
  assign n687 = ~Ni10 & ~n637;
  assign n688 = n686 & ~n687;
  assign n689 = ~n685 & n688;
  assign n690 = Ni8 & n689;
  assign n691 = ~Pi24 & Pi23;
  assign n692 = Ni10 & ~Ni8;
  assign n693 = ~Ni9 & n692;
  assign n694 = Ni7 & n693;
  assign n695 = n691 & n694;
  assign n696 = ~n690 & ~n695;
  assign n697 = P__cmxcl_1 & ~n696;
  assign n698 = ~Ni33 & ~n668;
  assign P__cmnxcp_0 = n697 | n698;
  assign n700 = Ni32 & Ni30;
  assign n701 = Ni43 & ~n700;
  assign P__cmndst1p0 = ~Ni42 & n701;
  assign n703 = ~Ni32 & Ni30;
  assign n704 = Ni38 & ~Ni37;
  assign P__cmndst0p0 = ~n703 & n704;
  assign n706 = Ni32 & ~Ni30;
  assign n707 = Ni31 & n706;
  assign n708 = ~Pi22 & ~n707;
  assign n709 = ~Ni47 & n708;
  assign n710 = Pi20 & n709;
  assign n711 = Ni48 & ~n709;
  assign n932 = n710 | n711;
  assign n713 = Ni32 & n662;
  assign n714 = Ni47 & ~n713;
  assign n937 = n708 | n714;
  assign n716 = ~Pi21 & Ni32;
  assign n717 = ~Pi21 & ~n659;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~Ni45 & ~n718;
  assign n720 = Pi20 & n719;
  assign n721 = Ni46 & ~n719;
  assign n942_1 = n720 | n721;
  assign n723 = ~Ni32 & n662;
  assign n724 = Ni45 & ~n723;
  assign n947_1 = ~n718 | n724;
  assign n726 = ~Ni31 & n700;
  assign n727 = ~Ni33 & n726;
  assign n728 = ~Ni44 & ~n726;
  assign n952_1 = ~n727 & ~n728;
  assign n730 = Pi19 & Pi17;
  assign n731 = ~Pi16 & n730;
  assign n732 = ~Pi20 & ~Ni44;
  assign n733 = Pi20 & Ni44;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n731 & ~n734;
  assign n736 = ~Pi19 & Pi17;
  assign n737 = Ni40 & n736;
  assign n738 = Pi19 & ~Pi17;
  assign n739 = ~Ni40 & n738;
  assign n740 = ~n737 & ~n739;
  assign n741 = n735 & n740;
  assign n742 = ~Ni41 & ~n741;
  assign n743 = Pi16 & Ni41;
  assign n744 = Pi16 & n730;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n742 & n745;
  assign n747 = ~Ni42 & n746;
  assign n748 = n701 & ~n747;
  assign n957_1 = n726 | n748;
  assign n750 = ~Ni38 & ~Ni37;
  assign n751 = ~n703 & n750;
  assign n752 = ~Ni44 & ~Ni39;
  assign n753 = Ni44 & Ni39;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n751 & ~n754;
  assign n756 = Ni43 & Ni42;
  assign n757 = ~n700 & ~n756;
  assign n758 = ~n755 & ~n757;
  assign n759 = Pi18 & ~Pi17;
  assign n760 = Ni40 & n759;
  assign n761 = ~n734 & n760;
  assign n762 = ~Ni41 & ~n761;
  assign n763 = Ni43 & ~n743;
  assign n764 = ~n762 & n763;
  assign n765 = ~Ni42 & ~n764;
  assign n766 = ~n700 & ~n765;
  assign n767 = ~n726 & ~n766;
  assign n962 = ~n758 & ~n767;
  assign n769 = ~Pi27 & Ni33;
  assign n770 = n584 & n769;
  assign n771 = ~Pi24 & ~Ni33;
  assign n772 = n617 & n771;
  assign n773 = ~n770 & ~n772;
  assign n774 = ~Ni6 & ~Ni4;
  assign n775 = ~Ni5 & n774;
  assign n776 = P__cmxcl_1 & n775;
  assign n777 = n726 & n776;
  assign n778 = ~n773 & n777;
  assign n779 = ~Ni33 & ~n617;
  assign n780 = Ni33 & ~n584;
  assign n781 = ~n779 & ~n780;
  assign n782 = n777 & n781;
  assign n783 = ~Ni41 & ~n782;
  assign n967_1 = ~n778 & ~n783;
  assign n785 = Ni40 & ~n726;
  assign n786 = Pi23 & n776;
  assign n787 = n727 & n786;
  assign n788 = ~n785 & ~n787;
  assign n789 = n617 & ~n788;
  assign n790 = Ni33 & n726;
  assign n791 = Pi26 & n775;
  assign n792 = P__cmx1ad_9 & n791;
  assign n793 = Ni40 & ~n584;
  assign n794 = ~n792 & ~n793;
  assign n795 = n790 & ~n794;
  assign n796 = P__cmx0ad_9 & n775;
  assign n797 = n776 & n790;
  assign n798 = Ni40 & ~n797;
  assign n799 = ~n796 & n798;
  assign n800 = ~n795 & ~n799;
  assign n972_1 = n789 | ~n800;
  assign n802 = ~Ni31 & n703;
  assign n803 = ~Ni33 & n802;
  assign n804 = ~Ni39 & ~n802;
  assign n977 = ~n803 & ~n804;
  assign n806 = ~Pi20 & ~Ni39;
  assign n807 = Pi20 & Ni39;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~Ni37 & ~Ni36;
  assign n810 = ~Pi19 & ~Ni35;
  assign n811 = ~Pi17 & Ni35;
  assign n812 = ~n810 & ~n811;
  assign n813 = n809 & ~n812;
  assign n814 = ~n808 & n813;
  assign n815 = Ni38 & ~n703;
  assign n816 = ~Ni37 & Ni36;
  assign n817 = ~Pi15 & n816;
  assign n818 = n815 & ~n817;
  assign n819 = ~n814 & n818;
  assign n982_1 = n802 | n819;
  assign n821 = ~Ni37 & n759;
  assign n822 = ~Ni36 & Ni35;
  assign n823 = ~n808 & n822;
  assign n824 = n821 & n823;
  assign n825 = ~n817 & ~n824;
  assign n826 = n815 & ~n825;
  assign n827 = ~Ni43 & ~Ni42;
  assign n828 = ~Ni30 & n827;
  assign n829 = ~n754 & ~n828;
  assign n830 = Ni38 & ~n829;
  assign n831 = Ni37 & ~n703;
  assign n832 = ~n754 & n802;
  assign n833 = ~n827 & n832;
  assign n834 = ~n831 & ~n833;
  assign n835 = ~n830 & ~n834;
  assign n987_1 = n826 | n835;
  assign n837 = Ni33 & n802;
  assign n838 = n617 & ~n837;
  assign n839 = ~n584 & ~n838;
  assign n840 = n776 & n802;
  assign n841 = ~n779 & n840;
  assign n842 = ~n839 & n841;
  assign n843 = Ni36 & ~n842;
  assign n844 = ~n771 & ~n780;
  assign n845 = n841 & n844;
  assign n846 = ~n769 & n845;
  assign n992 = n843 | n846;
  assign n848 = n792 & n837;
  assign n849 = n584 & ~n803;
  assign n850 = ~n617 & ~n849;
  assign n851 = n840 & ~n850;
  assign n852 = Ni35 & ~n851;
  assign n853 = Pi23 & n803;
  assign n854 = Ni33 & Ni30;
  assign n855 = ~Ni31 & n854;
  assign n856 = Ni35 & ~Ni32;
  assign n857 = n855 & n856;
  assign n858 = ~n584 & n857;
  assign n859 = ~n853 & ~n858;
  assign n860 = n796 & ~n859;
  assign n861 = ~n852 & ~n860;
  assign n997_1 = n848 | ~n861;
  assign n863 = ~Ni10 & ~n570;
  assign n864 = Pi22 & Pi21;
  assign n865 = Pi25 & n864;
  assign n866 = Ni34 & ~n865;
  assign n867 = ~Pi20 & n864;
  assign n868 = Pi25 & n867;
  assign n869 = ~Pi16 & n736;
  assign n870 = ~Ni31 & ~Ni30;
  assign n871 = ~Ni32 & n870;
  assign n872 = ~Ni47 & ~Ni45;
  assign n873 = ~Ni38 & Ni37;
  assign n874 = ~Ni43 & Ni42;
  assign n875 = ~n873 & ~n874;
  assign n876 = n872 & n875;
  assign n877 = ~Ni47 & n827;
  assign n878 = ~Ni41 & n877;
  assign n879 = ~Ni45 & n878;
  assign n880 = ~Ni43 & n872;
  assign n881 = Ni44 & n880;
  assign n882 = ~Ni40 & ~n881;
  assign n883 = n879 & ~n882;
  assign n884 = Ni38 & ~n883;
  assign n885 = n876 & ~n884;
  assign n886 = n822 & ~n885;
  assign n887 = n872 & ~n874;
  assign n888 = ~Ni35 & ~n887;
  assign n889 = ~Ni36 & n704;
  assign n890 = ~Ni39 & ~Ni36;
  assign n891 = ~Ni37 & n890;
  assign n892 = ~n889 & ~n891;
  assign n893 = ~Ni35 & ~n892;
  assign n894 = ~n883 & n893;
  assign n895 = ~n888 & ~n894;
  assign n896 = ~n809 & ~n883;
  assign n897 = ~n873 & ~n896;
  assign n898 = n895 & n897;
  assign n899 = ~n886 & n898;
  assign n900 = n871 & n899;
  assign n901 = ~Ni34 & ~n900;
  assign n902 = n869 & ~n901;
  assign n903 = ~Pi16 & n738;
  assign n904 = Ni40 & ~n881;
  assign n905 = n879 & ~n904;
  assign n906 = Ni38 & ~n905;
  assign n907 = n876 & ~n906;
  assign n908 = ~Ni36 & ~Ni35;
  assign n909 = ~n907 & n908;
  assign n910 = Ni35 & ~n887;
  assign n911 = Ni35 & ~n892;
  assign n912 = ~n905 & n911;
  assign n913 = ~n910 & ~n912;
  assign n914 = ~n809 & ~n905;
  assign n915 = ~n873 & ~n914;
  assign n916 = n913 & n915;
  assign n917 = ~n909 & n916;
  assign n918 = n871 & n917;
  assign n919 = ~Ni34 & ~n918;
  assign n920 = n903 & ~n919;
  assign n921 = ~n902 & ~n920;
  assign n922 = n868 & ~n921;
  assign n923 = ~Pi19 & ~Pi17;
  assign n924 = Pi16 & n923;
  assign n925 = ~n750 & ~n816;
  assign n926 = ~n890 & ~n925;
  assign n927 = ~Ni44 & ~Ni41;
  assign n928 = ~Ni45 & n827;
  assign n929 = ~n927 & n928;
  assign n930 = ~Ni47 & n929;
  assign n931 = ~n926 & ~n930;
  assign n932_1 = n876 & ~n931;
  assign n933 = n816 & ~n930;
  assign n934 = n932_1 & ~n933;
  assign n935 = n871 & n934;
  assign n936 = ~Ni34 & ~n935;
  assign n937_1 = n868 & ~n936;
  assign n938 = Ni39 & n809;
  assign n939 = ~n925 & ~n938;
  assign n940 = Ni44 & ~Ni41;
  assign n941 = n928 & ~n940;
  assign n942 = ~Ni47 & n941;
  assign n943 = ~n939 & ~n942;
  assign n944 = n876 & ~n943;
  assign n945 = n816 & ~n942;
  assign n946 = n944 & ~n945;
  assign n947 = n871 & n946;
  assign n948 = ~Ni34 & ~n947;
  assign n949 = Pi20 & n864;
  assign n950 = Pi25 & n949;
  assign n951 = ~n948 & n950;
  assign n952 = ~n937_1 & ~n951;
  assign n953 = n924 & ~n952;
  assign n954 = ~n922 & ~n953;
  assign n955 = Pi16 & n738;
  assign n956 = ~Ni44 & Ni40;
  assign n957 = ~Ni41 & n956;
  assign n958 = n928 & ~n957;
  assign n959 = ~Ni47 & n958;
  assign n960 = Ni38 & ~n959;
  assign n961 = n876 & ~n960;
  assign n962_1 = n908 & ~n961;
  assign n963 = n911 & ~n959;
  assign n964 = ~n910 & ~n963;
  assign n965 = ~n873 & n958;
  assign n966 = ~Ni47 & n965;
  assign n967 = ~n809 & ~n966;
  assign n968 = n964 & ~n967;
  assign n969 = ~n962_1 & n968;
  assign n970 = n871 & n969;
  assign n971 = ~Ni34 & ~n970;
  assign n972 = n868 & ~n971;
  assign n973 = Ni44 & Ni40;
  assign n974 = ~Ni41 & n973;
  assign n975 = n928 & ~n974;
  assign n976 = ~Ni47 & n975;
  assign n977_1 = Ni38 & ~n976;
  assign n978 = n876 & ~n977_1;
  assign n979 = n908 & ~n978;
  assign n980 = ~n889 & ~n938;
  assign n981 = Ni35 & ~n980;
  assign n982 = ~n976 & n981;
  assign n983 = ~n910 & ~n982;
  assign n984 = ~n873 & n975;
  assign n985 = ~Ni47 & n984;
  assign n986 = ~n809 & ~n985;
  assign n987 = n983 & ~n986;
  assign n988 = ~n979 & n987;
  assign n989 = n871 & n988;
  assign n990 = ~Ni34 & ~n989;
  assign n991 = n950 & ~n990;
  assign n992_1 = ~n972 & ~n991;
  assign n993 = n955 & ~n992_1;
  assign n994 = ~Pi16 & n923;
  assign n995 = ~Ni41 & n928;
  assign n996 = Ni44 & n995;
  assign n997 = ~Ni47 & n996;
  assign n998 = ~n926 & ~n997;
  assign n999 = n876 & ~n998;
  assign n1000 = n816 & ~n997;
  assign n1001 = n999 & ~n1000;
  assign n1002_1 = n871 & n1001;
  assign n1003 = ~Ni34 & ~n1002_1;
  assign n1004 = n868 & ~n1003;
  assign n1005 = ~Ni42 & n927;
  assign n1006 = n880 & n1005;
  assign n1007 = ~n939 & ~n1006;
  assign n1008 = n876 & ~n1007;
  assign n1009 = n816 & ~n1006;
  assign n1010 = n1008 & ~n1009;
  assign n1011 = n871 & n1010;
  assign n1012_1 = ~Ni34 & ~n1011;
  assign n1013 = n950 & ~n1012_1;
  assign n1014 = ~n1004 & ~n1013;
  assign n1015 = n994 & ~n1014;
  assign n1016 = Ni38 & ~n879;
  assign n1017 = n876 & ~n1016;
  assign n1018 = Ni36 & ~n879;
  assign n1019 = n1017 & ~n1018;
  assign n1020 = n871 & n1019;
  assign n1021 = ~Ni34 & ~n1020;
  assign n1022 = ~Pi16 & n1021;
  assign n1023 = ~Ni47 & n928;
  assign n1024 = Ni38 & ~n1023;
  assign n1025 = n876 & ~n1024;
  assign n1026 = Ni36 & ~n1023;
  assign n1027_1 = n1025 & ~n1026;
  assign n1028 = n871 & n1027_1;
  assign n1029 = ~Ni34 & ~n1028;
  assign n1030 = n730 & n864;
  assign n1031 = Pi25 & n1030;
  assign n1032 = ~n1029 & n1031;
  assign n1033 = ~n1022 & n1032;
  assign n1034 = ~n1015 & ~n1033;
  assign n1035 = Pi16 & n736;
  assign n1036 = ~Ni44 & ~Ni40;
  assign n1037 = ~Ni41 & n1036;
  assign n1038 = n928 & ~n1037;
  assign n1039 = ~Ni47 & n1038;
  assign n1040 = Ni38 & ~n1039;
  assign n1041 = n876 & ~n1040;
  assign n1042_1 = n822 & ~n1041;
  assign n1043 = n893 & ~n1039;
  assign n1044 = ~n888 & ~n1043;
  assign n1045 = ~n873 & n1038;
  assign n1046 = ~Ni47 & n1045;
  assign n1047 = ~n809 & ~n1046;
  assign n1048 = n1044 & ~n1047;
  assign n1049 = ~n1042_1 & n1048;
  assign n1050 = n871 & n1049;
  assign n1051 = ~Ni34 & ~n1050;
  assign n1052 = n868 & ~n1051;
  assign n1053 = Ni44 & ~Ni40;
  assign n1054 = ~Ni41 & n1053;
  assign n1055 = n928 & ~n1054;
  assign n1056 = ~Ni47 & n1055;
  assign n1057_1 = Ni38 & ~n1056;
  assign n1058 = n876 & ~n1057_1;
  assign n1059 = n822 & ~n1058;
  assign n1060 = ~Ni35 & ~n980;
  assign n1061 = ~n1056 & n1060;
  assign n1062 = ~n888 & ~n1061;
  assign n1063 = ~n873 & n1055;
  assign n1064 = ~Ni47 & n1063;
  assign n1065 = ~n809 & ~n1064;
  assign n1066 = n1062 & ~n1065;
  assign n1067 = ~n1059 & n1066;
  assign n1068 = n871 & n1067;
  assign n1069 = ~Ni34 & ~n1068;
  assign n1070 = n950 & ~n1069;
  assign n1071 = ~n1052 & ~n1070;
  assign n1072_1 = n1035 & ~n1071;
  assign n1073 = n1034 & ~n1072_1;
  assign n1074 = ~n993 & n1073;
  assign n1075 = ~Ni44 & n880;
  assign n1076 = ~Ni40 & ~n1075;
  assign n1077_1 = n879 & ~n1076;
  assign n1078 = Ni38 & ~n1077_1;
  assign n1079 = n876 & ~n1078;
  assign n1080 = n822 & ~n1079;
  assign n1081 = n1060 & ~n1077_1;
  assign n1082_1 = ~n888 & ~n1081;
  assign n1083 = ~n809 & ~n1077_1;
  assign n1084 = ~n873 & ~n1083;
  assign n1085 = n1082_1 & n1084;
  assign n1086_1 = ~n1080 & n1085;
  assign n1087 = n871 & n1086_1;
  assign n1088 = ~Ni34 & ~n1087;
  assign n1089 = n869 & ~n1088;
  assign n1090 = Ni40 & ~n1075;
  assign n1091 = n879 & ~n1090;
  assign n1092 = Ni38 & ~n1091;
  assign n1093 = n876 & ~n1092;
  assign n1094 = n908 & ~n1093;
  assign n1095 = n981 & ~n1091;
  assign n1096 = ~n910 & ~n1095;
  assign n1097 = ~n809 & ~n1091;
  assign n1098 = ~n873 & ~n1097;
  assign n1099 = n1096 & n1098;
  assign n1100 = ~n1094 & n1099;
  assign n1101 = n871 & n1100;
  assign n1102 = ~Ni34 & ~n1101;
  assign n1103 = n903 & ~n1102;
  assign n1104 = ~n1089 & ~n1103;
  assign n1105 = n950 & ~n1104;
  assign n1106 = ~Pi15 & ~n1105;
  assign n1107 = n1074 & n1106;
  assign n1108 = n954 & n1107;
  assign n1109 = ~Ni38 & n999;
  assign n1110 = ~n1001 & ~n1109;
  assign n1111 = n871 & ~n1110;
  assign n1112 = ~Ni34 & ~n1111;
  assign n1113 = n868 & ~n1112;
  assign n1114 = ~Ni38 & n1008;
  assign n1115 = ~n1010 & ~n1114;
  assign n1116 = n871 & ~n1115;
  assign n1117 = ~Ni34 & ~n1116;
  assign n1118 = n950 & ~n1117;
  assign n1119 = ~n1113 & ~n1118;
  assign n1120 = n994 & ~n1119;
  assign n1121 = n907 & n913;
  assign n1122 = n871 & n1121;
  assign n1123 = ~Ni34 & ~n1122;
  assign n1124 = n903 & ~n1123;
  assign n1125 = n885 & n895;
  assign n1126 = n871 & n1125;
  assign n1127 = ~Ni34 & ~n1126;
  assign n1128 = n869 & ~n1127;
  assign n1129 = ~n1124 & ~n1128;
  assign n1130 = Ni38 & n933;
  assign n1131 = n932_1 & ~n1130;
  assign n1132 = n871 & n1131;
  assign n1133 = ~Ni34 & ~n1132;
  assign n1134 = n924 & ~n1133;
  assign n1135 = n1129 & ~n1134;
  assign n1136 = n868 & ~n1135;
  assign n1137 = n1079 & n1082_1;
  assign n1138 = n871 & n1137;
  assign n1139 = ~Ni34 & ~n1138;
  assign n1140 = n869 & ~n1139;
  assign n1141 = n1093 & n1096;
  assign n1142 = n871 & n1141;
  assign n1143 = ~Ni34 & ~n1142;
  assign n1144 = n903 & ~n1143;
  assign n1145 = ~Ni38 & n944;
  assign n1146 = ~n946 & ~n1145;
  assign n1147 = n871 & ~n1146;
  assign n1148 = ~Ni34 & ~n1147;
  assign n1149 = n924 & ~n1148;
  assign n1150 = ~n1144 & ~n1149;
  assign n1151 = ~n1140 & n1150;
  assign n1152 = n950 & ~n1151;
  assign n1153 = ~n1136 & ~n1152;
  assign n1154 = n961 & n964;
  assign n1155 = n871 & n1154;
  assign n1156 = ~Ni34 & ~n1155;
  assign n1157 = n868 & ~n1156;
  assign n1158 = n978 & n983;
  assign n1159 = n871 & n1158;
  assign n1160 = ~Ni34 & ~n1159;
  assign n1161 = n950 & ~n1160;
  assign n1162 = ~n1157 & ~n1161;
  assign n1163 = n955 & ~n1162;
  assign n1164 = n1041 & n1044;
  assign n1165 = n871 & n1164;
  assign n1166 = ~Ni34 & ~n1165;
  assign n1167 = n868 & ~n1166;
  assign n1168 = n1058 & n1062;
  assign n1169 = n871 & n1168;
  assign n1170 = ~Ni34 & ~n1169;
  assign n1171 = n950 & ~n1170;
  assign n1172 = ~n1167 & ~n1171;
  assign n1173 = n1035 & ~n1172;
  assign n1174 = n871 & n1025;
  assign n1175 = ~Ni34 & ~n1174;
  assign n1176 = n1031 & ~n1175;
  assign n1177 = Pi15 & ~n1176;
  assign n1178 = ~Pi16 & Pi15;
  assign n1179 = n871 & n1017;
  assign n1180 = ~Ni34 & ~n1179;
  assign n1181 = n1178 & n1180;
  assign n1182 = ~n1177 & ~n1181;
  assign n1183 = ~n1173 & ~n1182;
  assign n1184 = ~n1163 & n1183;
  assign n1185 = n1153 & n1184;
  assign n1186 = ~n1120 & n1185;
  assign n1187 = ~n1108 & ~n1186;
  assign n1188 = ~n866 & ~n1187;
  assign n1189 = n863 & ~n1188;
  assign n1190 = ~Pi15 & n570;
  assign n1191 = ~n18 & n864;
  assign n1192 = ~n1051 & n1191;
  assign n1193 = Ni34 & n1049;
  assign n1194 = n1192 & ~n1193;
  assign n1195 = n864 & n871;
  assign n1196 = Ni34 & ~n1195;
  assign n1197 = Ni34 & P__cmxig_0;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = n18 & n1195;
  assign n1200 = ~Ni34 & ~n1049;
  assign n1201 = Ni33 & ~n1200;
  assign n1202 = n1199 & n1201;
  assign n1203 = n1198 & ~n1202;
  assign n1204 = n1049 & ~n1202;
  assign n1205 = ~n1196 & n1204;
  assign n1206 = ~n1203 & ~n1205;
  assign n1207 = ~n1194 & ~n1206;
  assign n1208 = n1035 & ~n1207;
  assign n1209 = ~n971 & n1191;
  assign n1210 = Ni34 & Ni33;
  assign n1211 = Ni33 & n969;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = n1199 & ~n1212;
  assign n1214 = n1198 & ~n1213;
  assign n1215 = ~n1209 & n1214;
  assign n1216 = n955 & ~n1215;
  assign n1217 = ~Ni34 & n871;
  assign n1218 = n1191 & n1217;
  assign n1219 = ~n1196 & ~n1218;
  assign n1220 = n969 & ~n1213;
  assign n1221 = n1219 & n1220;
  assign n1222 = n1216 & ~n1221;
  assign n1223 = ~Ni34 & ~n934;
  assign n1224 = Ni33 & ~n1223;
  assign n1225 = n1199 & n1224;
  assign n1226 = ~n1196 & ~n1225;
  assign n1227 = ~n1191 & ~n1197;
  assign n1228 = ~n936 & ~n1227;
  assign n1229 = n1226 & ~n1228;
  assign n1230 = n924 & ~n1229;
  assign n1231 = Ni34 & n934;
  assign n1232 = n1226 & n1231;
  assign n1233 = n1230 & ~n1232;
  assign n1234 = Ni34 & n917;
  assign n1235 = ~n919 & ~n1234;
  assign n1236 = n903 & n1191;
  assign n1237 = n1235 & n1236;
  assign n1238 = ~Pi20 & ~n1237;
  assign n1239 = ~n1233 & n1238;
  assign n1240 = ~n1222 & n1239;
  assign n1241 = ~n1208 & n1240;
  assign n1242 = n1195 & n1197;
  assign n1243 = ~n899 & n1242;
  assign n1244 = ~Ni34 & ~n899;
  assign n1245 = Ni33 & ~n1244;
  assign n1246 = n1199 & n1245;
  assign n1247 = ~n1196 & ~n1246;
  assign n1248 = Ni34 & n899;
  assign n1249 = ~n901 & ~n1248;
  assign n1250 = n1191 & n1249;
  assign n1251 = n1247 & ~n1250;
  assign n1252 = ~n1243 & n1251;
  assign n1253 = n869 & ~n1252;
  assign n1254 = Ni33 & n917;
  assign n1255 = ~n1210 & ~n1254;
  assign n1256 = n1199 & ~n1255;
  assign n1257 = ~n917 & n1197;
  assign n1258 = ~n1196 & ~n1257;
  assign n1259 = ~n1256 & n1258;
  assign n1260 = n903 & ~n1259;
  assign n1261 = ~n1003 & n1191;
  assign n1262 = ~Ni34 & ~n1001;
  assign n1263 = Ni33 & ~n1262;
  assign n1264 = n1199 & n1263;
  assign n1265 = n1198 & ~n1264;
  assign n1266 = ~n1261 & n1265;
  assign n1267 = n994 & ~n1266;
  assign n1268 = n1001 & n1219;
  assign n1269 = ~n1264 & n1268;
  assign n1270 = n1267 & ~n1269;
  assign n1271 = ~n1260 & ~n1270;
  assign n1272 = ~n1253 & n1271;
  assign n1273 = n1241 & n1272;
  assign n1274 = Ni34 & n1086_1;
  assign n1275 = ~n1088 & n1191;
  assign n1276 = ~n1274 & n1275;
  assign n1277 = Ni33 & n1086_1;
  assign n1278 = ~n1210 & ~n1277;
  assign n1279 = n1199 & ~n1278;
  assign n1280 = ~n1086_1 & n1197;
  assign n1281 = ~n1196 & ~n1280;
  assign n1282 = ~n1279 & n1281;
  assign n1283 = ~n1276 & n1282;
  assign n1284 = n869 & ~n1283;
  assign n1285 = ~Ni34 & ~n1100;
  assign n1286 = Ni33 & ~n1285;
  assign n1287 = n1199 & n1286;
  assign n1288 = ~n1196 & ~n1287;
  assign n1289 = Ni34 & n1100;
  assign n1290 = ~n1102 & n1191;
  assign n1291 = ~n1100 & n1242;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = ~n1289 & ~n1292;
  assign n1294 = n1288 & ~n1293;
  assign n1295 = n903 & ~n1294;
  assign n1296 = ~Ni34 & ~n946;
  assign n1297 = Ni33 & ~n1296;
  assign n1298 = n1199 & n1297;
  assign n1299 = ~n1196 & ~n1298;
  assign n1300 = ~n948 & ~n1227;
  assign n1301 = n1299 & ~n1300;
  assign n1302 = n924 & ~n1301;
  assign n1303 = Ni34 & n946;
  assign n1304 = n1299 & n1303;
  assign n1305 = n1302 & ~n1304;
  assign n1306 = Ni33 & n1010;
  assign n1307 = ~n1210 & ~n1306;
  assign n1308 = n1199 & ~n1307;
  assign n1309 = ~n1196 & ~n1308;
  assign n1310 = ~n1012_1 & ~n1227;
  assign n1311 = n1309 & ~n1310;
  assign n1312 = n994 & ~n1311;
  assign n1313 = Ni34 & n1010;
  assign n1314 = n1309 & n1313;
  assign n1315 = n1312 & ~n1314;
  assign n1316 = n955 & n988;
  assign n1317 = n1218 & n1316;
  assign n1318 = Pi20 & ~n1317;
  assign n1319 = ~n1315 & n1318;
  assign n1320 = ~n1305 & n1319;
  assign n1321 = ~n1069 & ~n1227;
  assign n1322 = ~Ni34 & ~n1067;
  assign n1323 = Ni33 & ~n1322;
  assign n1324 = n1199 & n1323;
  assign n1325 = ~n1196 & ~n1324;
  assign n1326 = ~n1321 & n1325;
  assign n1327 = n1035 & ~n1326;
  assign n1328 = Ni34 & n1067;
  assign n1329 = n1325 & n1328;
  assign n1330 = n1327 & ~n1329;
  assign n1331 = ~n990 & n1191;
  assign n1332 = Ni33 & n988;
  assign n1333 = ~n1210 & ~n1332;
  assign n1334 = n1199 & ~n1333;
  assign n1335 = n1198 & ~n1334;
  assign n1336 = ~n1331 & n1335;
  assign n1337 = n955 & ~n1336;
  assign n1338 = n988 & ~n1334;
  assign n1339 = ~n1196 & n1338;
  assign n1340 = n1337 & ~n1339;
  assign n1341 = ~n1330 & ~n1340;
  assign n1342 = n1320 & n1341;
  assign n1343 = ~n1295 & n1342;
  assign n1344 = ~n1284 & n1343;
  assign n1345 = ~n1273 & ~n1344;
  assign n1346 = ~n18 & n1026;
  assign n1347 = ~n18 & n1217;
  assign n1348 = ~n18 & ~n1025;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1346 & n1349;
  assign n1351 = ~n1029 & ~n1350;
  assign n1352 = n864 & n1351;
  assign n1353 = n1026 & ~n1210;
  assign n1354 = Ni33 & n1025;
  assign n1355 = ~n1210 & ~n1354;
  assign n1356 = n1199 & ~n1355;
  assign n1357 = ~n1353 & n1356;
  assign n1358 = ~n1027_1 & n1197;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1352 & n1359;
  assign n1361 = ~n1196 & n1360;
  assign n1362 = n744 & ~n1361;
  assign n1363 = Ni33 & n1017;
  assign n1364 = ~n1210 & ~n1363;
  assign n1365 = n1199 & ~n1364;
  assign n1366 = ~n1196 & ~n1365;
  assign n1367 = n1018 & ~n1210;
  assign n1368 = n1365 & ~n1367;
  assign n1369 = n1198 & ~n1368;
  assign n1370 = ~n1366 & ~n1369;
  assign n1371 = ~n1021 & n1191;
  assign n1372 = n1217 & n1371;
  assign n1373 = ~n1370 & ~n1372;
  assign n1374 = n1369 & ~n1371;
  assign n1375 = ~n1019 & ~n1374;
  assign n1376 = n1373 & ~n1375;
  assign n1377 = n731 & ~n1376;
  assign n1378 = ~n1362 & ~n1377;
  assign n1379 = ~n1345 & n1378;
  assign n1380 = n1190 & ~n1379;
  assign n1381 = Pi15 & n570;
  assign n1382 = ~n1017 & n1197;
  assign n1383 = ~n1180 & n1191;
  assign n1384 = n1017 & ~n1347;
  assign n1385 = n1383 & ~n1384;
  assign n1386 = n1366 & ~n1385;
  assign n1387 = ~n1382 & n1386;
  assign n1388 = n731 & ~n1387;
  assign n1389 = Ni33 & n1137;
  assign n1390 = ~n1210 & ~n1389;
  assign n1391 = n1199 & ~n1390;
  assign n1392 = ~n1196 & ~n1391;
  assign n1393 = n869 & ~n1392;
  assign n1394 = n1140 & ~n1227;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = n1137 & n1392;
  assign n1397 = Ni34 & n1396;
  assign n1398 = ~n1395 & ~n1397;
  assign n1399 = ~n1148 & ~n1227;
  assign n1400 = n1146 & n1399;
  assign n1401 = ~n1145 & n1296;
  assign n1402 = Ni33 & ~n1401;
  assign n1403 = n1199 & n1402;
  assign n1404 = ~n1196 & ~n1403;
  assign n1405 = ~n1146 & n1218;
  assign n1406 = n1404 & ~n1405;
  assign n1407 = ~n1400 & n1406;
  assign n1408 = n924 & ~n1407;
  assign n1409 = ~n1398 & ~n1408;
  assign n1410 = Ni33 & n1141;
  assign n1411 = ~n1210 & ~n1410;
  assign n1412 = n1199 & ~n1411;
  assign n1413 = n1198 & ~n1412;
  assign n1414 = n903 & ~n1413;
  assign n1415 = n1144 & n1191;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = n1219 & ~n1412;
  assign n1418 = n1141 & n1417;
  assign n1419 = ~n1416 & ~n1418;
  assign n1420 = Ni33 & n1168;
  assign n1421 = ~n1210 & ~n1420;
  assign n1422 = n1199 & ~n1421;
  assign n1423 = ~n1196 & ~n1422;
  assign n1424 = ~n1170 & ~n1227;
  assign n1425 = n1423 & ~n1424;
  assign n1426 = n1035 & ~n1425;
  assign n1427 = Ni34 & n1168;
  assign n1428 = n1423 & n1427;
  assign n1429 = n1426 & ~n1428;
  assign n1430 = Ni33 & ~n1115;
  assign n1431 = ~n1210 & ~n1430;
  assign n1432 = n1199 & ~n1431;
  assign n1433 = ~n1196 & ~n1432;
  assign n1434 = ~n1117 & ~n1227;
  assign n1435 = n1433 & ~n1434;
  assign n1436 = n994 & ~n1435;
  assign n1437 = Ni34 & ~n1115;
  assign n1438 = n1433 & n1437;
  assign n1439 = n1436 & ~n1438;
  assign n1440 = ~n1429 & ~n1439;
  assign n1441 = ~n1419 & n1440;
  assign n1442 = ~n1160 & n1191;
  assign n1443 = Ni33 & n1158;
  assign n1444 = ~n1210 & ~n1443;
  assign n1445 = n1199 & ~n1444;
  assign n1446 = n1198 & ~n1445;
  assign n1447 = ~n1442 & n1446;
  assign n1448 = n955 & ~n1447;
  assign n1449 = n1219 & ~n1445;
  assign n1450 = n1158 & n1449;
  assign n1451 = n1448 & ~n1450;
  assign n1452 = Pi20 & ~n1451;
  assign n1453 = n1441 & n1452;
  assign n1454 = n1409 & n1453;
  assign n1455 = Ni33 & ~n1110;
  assign n1456 = ~n1210 & ~n1455;
  assign n1457 = n1199 & ~n1456;
  assign n1458 = ~n1196 & ~n1457;
  assign n1459 = ~n1112 & ~n1227;
  assign n1460 = n1458 & ~n1459;
  assign n1461 = n994 & ~n1460;
  assign n1462 = Ni34 & ~n1110;
  assign n1463 = n1458 & n1462;
  assign n1464 = n1461 & ~n1463;
  assign n1465 = ~Ni34 & ~n1125;
  assign n1466 = Ni33 & ~n1465;
  assign n1467 = n1199 & n1466;
  assign n1468 = n1198 & ~n1467;
  assign n1469 = n869 & ~n1468;
  assign n1470 = n1125 & ~n1467;
  assign n1471 = ~n1196 & n1470;
  assign n1472 = n1469 & ~n1471;
  assign n1473 = Ni33 & n1121;
  assign n1474 = ~n1210 & ~n1473;
  assign n1475 = n1199 & ~n1474;
  assign n1476 = n1198 & ~n1475;
  assign n1477 = n903 & ~n1476;
  assign n1478 = n1121 & ~n1475;
  assign n1479 = ~n1196 & n1478;
  assign n1480 = n1477 & ~n1479;
  assign n1481 = ~n1472 & ~n1480;
  assign n1482 = ~n1133 & n1191;
  assign n1483 = Ni34 & n1131;
  assign n1484 = n1482 & ~n1483;
  assign n1485 = Ni33 & n1131;
  assign n1486 = ~n1210 & ~n1485;
  assign n1487 = n1199 & ~n1486;
  assign n1488 = ~n1131 & n1197;
  assign n1489 = ~n1196 & ~n1488;
  assign n1490 = ~n1487 & n1489;
  assign n1491 = ~n1484 & n1490;
  assign n1492 = n924 & ~n1491;
  assign n1493 = Ni34 & n1121;
  assign n1494 = ~n1123 & ~n1493;
  assign n1495 = n1236 & n1494;
  assign n1496 = n1125 & ~n1217;
  assign n1497 = ~n1465 & ~n1496;
  assign n1498 = n869 & n1191;
  assign n1499 = n1497 & n1498;
  assign n1500 = ~n1495 & ~n1499;
  assign n1501 = ~Pi20 & n1500;
  assign n1502 = ~n1492 & n1501;
  assign n1503 = ~n1156 & ~n1227;
  assign n1504 = Ni33 & n1154;
  assign n1505 = ~n1210 & ~n1504;
  assign n1506 = n1199 & ~n1505;
  assign n1507 = ~n1196 & ~n1506;
  assign n1508 = ~n1503 & n1507;
  assign n1509 = n955 & ~n1508;
  assign n1510 = Ni34 & n1154;
  assign n1511 = n1507 & n1510;
  assign n1512 = n1509 & ~n1511;
  assign n1513 = ~Ni34 & ~n1164;
  assign n1514 = Ni33 & ~n1513;
  assign n1515 = n1199 & n1514;
  assign n1516 = ~n1196 & ~n1515;
  assign n1517 = ~n1166 & ~n1227;
  assign n1518 = n1516 & ~n1517;
  assign n1519 = n1035 & ~n1518;
  assign n1520 = Ni34 & n1164;
  assign n1521 = n1516 & n1520;
  assign n1522 = n1519 & ~n1521;
  assign n1523 = ~n1512 & ~n1522;
  assign n1524 = n1502 & n1523;
  assign n1525 = n1481 & n1524;
  assign n1526 = ~n1464 & n1525;
  assign n1527 = ~n1454 & ~n1526;
  assign n1528 = n744 & n864;
  assign n1529 = ~n1175 & ~n1349;
  assign n1530 = n1528 & n1529;
  assign n1531 = ~n1196 & ~n1356;
  assign n1532 = ~n1197 & n1531;
  assign n1533 = n744 & ~n1532;
  assign n1534 = n1025 & n1531;
  assign n1535 = n1533 & ~n1534;
  assign n1536 = ~n1530 & ~n1535;
  assign n1537 = ~n1527 & n1536;
  assign n1538 = ~n1388 & n1537;
  assign n1539 = n1381 & ~n1538;
  assign n1540 = ~n1192 & n1203;
  assign n1541 = n1035 & ~n1540;
  assign n1542 = n869 & ~n1247;
  assign n1543 = n902 & ~n1227;
  assign n1544 = ~n1230 & ~n1543;
  assign n1545 = ~n1542 & n1544;
  assign n1546 = ~n1541 & n1545;
  assign n1547 = ~n919 & n1191;
  assign n1548 = n1198 & ~n1256;
  assign n1549 = ~n1547 & n1548;
  assign n1550 = n903 & ~n1549;
  assign n1551 = ~Pi20 & ~n1267;
  assign n1552 = ~n1216 & n1551;
  assign n1553 = ~n1550 & n1552;
  assign n1554 = n1546 & n1553;
  assign n1555 = n1198 & ~n1290;
  assign n1556 = ~n1287 & n1555;
  assign n1557 = n903 & ~n1556;
  assign n1558 = Pi20 & ~n1302;
  assign n1559 = ~n1327 & n1558;
  assign n1560 = n1198 & ~n1279;
  assign n1561 = ~n1275 & n1560;
  assign n1562 = n869 & ~n1561;
  assign n1563 = ~n1312 & ~n1337;
  assign n1564 = ~n1562 & n1563;
  assign n1565 = n1559 & n1564;
  assign n1566 = ~n1557 & n1565;
  assign n1567 = ~n1554 & ~n1566;
  assign n1568 = n731 & ~n1374;
  assign n1569 = ~n1029 & n1191;
  assign n1570 = n1198 & ~n1357;
  assign n1571 = ~n1569 & n1570;
  assign n1572 = n744 & ~n1571;
  assign n1573 = ~Pi15 & ~n1572;
  assign n1574 = ~n1568 & n1573;
  assign n1575 = ~n1567 & n1574;
  assign n1576 = n1198 & ~n1365;
  assign n1577 = ~n1383 & n1576;
  assign n1578 = n731 & ~n1577;
  assign n1579 = Pi20 & n1416;
  assign n1580 = ~n1436 & n1579;
  assign n1581 = ~n1426 & ~n1448;
  assign n1582 = ~n1399 & n1404;
  assign n1583 = n924 & ~n1582;
  assign n1584 = n1395 & ~n1583;
  assign n1585 = n1581 & n1584;
  assign n1586 = n1580 & n1585;
  assign n1587 = ~n1477 & ~n1519;
  assign n1588 = n1198 & ~n1487;
  assign n1589 = ~n1482 & n1588;
  assign n1590 = n924 & ~n1589;
  assign n1591 = ~Pi20 & ~n1590;
  assign n1592 = n1587 & n1591;
  assign n1593 = ~n1469 & ~n1509;
  assign n1594 = ~n1129 & n1191;
  assign n1595 = n1593 & ~n1594;
  assign n1596 = n1592 & n1595;
  assign n1597 = ~n1461 & n1596;
  assign n1598 = ~n1586 & ~n1597;
  assign n1599 = ~n18 & n1528;
  assign n1600 = ~n1175 & n1599;
  assign n1601 = ~n1533 & ~n1600;
  assign n1602 = Pi15 & n1601;
  assign n1603 = ~n1598 & n1602;
  assign n1604 = ~n1578 & n1603;
  assign n1605 = ~n1575 & ~n1604;
  assign n1606 = ~n570 & n1605;
  assign n1607 = ~n1539 & ~n1606;
  assign n1608 = ~n1380 & n1607;
  assign n1609 = Ni10 & ~n1608;
  assign n1610 = ~Pi16 & ~Pi15;
  assign n1611 = Pi19 & n949;
  assign n1612 = Pi25 & n1217;
  assign n1613 = P__cmxig_0 & n1612;
  assign n1614 = n1100 & n1613;
  assign n1615 = Pi25 & ~n18;
  assign n1616 = ~n1289 & n1615;
  assign n1617 = ~n1102 & n1616;
  assign n1618 = n18 & n871;
  assign n1619 = Pi25 & n1618;
  assign n1620 = n1286 & n1619;
  assign n1621 = ~n1617 & ~n1620;
  assign n1622 = ~n1614 & n1621;
  assign n1623 = n1611 & ~n1622;
  assign n1624 = ~Pi19 & n864;
  assign n1625 = ~Pi20 & n1624;
  assign n1626 = n1263 & n1619;
  assign n1627 = n1001 & ~n1217;
  assign n1628 = n1615 & ~n1627;
  assign n1629 = ~n1262 & n1628;
  assign n1630 = n1001 & n1613;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n1626 & n1631;
  assign n1633 = n1625 & ~n1632;
  assign n1634 = ~n1623 & ~n1633;
  assign n1635 = ~n1002_1 & n1625;
  assign n1636 = Pi19 & n867;
  assign n1637 = ~n918 & n1636;
  assign n1638 = ~n1101 & n1611;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n1635 & n1639;
  assign n1641 = Ni34 & ~n1640;
  assign n1642 = Ni34 & ~n864;
  assign n1643 = Pi20 & n1624;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = n1210 & n1618;
  assign n1646 = ~n1642 & ~n1645;
  assign n1647 = Ni34 & ~n1011;
  assign n1648 = n1646 & ~n1647;
  assign n1649 = ~n1644 & ~n1648;
  assign n1650 = Pi20 & ~Pi19;
  assign n1651 = n1210 & ~n1650;
  assign n1652 = n1199 & n1651;
  assign n1653 = ~n1649 & ~n1652;
  assign n1654 = ~n1641 & n1653;
  assign n1655 = ~n1255 & n1619;
  assign n1656 = n1235 & n1615;
  assign n1657 = n917 & n1613;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1655 & n1658;
  assign n1660 = n1636 & ~n1659;
  assign n1661 = n1010 & n1613;
  assign n1662 = ~n1307 & n1619;
  assign n1663 = ~n1313 & n1615;
  assign n1664 = ~n1012_1 & n1663;
  assign n1665 = ~n1662 & ~n1664;
  assign n1666 = ~n1661 & n1665;
  assign n1667 = n1643 & ~n1666;
  assign n1668 = ~n1660 & ~n1667;
  assign n1669 = n1654 & n1668;
  assign n1670 = n1634 & n1669;
  assign n1671 = n1610 & ~n1670;
  assign n1672 = Pi16 & ~Pi15;
  assign n1673 = Ni34 & n969;
  assign n1674 = ~n971 & n1615;
  assign n1675 = ~n1673 & n1674;
  assign n1676 = n969 & n1613;
  assign n1677 = ~n1212 & n1619;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1675 & n1678;
  assign n1680 = n1636 & ~n1679;
  assign n1681 = n934 & n1613;
  assign n1682 = n1224 & n1619;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1231 & n1615;
  assign n1685 = ~n936 & n1684;
  assign n1686 = n1683 & ~n1685;
  assign n1687 = n1625 & ~n1686;
  assign n1688 = ~n1611 & ~n1642;
  assign n1689 = Ni34 & ~n989;
  assign n1690 = n1646 & ~n1689;
  assign n1691 = ~n1688 & ~n1690;
  assign n1692 = Ni34 & ~n935;
  assign n1693 = ~n1645 & ~n1692;
  assign n1694 = n1625 & ~n1693;
  assign n1695 = Ni34 & ~n947;
  assign n1696 = ~n1645 & ~n1695;
  assign n1697 = n1643 & ~n1696;
  assign n1698 = ~n1694 & ~n1697;
  assign n1699 = ~n1691 & n1698;
  assign n1700 = n1297 & n1619;
  assign n1701 = n946 & n1613;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1303 & n1615;
  assign n1704 = ~n948 & n1703;
  assign n1705 = n1702 & ~n1704;
  assign n1706 = n1643 & ~n1705;
  assign n1707 = n1699 & ~n1706;
  assign n1708 = ~n1687 & n1707;
  assign n1709 = Ni34 & ~n970;
  assign n1710 = ~n1645 & ~n1709;
  assign n1711 = n1636 & ~n1710;
  assign n1712 = ~P__cmxig_1 & n1612;
  assign n1713 = n988 & n1712;
  assign n1714 = ~n1333 & n1619;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = n1611 & ~n1715;
  assign n1717 = ~n1711 & ~n1716;
  assign n1718 = n1708 & n1717;
  assign n1719 = ~n1680 & n1718;
  assign n1720 = n1672 & ~n1719;
  assign n1721 = ~n1110 & n1613;
  assign n1722 = Ni34 & ~n1111;
  assign n1723 = ~n1645 & ~n1722;
  assign n1724 = ~n1456 & n1619;
  assign n1725 = ~n1462 & n1615;
  assign n1726 = ~n1112 & n1725;
  assign n1727 = ~n1724 & ~n1726;
  assign n1728 = n1723 & n1727;
  assign n1729 = ~n1721 & n1728;
  assign n1730 = n1625 & ~n1729;
  assign n1731 = Ni34 & ~n1116;
  assign n1732 = n1646 & ~n1731;
  assign n1733 = ~n1644 & ~n1732;
  assign n1734 = Ni34 & ~n1142;
  assign n1735 = ~n1645 & ~n1734;
  assign n1736 = n1611 & ~n1735;
  assign n1737 = Ni34 & ~n1122;
  assign n1738 = ~n1645 & ~n1737;
  assign n1739 = n1636 & ~n1738;
  assign n1740 = ~n1736 & ~n1739;
  assign n1741 = ~n1733 & n1740;
  assign n1742 = n1141 & n1613;
  assign n1743 = Ni34 & n1141;
  assign n1744 = n1615 & ~n1743;
  assign n1745 = ~n1143 & n1744;
  assign n1746 = ~n1411 & n1619;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n1742 & n1747;
  assign n1749 = n1611 & ~n1748;
  assign n1750 = n1741 & ~n1749;
  assign n1751 = ~n1115 & n1613;
  assign n1752 = ~n1431 & n1619;
  assign n1753 = ~n1437 & n1615;
  assign n1754 = ~n1117 & n1753;
  assign n1755 = ~n1752 & ~n1754;
  assign n1756 = ~n1751 & n1755;
  assign n1757 = n1643 & ~n1756;
  assign n1758 = n1494 & n1615;
  assign n1759 = ~n1474 & n1619;
  assign n1760 = n1121 & n1613;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n1758 & n1761;
  assign n1763 = n1636 & ~n1762;
  assign n1764 = ~n1757 & ~n1763;
  assign n1765 = n1750 & n1764;
  assign n1766 = ~n1730 & n1765;
  assign n1767 = n1178 & ~n1766;
  assign n1768 = ~n1720 & ~n1767;
  assign n1769 = Pi16 & Pi15;
  assign n1770 = ~n1483 & n1615;
  assign n1771 = ~n1133 & n1770;
  assign n1772 = n1131 & n1613;
  assign n1773 = ~n1486 & n1619;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1771 & n1774;
  assign n1776 = n1625 & ~n1775;
  assign n1777 = ~n1444 & n1619;
  assign n1778 = n1158 & n1712;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = n1611 & ~n1779;
  assign n1781 = ~n1776 & ~n1780;
  assign n1782 = Ni34 & ~n1132;
  assign n1783 = ~n1645 & ~n1782;
  assign n1784 = n1625 & ~n1783;
  assign n1785 = Ni34 & ~n1159;
  assign n1786 = n1646 & ~n1785;
  assign n1787 = ~n1688 & ~n1786;
  assign n1788 = ~n1784 & ~n1787;
  assign n1789 = ~n1146 & n1712;
  assign n1790 = Ni34 & ~n1147;
  assign n1791 = ~n1645 & ~n1790;
  assign n1792 = n1402 & n1619;
  assign n1793 = n1791 & ~n1792;
  assign n1794 = ~n1789 & n1793;
  assign n1795 = n1643 & ~n1794;
  assign n1796 = ~n1505 & n1619;
  assign n1797 = Ni34 & ~n1155;
  assign n1798 = ~n1645 & ~n1797;
  assign n1799 = ~n1510 & n1615;
  assign n1800 = ~n1156 & n1799;
  assign n1801 = n1154 & n1613;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n1798 & n1802;
  assign n1804 = ~n1796 & n1803;
  assign n1805 = n1636 & ~n1804;
  assign n1806 = ~n1795 & ~n1805;
  assign n1807 = n1788 & n1806;
  assign n1808 = n1781 & n1807;
  assign n1809 = n1769 & ~n1808;
  assign n1810 = ~Pi17 & ~n1809;
  assign n1811 = n1768 & n1810;
  assign n1812 = ~n1671 & n1811;
  assign n1813 = ~Ni10 & n570;
  assign n1814 = Pi19 & n864;
  assign n1815 = ~n1642 & ~n1814;
  assign n1816 = ~n1364 & n1619;
  assign n1817 = n1017 & n1712;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1815 & ~n1818;
  assign n1820 = Ni34 & ~n1126;
  assign n1821 = ~n1645 & ~n1820;
  assign n1822 = n1625 & ~n1821;
  assign n1823 = Ni34 & ~n1179;
  assign n1824 = n1646 & ~n1823;
  assign n1825 = ~n1815 & ~n1824;
  assign n1826 = Ni34 & ~n1138;
  assign n1827 = ~n1645 & ~n1826;
  assign n1828 = n1643 & ~n1827;
  assign n1829 = ~n1825 & ~n1828;
  assign n1830 = ~n1822 & n1829;
  assign n1831 = ~n1390 & n1619;
  assign n1832 = n1137 & n1712;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = n1643 & ~n1833;
  assign n1835 = n1125 & n1613;
  assign n1836 = n1497 & n1615;
  assign n1837 = n1466 & n1619;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = ~n1835 & n1838;
  assign n1840 = n1625 & ~n1839;
  assign n1841 = ~n1834 & ~n1840;
  assign n1842 = n1830 & n1841;
  assign n1843 = ~n1819 & n1842;
  assign n1844 = n1178 & ~n1843;
  assign n1845 = n1514 & n1619;
  assign n1846 = Ni34 & ~n1165;
  assign n1847 = ~n1645 & ~n1846;
  assign n1848 = n1164 & n1613;
  assign n1849 = ~n1520 & n1615;
  assign n1850 = ~n1166 & n1849;
  assign n1851 = ~n1848 & ~n1850;
  assign n1852 = n1847 & n1851;
  assign n1853 = ~n1845 & n1852;
  assign n1854 = n1625 & ~n1853;
  assign n1855 = ~n1427 & n1615;
  assign n1856 = ~n1170 & n1855;
  assign n1857 = n1168 & n1613;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = Ni34 & ~n1169;
  assign n1860 = ~n1645 & ~n1859;
  assign n1861 = ~n1421 & n1619;
  assign n1862 = n1860 & ~n1861;
  assign n1863 = n1858 & n1862;
  assign n1864 = n1643 & ~n1863;
  assign n1865 = Pi25 & n1529;
  assign n1866 = ~n1355 & n1619;
  assign n1867 = Ni34 & ~n1174;
  assign n1868 = n1646 & ~n1867;
  assign n1869 = n1025 & n1613;
  assign n1870 = n1868 & ~n1869;
  assign n1871 = ~n1866 & n1870;
  assign n1872 = ~n1865 & n1871;
  assign n1873 = ~n1815 & ~n1872;
  assign n1874 = ~n1864 & ~n1873;
  assign n1875 = ~n1854 & n1874;
  assign n1876 = n1769 & ~n1875;
  assign n1877 = ~n1844 & ~n1876;
  assign n1878 = n1672 & n1814;
  assign n1879 = ~n1026 & n1869;
  assign n1880 = Pi25 & n1351;
  assign n1881 = ~n1353 & n1866;
  assign n1882 = ~n1880 & ~n1881;
  assign n1883 = ~n1879 & n1882;
  assign n1884 = n1878 & ~n1883;
  assign n1885 = n1245 & n1619;
  assign n1886 = n1249 & n1615;
  assign n1887 = Ni34 & ~n900;
  assign n1888 = ~n1645 & ~n1887;
  assign n1889 = n899 & n1613;
  assign n1890 = n1888 & ~n1889;
  assign n1891 = ~n1886 & n1890;
  assign n1892 = ~n1885 & n1891;
  assign n1893 = n1625 & ~n1892;
  assign n1894 = n1086_1 & n1613;
  assign n1895 = ~n1274 & n1615;
  assign n1896 = ~n1088 & n1895;
  assign n1897 = ~n1894 & ~n1896;
  assign n1898 = Ni34 & ~n1087;
  assign n1899 = ~n1645 & ~n1898;
  assign n1900 = ~n1278 & n1619;
  assign n1901 = n1899 & ~n1900;
  assign n1902 = n1897 & n1901;
  assign n1903 = n1643 & ~n1902;
  assign n1904 = ~n1367 & n1816;
  assign n1905 = n1020 & n1347;
  assign n1906 = Pi25 & n1905;
  assign n1907 = ~n1904 & ~n1906;
  assign n1908 = Ni34 & ~n1020;
  assign n1909 = n1019 & n1613;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1646 & n1910;
  assign n1912 = n1907 & n1911;
  assign n1913 = ~n1815 & ~n1912;
  assign n1914 = ~n1903 & ~n1913;
  assign n1915 = ~n1893 & n1914;
  assign n1916 = n1610 & ~n1915;
  assign n1917 = ~n1884 & ~n1916;
  assign n1918 = Ni34 & ~n1027_1;
  assign n1919 = ~n1196 & ~n1645;
  assign n1920 = ~n1918 & n1919;
  assign n1921 = ~n1815 & ~n1920;
  assign n1922 = n1049 & n1712;
  assign n1923 = Ni34 & ~n1050;
  assign n1924 = ~n1645 & ~n1923;
  assign n1925 = n1201 & n1619;
  assign n1926 = n1924 & ~n1925;
  assign n1927 = ~n1922 & n1926;
  assign n1928 = n1625 & ~n1927;
  assign n1929 = n1067 & n1613;
  assign n1930 = Ni34 & ~n1068;
  assign n1931 = ~n1645 & ~n1930;
  assign n1932 = ~n1328 & n1615;
  assign n1933 = ~n1069 & n1932;
  assign n1934 = n1323 & n1619;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = n1931 & n1935;
  assign n1937 = ~n1929 & n1936;
  assign n1938 = n1643 & ~n1937;
  assign n1939 = ~n1928 & ~n1938;
  assign n1940 = ~n1921 & n1939;
  assign n1941 = n1672 & ~n1940;
  assign n1942 = Pi17 & ~n1941;
  assign n1943 = n1917 & n1942;
  assign n1944 = n1877 & n1943;
  assign n1945 = n1813 & ~n1944;
  assign n1946 = ~n1812 & n1945;
  assign n1947 = ~n1609 & ~n1946;
  assign n1948 = ~n1189 & n1947;
  assign n1949 = n580 & ~n1948;
  assign n1950 = n1625 & ~n1723;
  assign n1951 = n1741 & ~n1950;
  assign n1952 = n1178 & ~n1951;
  assign n1953 = n1699 & ~n1711;
  assign n1954 = n1672 & ~n1953;
  assign n1955 = ~n1952 & ~n1954;
  assign n1956 = n1610 & ~n1654;
  assign n1957 = n1636 & ~n1798;
  assign n1958 = n1643 & ~n1791;
  assign n1959 = n1788 & ~n1958;
  assign n1960 = ~n1957 & n1959;
  assign n1961 = n1769 & ~n1960;
  assign n1962 = ~Pi17 & ~n1961;
  assign n1963 = ~n1956 & n1962;
  assign n1964 = n1955 & n1963;
  assign n1965 = n864 & ~n1645;
  assign n1966 = ~n1908 & n1965;
  assign n1967 = ~n1624 & ~n1966;
  assign n1968 = ~Pi20 & ~Pi19;
  assign n1969 = ~n1888 & n1968;
  assign n1970 = n1650 & ~n1899;
  assign n1971 = ~n1969 & ~n1970;
  assign n1972 = ~n1967 & n1971;
  assign n1973 = n1610 & ~n1972;
  assign n1974 = n1178 & ~n1830;
  assign n1975 = n1643 & ~n1860;
  assign n1976 = ~n1815 & ~n1868;
  assign n1977 = n1625 & ~n1847;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1975 & n1978;
  assign n1980 = n1769 & ~n1979;
  assign n1981 = n1643 & ~n1931;
  assign n1982 = n1625 & ~n1924;
  assign n1983 = ~n1921 & ~n1982;
  assign n1984 = ~n1981 & n1983;
  assign n1985 = n1672 & ~n1984;
  assign n1986 = ~n1980 & ~n1985;
  assign n1987 = ~n1974 & n1986;
  assign n1988 = Pi17 & n1987;
  assign n1989 = ~n1973 & n1988;
  assign n1990 = ~n1964 & ~n1989;
  assign n1991 = n571 & ~n1990;
  assign n1992 = Ni34 & ~n1991;
  assign n1993 = ~n580 & n1992;
  assign n1002 = n1949 | n1993;
  assign n1995 = Ni33 & ~n871;
  assign n1996 = Ni46 & Ni45;
  assign n1997 = n871 & n1996;
  assign n1998 = ~n1995 & ~n1997;
  assign n1999 = ~Pi21 & ~n1998;
  assign n2000 = ~Pi22 & Pi21;
  assign n2001 = Ni48 & Ni47;
  assign n2002 = ~Ni45 & n2001;
  assign n2003 = ~n1996 & ~n2002;
  assign n2004 = n871 & ~n2003;
  assign n2005 = ~n1995 & ~n2004;
  assign n2006 = n2000 & ~n2005;
  assign n2007 = ~n1999 & ~n2006;
  assign n2008 = ~n864 & n1995;
  assign n2009 = ~n872 & n2003;
  assign n2010 = ~Pi22 & ~n2009;
  assign n2011 = ~Ni46 & Ni45;
  assign n2012 = ~Pi21 & ~n2011;
  assign n2013 = ~n2010 & ~n2012;
  assign n2014 = n871 & ~n2013;
  assign n2015 = ~n2008 & ~n2014;
  assign n2016 = Pi20 & ~n2015;
  assign n2017 = n2007 & ~n2016;
  assign n2018 = ~Ni33 & n870;
  assign n2019 = ~Ni32 & n2018;
  assign n2020 = Ni39 & n872;
  assign n2021 = n2003 & ~n2020;
  assign n2022 = n873 & ~n2021;
  assign n2023 = ~n881 & n2003;
  assign n2024 = ~Ni42 & n2003;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n873 & n2025;
  assign n2027 = ~n2022 & ~n2026;
  assign n2028 = n2019 & ~n2027;
  assign n2029 = ~Ni44 & ~Ni43;
  assign n2030 = n872 & ~n2029;
  assign n2031 = n2003 & ~n2030;
  assign n2032 = ~Ni42 & n872;
  assign n2033 = n2031 & ~n2032;
  assign n2034 = ~n873 & ~n2033;
  assign n2035 = n871 & ~n2022;
  assign n2036 = ~n2034 & n2035;
  assign n2037 = Ni33 & ~n2036;
  assign n2038 = ~n2028 & ~n2037;
  assign n2039 = n864 & ~n2038;
  assign n2040 = n2017 & ~n2039;
  assign n2041 = ~n570 & ~n2040;
  assign n2042 = Ni34 & n2019;
  assign n2043 = n864 & n2042;
  assign n2044 = ~n1006 & ~n2025;
  assign n2045 = Ni41 & ~n2025;
  assign n2046 = ~n1023 & n2023;
  assign n2047 = ~Ni40 & ~n2046;
  assign n2048 = ~n2045 & n2047;
  assign n2049 = n2044 & ~n2048;
  assign n2050 = n816 & ~n2049;
  assign n2051 = n750 & ~n2033;
  assign n2052 = n704 & ~n2049;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = n908 & ~n2053;
  assign n2055 = ~n2022 & ~n2051;
  assign n2056 = ~n890 & ~n2022;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = Ni38 & ~n816;
  assign n2059 = ~n938 & ~n2058;
  assign n2060 = ~n2049 & ~n2059;
  assign n2061 = ~n2057 & ~n2060;
  assign n2062 = ~n2054 & n2061;
  assign n2063 = ~n2050 & n2062;
  assign n2064 = n903 & ~n2063;
  assign n2065 = Ni41 & ~n2046;
  assign n2066 = ~Ni41 & ~n2044;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = ~n2047 & n2067;
  assign n2069 = n816 & ~n2068;
  assign n2070 = n704 & ~n2068;
  assign n2071 = ~n2051 & ~n2070;
  assign n2072 = n908 & ~n2071;
  assign n2073 = ~n2059 & ~n2068;
  assign n2074 = ~n2057 & ~n2073;
  assign n2075 = ~n2072 & n2074;
  assign n2076 = ~n2069 & n2075;
  assign n2077 = n955 & ~n2076;
  assign n2078 = ~n2064 & ~n2077;
  assign n2079 = ~n2044 & ~n2059;
  assign n2080 = ~n2057 & ~n2079;
  assign n2081 = n816 & ~n2044;
  assign n2082 = n2080 & ~n2081;
  assign n2083 = n994 & ~n2082;
  assign n2084 = n816 & ~n2067;
  assign n2085 = ~n2059 & ~n2067;
  assign n2086 = ~n2057 & ~n2085;
  assign n2087 = ~n2084 & n2086;
  assign n2088 = n924 & ~n2087;
  assign n2089 = ~n2083 & ~n2088;
  assign n2090 = n2078 & n2089;
  assign n2091 = Pi20 & ~n2090;
  assign n2092 = n2023 & ~n2065;
  assign n2093 = ~n2047 & n2092;
  assign n2094 = n816 & ~n2093;
  assign n2095 = n704 & ~n2093;
  assign n2096 = ~n2051 & ~n2095;
  assign n2097 = n908 & ~n2096;
  assign n2098 = ~Ni38 & n938;
  assign n2099 = ~n2033 & n2098;
  assign n2100 = ~n2022 & ~n2099;
  assign n2101 = ~n891 & ~n2058;
  assign n2102 = ~n2093 & ~n2101;
  assign n2103 = n2100 & ~n2102;
  assign n2104 = ~n2097 & n2103;
  assign n2105 = ~n2094 & n2104;
  assign n2106 = n955 & ~n2105;
  assign n2107 = ~Ni42 & Ni41;
  assign n2108 = n2003 & n2107;
  assign n2109 = ~n2023 & ~n2108;
  assign n2110 = ~n2048 & ~n2109;
  assign n2111 = n816 & ~n2110;
  assign n2112 = n704 & ~n2110;
  assign n2113 = ~n2051 & ~n2112;
  assign n2114 = n908 & ~n2113;
  assign n2115 = ~n2101 & ~n2110;
  assign n2116 = n2100 & ~n2115;
  assign n2117 = ~n2114 & n2116;
  assign n2118 = ~n2111 & n2117;
  assign n2119 = n903 & ~n2118;
  assign n2120 = ~n2106 & ~n2119;
  assign n2121 = ~n2101 & n2109;
  assign n2122 = n2100 & ~n2121;
  assign n2123 = n816 & n2109;
  assign n2124 = n2122 & ~n2123;
  assign n2125 = n994 & ~n2124;
  assign n2126 = n816 & ~n2092;
  assign n2127 = ~n2092 & ~n2101;
  assign n2128 = n2100 & ~n2127;
  assign n2129 = ~n2126 & n2128;
  assign n2130 = n924 & ~n2129;
  assign n2131 = ~n2125 & ~n2130;
  assign n2132 = n2120 & n2131;
  assign n2133 = ~Pi20 & ~n2132;
  assign n2134 = Pi17 & ~Pi16;
  assign n2135 = Ni40 & ~n2046;
  assign n2136 = ~n2045 & n2135;
  assign n2137 = ~n2109 & ~n2136;
  assign n2138 = n816 & ~n2137;
  assign n2139 = n704 & ~n2137;
  assign n2140 = ~n2051 & ~n2139;
  assign n2141 = n822 & ~n2140;
  assign n2142 = ~n2101 & ~n2137;
  assign n2143 = n2100 & ~n2142;
  assign n2144 = ~n2141 & n2143;
  assign n2145 = ~n2138 & n2144;
  assign n2146 = n1968 & ~n2145;
  assign n2147 = n2044 & ~n2136;
  assign n2148 = n816 & ~n2147;
  assign n2149 = n704 & ~n2147;
  assign n2150 = ~n2051 & ~n2149;
  assign n2151 = n822 & ~n2150;
  assign n2152 = ~n2059 & ~n2147;
  assign n2153 = ~n2057 & ~n2152;
  assign n2154 = ~n2151 & n2153;
  assign n2155 = ~n2148 & n2154;
  assign n2156 = n1650 & ~n2155;
  assign n2157 = ~n2146 & ~n2156;
  assign n2158 = n2134 & ~n2157;
  assign n2159 = Pi17 & Pi16;
  assign n2160 = n2092 & ~n2135;
  assign n2161 = n816 & ~n2160;
  assign n2162 = n704 & ~n2160;
  assign n2163 = ~n2051 & ~n2162;
  assign n2164 = n822 & ~n2163;
  assign n2165 = ~n2101 & ~n2160;
  assign n2166 = n2100 & ~n2165;
  assign n2167 = ~n2164 & n2166;
  assign n2168 = ~n2161 & n2167;
  assign n2169 = n1968 & ~n2168;
  assign n2170 = n2067 & ~n2135;
  assign n2171 = n816 & ~n2170;
  assign n2172 = n704 & ~n2170;
  assign n2173 = ~n2051 & ~n2172;
  assign n2174 = n822 & ~n2173;
  assign n2175 = ~n2059 & ~n2170;
  assign n2176 = ~n2057 & ~n2175;
  assign n2177 = ~n2174 & n2176;
  assign n2178 = ~n2171 & n2177;
  assign n2179 = n1650 & ~n2178;
  assign n2180 = ~n2169 & ~n2179;
  assign n2181 = n2159 & ~n2180;
  assign n2182 = ~n2158 & ~n2181;
  assign n2183 = ~n2133 & n2182;
  assign n2184 = ~n2091 & n2183;
  assign n2185 = n2043 & ~n2184;
  assign n2186 = ~Pi20 & ~n2007;
  assign n2187 = ~Ni34 & n2028;
  assign n2188 = ~n2037 & ~n2187;
  assign n2189 = n864 & ~n2188;
  assign n2190 = ~n2016 & ~n2189;
  assign n2191 = ~n2186 & n2190;
  assign n2192 = Ni36 & ~n873;
  assign n2193 = ~n2046 & n2192;
  assign n2194 = Ni38 & ~n2046;
  assign n2195 = n2055 & ~n2194;
  assign n2196 = Ni36 & ~n2022;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = ~n2193 & ~n2197;
  assign n2199 = n2042 & ~n2198;
  assign n2200 = n2188 & ~n2199;
  assign n2201 = n1528 & ~n2200;
  assign n2202 = ~n2055 & n2197;
  assign n2203 = n2045 & ~n2202;
  assign n2204 = n2199 & ~n2203;
  assign n2205 = n731 & n864;
  assign n2206 = n2204 & n2205;
  assign n2207 = ~n2201 & ~n2206;
  assign n2208 = n2191 & n2207;
  assign n2209 = ~n2185 & n2208;
  assign n2210 = n1190 & ~n2209;
  assign n2211 = n2042 & ~n2195;
  assign n2212 = n2045 & n2055;
  assign n2213 = ~Pi16 & n2212;
  assign n2214 = n2211 & ~n2213;
  assign n2215 = n2188 & ~n2214;
  assign n2216 = n1030 & ~n2215;
  assign n2217 = ~n822 & ~n2053;
  assign n2218 = n2061 & ~n2217;
  assign n2219 = n903 & ~n2218;
  assign n2220 = ~n822 & ~n2071;
  assign n2221 = n2074 & ~n2220;
  assign n2222 = n955 & ~n2221;
  assign n2223 = ~n2219 & ~n2222;
  assign n2224 = Ni36 & n2051;
  assign n2225 = Ni38 & n2084;
  assign n2226 = n2086 & ~n2225;
  assign n2227 = ~n2224 & n2226;
  assign n2228 = n924 & ~n2227;
  assign n2229 = Ni38 & n2081;
  assign n2230 = n2080 & ~n2224;
  assign n2231 = ~n2229 & n2230;
  assign n2232 = n994 & ~n2231;
  assign n2233 = ~n2228 & ~n2232;
  assign n2234 = n2223 & n2233;
  assign n2235 = Pi20 & ~n2234;
  assign n2236 = ~n822 & ~n2113;
  assign n2237 = n2116 & ~n2236;
  assign n2238 = n903 & ~n2237;
  assign n2239 = ~n822 & ~n2096;
  assign n2240 = n2103 & ~n2239;
  assign n2241 = n955 & ~n2240;
  assign n2242 = ~n2238 & ~n2241;
  assign n2243 = Ni38 & n2126;
  assign n2244 = n2128 & ~n2243;
  assign n2245 = ~n2224 & n2244;
  assign n2246 = n924 & ~n2245;
  assign n2247 = Ni38 & n2123;
  assign n2248 = n2122 & ~n2224;
  assign n2249 = ~n2247 & n2248;
  assign n2250 = n994 & ~n2249;
  assign n2251 = ~n2246 & ~n2250;
  assign n2252 = n2242 & n2251;
  assign n2253 = ~Pi20 & ~n2252;
  assign n2254 = ~n908 & ~n2140;
  assign n2255 = n2143 & ~n2254;
  assign n2256 = n1968 & ~n2255;
  assign n2257 = ~n908 & ~n2150;
  assign n2258 = n2153 & ~n2257;
  assign n2259 = n1650 & ~n2258;
  assign n2260 = ~n2256 & ~n2259;
  assign n2261 = n2134 & ~n2260;
  assign n2262 = ~n908 & ~n2163;
  assign n2263 = n2166 & ~n2262;
  assign n2264 = n1968 & ~n2263;
  assign n2265 = ~n908 & ~n2173;
  assign n2266 = n2176 & ~n2265;
  assign n2267 = n1650 & ~n2266;
  assign n2268 = ~n2264 & ~n2267;
  assign n2269 = n2159 & ~n2268;
  assign n2270 = ~n2261 & ~n2269;
  assign n2271 = ~n2253 & n2270;
  assign n2272 = ~n2235 & n2271;
  assign n2273 = n2043 & ~n2272;
  assign n2274 = n2191 & ~n2273;
  assign n2275 = ~n2216 & n2274;
  assign n2276 = n1381 & ~n2275;
  assign n2277 = ~n2210 & ~n2276;
  assign n2278 = ~n2041 & n2277;
  assign n2279 = P__cmxcl_1 & ~n579;
  assign n2280 = ~n2278 & n2279;
  assign n2281 = Ni33 & ~P__cmxcl_1;
  assign n2282 = ~Pi25 & n864;
  assign n2283 = n2037 & n2282;
  assign n2284 = n2015 & ~n2283;
  assign n2285 = Ni33 & n816;
  assign n2286 = ~n827 & n2030;
  assign n2287 = n2003 & ~n2286;
  assign n2288 = Ni40 & n2287;
  assign n2289 = ~Ni41 & ~n2031;
  assign n2290 = n2287 & ~n2289;
  assign n2291 = ~n2288 & ~n2290;
  assign n2292 = n2285 & n2291;
  assign n2293 = ~Ni34 & n2292;
  assign n2294 = n750 & n2025;
  assign n2295 = ~n2022 & ~n2294;
  assign n2296 = Ni33 & ~n2295;
  assign n2297 = ~Ni38 & ~n1060;
  assign n2298 = Ni33 & ~n2297;
  assign n2299 = n2291 & n2298;
  assign n2300 = ~n2296 & ~n2299;
  assign n2301 = ~Ni34 & ~n2300;
  assign n2302 = ~n1217 & n2037;
  assign n2303 = ~n2187 & ~n2302;
  assign n2304 = ~n2301 & n2303;
  assign n2305 = n2042 & ~n2178;
  assign n2306 = n2304 & ~n2305;
  assign n2307 = ~n2293 & n2306;
  assign n2308 = n865 & ~n2307;
  assign n2309 = n2284 & ~n2308;
  assign n2310 = n1650 & ~n2309;
  assign n2311 = ~Pi25 & n2037;
  assign n2312 = ~Pi25 & n2019;
  assign n2313 = ~n2198 & n2312;
  assign n2314 = ~n2311 & ~n2313;
  assign n2315 = n1814 & ~n2314;
  assign n2316 = Ni33 & ~n2287;
  assign n2317 = n2192 & n2316;
  assign n2318 = ~Ni34 & n2317;
  assign n2319 = Ni38 & n2316;
  assign n2320 = ~n2296 & ~n2319;
  assign n2321 = ~Ni34 & ~n2320;
  assign n2322 = n2303 & ~n2321;
  assign n2323 = ~n2318 & n2322;
  assign n2324 = ~n2199 & n2323;
  assign n2325 = n1814 & ~n2324;
  assign n2326 = n2017 & ~n2325;
  assign n2327 = n864 & n2312;
  assign n2328 = ~n2180 & n2327;
  assign n2329 = n2326 & ~n2328;
  assign n2330 = ~n2315 & n2329;
  assign n2331 = n2007 & ~n2283;
  assign n2332 = n2042 & ~n2168;
  assign n2333 = ~Ni42 & ~Ni41;
  assign n2334 = Ni44 & ~Ni43;
  assign n2335 = n872 & ~n2334;
  assign n2336 = n2003 & ~n2335;
  assign n2337 = n2333 & ~n2336;
  assign n2338 = Ni42 & n2289;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = n2287 & n2339;
  assign n2341 = ~n2288 & ~n2340;
  assign n2342 = n2285 & n2341;
  assign n2343 = ~Ni34 & n2342;
  assign n2344 = ~Ni38 & ~n893;
  assign n2345 = Ni33 & ~n2344;
  assign n2346 = n2341 & n2345;
  assign n2347 = ~n2296 & ~n2346;
  assign n2348 = ~Ni34 & ~n2347;
  assign n2349 = n2303 & ~n2348;
  assign n2350 = ~n2343 & n2349;
  assign n2351 = ~n2332 & n2350;
  assign n2352 = n865 & ~n2351;
  assign n2353 = n2331 & ~n2352;
  assign n2354 = n1968 & ~n2353;
  assign n2355 = n2330 & ~n2354;
  assign n2356 = ~n2310 & n2355;
  assign n2357 = n2159 & ~n2356;
  assign n2358 = n2158 & n2327;
  assign n2359 = ~Pi15 & ~n2358;
  assign n2360 = ~n2090 & n2327;
  assign n2361 = n2042 & ~n2082;
  assign n2362 = Ni41 & ~n2033;
  assign n2363 = n2031 & ~n2362;
  assign n2364 = n816 & ~n2363;
  assign n2365 = ~n2056 & ~n2295;
  assign n2366 = ~n2059 & ~n2363;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n2364 & n2367;
  assign n2369 = Ni33 & ~n2368;
  assign n2370 = ~Ni34 & n2369;
  assign n2371 = n2303 & ~n2370;
  assign n2372 = ~n2361 & n2371;
  assign n2373 = n994 & ~n2372;
  assign n2374 = ~n2360 & ~n2373;
  assign n2375 = ~Ni40 & n2287;
  assign n2376 = ~n2290 & ~n2375;
  assign n2377 = n2285 & n2376;
  assign n2378 = ~Ni34 & n2377;
  assign n2379 = n2042 & ~n2076;
  assign n2380 = ~Ni38 & ~n981;
  assign n2381 = Ni33 & ~n2380;
  assign n2382 = n2376 & n2381;
  assign n2383 = ~n2296 & ~n2382;
  assign n2384 = ~Ni34 & ~n2383;
  assign n2385 = n2303 & ~n2384;
  assign n2386 = ~n2379 & n2385;
  assign n2387 = ~n2378 & n2386;
  assign n2388 = n865 & n955;
  assign n2389 = ~n2387 & n2388;
  assign n2390 = n2287 & ~n2362;
  assign n2391 = Ni40 & ~n2031;
  assign n2392 = n2390 & ~n2391;
  assign n2393 = n2285 & ~n2392;
  assign n2394 = ~Ni34 & n2393;
  assign n2395 = n2042 & ~n2063;
  assign n2396 = n2381 & ~n2392;
  assign n2397 = ~n2296 & ~n2396;
  assign n2398 = ~Ni34 & ~n2397;
  assign n2399 = n2303 & ~n2398;
  assign n2400 = ~n2395 & n2399;
  assign n2401 = ~n2394 & n2400;
  assign n2402 = n903 & ~n2401;
  assign n2403 = ~Pi17 & ~n2284;
  assign n2404 = Pi20 & ~n2403;
  assign n2405 = n816 & ~n2290;
  assign n2406 = ~n2059 & ~n2290;
  assign n2407 = ~n2365 & ~n2406;
  assign n2408 = ~n2405 & n2407;
  assign n2409 = Ni33 & ~n2408;
  assign n2410 = ~Ni34 & n2409;
  assign n2411 = n2042 & ~n2087;
  assign n2412 = n2303 & ~n2411;
  assign n2413 = ~n2410 & n2412;
  assign n2414 = n865 & n924;
  assign n2415 = ~n2413 & n2414;
  assign n2416 = n2404 & ~n2415;
  assign n2417 = ~n2402 & n2416;
  assign n2418 = ~n2389 & n2417;
  assign n2419 = n2374 & n2418;
  assign n2420 = ~Pi17 & ~n2331;
  assign n2421 = ~Pi20 & ~n2420;
  assign n2422 = ~Pi16 & n1968;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = n2042 & ~n2124;
  assign n2425 = n2339 & ~n2362;
  assign n2426 = n816 & ~n2425;
  assign n2427 = n2025 & n2098;
  assign n2428 = ~n2022 & ~n2427;
  assign n2429 = ~n2101 & ~n2425;
  assign n2430 = n2428 & ~n2429;
  assign n2431 = ~n2426 & n2430;
  assign n2432 = Ni33 & ~n2431;
  assign n2433 = ~Ni34 & n2432;
  assign n2434 = n2303 & ~n2433;
  assign n2435 = ~n2424 & n2434;
  assign n2436 = n865 & ~n2435;
  assign n2437 = n2331 & ~n2436;
  assign n2438 = n994 & ~n2437;
  assign n2439 = n2042 & ~n2129;
  assign n2440 = ~n2101 & ~n2340;
  assign n2441 = n2428 & ~n2440;
  assign n2442 = n816 & ~n2340;
  assign n2443 = n2441 & ~n2442;
  assign n2444 = Ni33 & ~n2443;
  assign n2445 = ~Ni34 & n2444;
  assign n2446 = n2303 & ~n2445;
  assign n2447 = ~n2439 & n2446;
  assign n2448 = n2414 & ~n2447;
  assign n2449 = ~n2340 & ~n2375;
  assign n2450 = ~n2362 & ~n2449;
  assign n2451 = n2285 & ~n2450;
  assign n2452 = ~Ni34 & n2451;
  assign n2453 = ~Ni38 & ~n911;
  assign n2454 = Ni33 & ~n2453;
  assign n2455 = ~n2450 & n2454;
  assign n2456 = ~n2296 & ~n2455;
  assign n2457 = ~Ni34 & ~n2456;
  assign n2458 = n2303 & ~n2457;
  assign n2459 = n2042 & ~n2118;
  assign n2460 = n2458 & ~n2459;
  assign n2461 = ~n2452 & n2460;
  assign n2462 = n865 & n903;
  assign n2463 = ~n2461 & n2462;
  assign n2464 = ~n2448 & ~n2463;
  assign n2465 = n2285 & n2449;
  assign n2466 = ~Ni34 & n2465;
  assign n2467 = n2042 & ~n2105;
  assign n2468 = n2449 & n2454;
  assign n2469 = ~n2296 & ~n2468;
  assign n2470 = ~Ni34 & ~n2469;
  assign n2471 = n2303 & ~n2470;
  assign n2472 = ~n2467 & n2471;
  assign n2473 = ~n2466 & n2472;
  assign n2474 = n2388 & ~n2473;
  assign n2475 = ~n2132 & n2327;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n2464 & n2476;
  assign n2478 = ~n2438 & n2477;
  assign n2479 = ~n2423 & n2478;
  assign n2480 = ~n2419 & ~n2479;
  assign n2481 = ~Ni40 & ~n2031;
  assign n2482 = n2390 & ~n2481;
  assign n2483 = n2298 & ~n2482;
  assign n2484 = ~n2296 & ~n2483;
  assign n2485 = ~Ni34 & ~n2484;
  assign n2486 = n2303 & ~n2485;
  assign n2487 = n2285 & ~n2482;
  assign n2488 = ~Ni34 & n2487;
  assign n2489 = n2042 & ~n2155;
  assign n2490 = ~n2488 & ~n2489;
  assign n2491 = n2486 & n2490;
  assign n2492 = n2284 & n2491;
  assign n2493 = n1650 & ~n2492;
  assign n2494 = ~n2341 & ~n2362;
  assign n2495 = n2285 & ~n2494;
  assign n2496 = ~Ni34 & n2495;
  assign n2497 = n2345 & ~n2494;
  assign n2498 = ~n2296 & ~n2497;
  assign n2499 = ~Ni34 & ~n2498;
  assign n2500 = n2303 & ~n2499;
  assign n2501 = n2042 & ~n2145;
  assign n2502 = n2500 & ~n2501;
  assign n2503 = ~n2496 & n2502;
  assign n2504 = n865 & ~n2503;
  assign n2505 = n2331 & ~n2504;
  assign n2506 = n1968 & ~n2505;
  assign n2507 = Ni33 & ~n2390;
  assign n2508 = n2192 & n2507;
  assign n2509 = ~Ni34 & n2508;
  assign n2510 = Ni38 & n2507;
  assign n2511 = ~n2296 & ~n2510;
  assign n2512 = ~Ni34 & ~n2511;
  assign n2513 = n2303 & ~n2512;
  assign n2514 = ~n2509 & n2513;
  assign n2515 = ~n2204 & n2514;
  assign n2516 = n1814 & ~n2515;
  assign n2517 = n2017 & ~n2516;
  assign n2518 = n2203 & ~n2311;
  assign n2519 = n2315 & ~n2518;
  assign n2520 = n2517 & ~n2519;
  assign n2521 = ~n2506 & n2520;
  assign n2522 = ~n2493 & n2521;
  assign n2523 = n2134 & ~n2522;
  assign n2524 = ~n2480 & ~n2523;
  assign n2525 = n2359 & n2524;
  assign n2526 = ~n2357 & n2525;
  assign n2527 = ~n2234 & n2327;
  assign n2528 = n2404 & ~n2527;
  assign n2529 = n2042 & ~n2218;
  assign n2530 = n2399 & ~n2529;
  assign n2531 = n903 & ~n2530;
  assign n2532 = n2042 & ~n2221;
  assign n2533 = n2385 & ~n2532;
  assign n2534 = n2388 & ~n2533;
  assign n2535 = ~n2531 & ~n2534;
  assign n2536 = n2042 & ~n2231;
  assign n2537 = Ni36 & n2294;
  assign n2538 = n2367 & ~n2537;
  assign n2539 = Ni38 & n2364;
  assign n2540 = n2538 & ~n2539;
  assign n2541 = Ni33 & ~n2540;
  assign n2542 = ~Ni34 & n2541;
  assign n2543 = n2303 & ~n2542;
  assign n2544 = ~n2536 & n2543;
  assign n2545 = n994 & ~n2544;
  assign n2546 = Ni38 & n2405;
  assign n2547 = n2407 & ~n2546;
  assign n2548 = ~n2537 & n2547;
  assign n2549 = Ni33 & ~n2548;
  assign n2550 = ~Ni34 & n2549;
  assign n2551 = n2042 & ~n2227;
  assign n2552 = n2303 & ~n2551;
  assign n2553 = ~n2550 & n2552;
  assign n2554 = n2414 & ~n2553;
  assign n2555 = ~n2545 & ~n2554;
  assign n2556 = n2535 & n2555;
  assign n2557 = n2528 & n2556;
  assign n2558 = n2042 & ~n2240;
  assign n2559 = n2471 & ~n2558;
  assign n2560 = n955 & ~n2559;
  assign n2561 = n2042 & ~n2245;
  assign n2562 = Ni38 & n2442;
  assign n2563 = n2441 & ~n2562;
  assign n2564 = ~n2537 & n2563;
  assign n2565 = Ni33 & ~n2564;
  assign n2566 = ~Ni34 & n2565;
  assign n2567 = n2303 & ~n2566;
  assign n2568 = ~n2561 & n2567;
  assign n2569 = n924 & ~n2568;
  assign n2570 = n2042 & ~n2237;
  assign n2571 = n2458 & ~n2570;
  assign n2572 = n903 & ~n2571;
  assign n2573 = n2042 & ~n2249;
  assign n2574 = Ni38 & n2426;
  assign n2575 = n2430 & ~n2537;
  assign n2576 = ~n2574 & n2575;
  assign n2577 = Ni33 & ~n2576;
  assign n2578 = ~Ni34 & n2577;
  assign n2579 = n2303 & ~n2578;
  assign n2580 = ~n2573 & n2579;
  assign n2581 = n994 & ~n2580;
  assign n2582 = ~n2572 & ~n2581;
  assign n2583 = ~n2569 & n2582;
  assign n2584 = ~n2560 & n2583;
  assign n2585 = n865 & ~n2584;
  assign n2586 = ~n2252 & n2327;
  assign n2587 = n2421 & ~n2586;
  assign n2588 = ~n2585 & n2587;
  assign n2589 = ~n2557 & ~n2588;
  assign n2590 = ~n2270 & n2327;
  assign n2591 = ~n1528 & n2212;
  assign n2592 = n2312 & ~n2591;
  assign n2593 = ~n2195 & n2592;
  assign n2594 = ~n2311 & ~n2593;
  assign n2595 = n1030 & ~n2594;
  assign n2596 = Pi15 & ~n2595;
  assign n2597 = ~n2590 & n2596;
  assign n2598 = n2042 & ~n2266;
  assign n2599 = n2304 & ~n2598;
  assign n2600 = n865 & ~n2599;
  assign n2601 = n2284 & ~n2600;
  assign n2602 = n1650 & ~n2601;
  assign n2603 = ~n2211 & n2322;
  assign n2604 = n1814 & ~n2603;
  assign n2605 = n2017 & ~n2604;
  assign n2606 = n2042 & ~n2263;
  assign n2607 = n2349 & ~n2606;
  assign n2608 = n865 & ~n2607;
  assign n2609 = n2331 & ~n2608;
  assign n2610 = n1968 & ~n2609;
  assign n2611 = n2605 & ~n2610;
  assign n2612 = ~n2602 & n2611;
  assign n2613 = n2159 & ~n2612;
  assign n2614 = n2042 & ~n2255;
  assign n2615 = n2500 & ~n2614;
  assign n2616 = n865 & ~n2615;
  assign n2617 = n2331 & ~n2616;
  assign n2618 = n1968 & ~n2617;
  assign n2619 = n2211 & ~n2212;
  assign n2620 = n2513 & ~n2619;
  assign n2621 = n1814 & ~n2620;
  assign n2622 = n2017 & ~n2621;
  assign n2623 = n2042 & ~n2258;
  assign n2624 = n2486 & ~n2623;
  assign n2625 = n2284 & n2624;
  assign n2626 = n1650 & ~n2625;
  assign n2627 = n2622 & ~n2626;
  assign n2628 = ~n2618 & n2627;
  assign n2629 = n2134 & ~n2628;
  assign n2630 = ~n2613 & ~n2629;
  assign n2631 = n2597 & n2630;
  assign n2632 = ~n2589 & n2631;
  assign n2633 = n570 & ~n2632;
  assign n2634 = ~n2526 & n2633;
  assign n2635 = ~Ni14 & ~Ni13;
  assign n2636 = n582 & n2635;
  assign n2637 = ~n1995 & ~n2028;
  assign n2638 = n2300 & n2637;
  assign n2639 = n950 & ~n2638;
  assign n2640 = ~n2038 & n2282;
  assign n2641 = n2017 & ~n2640;
  assign n2642 = n2347 & n2637;
  assign n2643 = n868 & ~n2642;
  assign n2644 = n2641 & ~n2643;
  assign n2645 = ~n2639 & n2644;
  assign n2646 = n1035 & ~n2645;
  assign n2647 = n2383 & n2637;
  assign n2648 = n950 & ~n2647;
  assign n2649 = n2469 & n2637;
  assign n2650 = n868 & ~n2649;
  assign n2651 = n2641 & ~n2650;
  assign n2652 = ~n2648 & n2651;
  assign n2653 = n955 & ~n2652;
  assign n2654 = n730 & ~n2641;
  assign n2655 = Pi15 & ~n2654;
  assign n2656 = ~n2577 & n2637;
  assign n2657 = n868 & ~n2656;
  assign n2658 = ~n2541 & n2637;
  assign n2659 = n950 & ~n2658;
  assign n2660 = n2641 & ~n2659;
  assign n2661 = ~n2657 & n2660;
  assign n2662 = n994 & ~n2661;
  assign n2663 = n2655 & ~n2662;
  assign n2664 = ~n2653 & n2663;
  assign n2665 = n2320 & n2637;
  assign n2666 = n744 & ~n2665;
  assign n2667 = n2511 & n2637;
  assign n2668 = n731 & ~n2667;
  assign n2669 = ~n2666 & ~n2668;
  assign n2670 = n865 & ~n2669;
  assign n2671 = n2498 & n2637;
  assign n2672 = n868 & ~n2671;
  assign n2673 = n2484 & n2637;
  assign n2674 = n950 & ~n2673;
  assign n2675 = n2641 & ~n2674;
  assign n2676 = ~n2672 & n2675;
  assign n2677 = n869 & ~n2676;
  assign n2678 = ~n2670 & ~n2677;
  assign n2679 = ~n2565 & n2637;
  assign n2680 = n868 & ~n2679;
  assign n2681 = ~n2549 & n2637;
  assign n2682 = n950 & ~n2681;
  assign n2683 = n2641 & ~n2682;
  assign n2684 = ~n2680 & n2683;
  assign n2685 = n924 & ~n2684;
  assign n2686 = n2456 & n2637;
  assign n2687 = n868 & ~n2686;
  assign n2688 = n2397 & n2637;
  assign n2689 = n950 & ~n2688;
  assign n2690 = n2641 & ~n2689;
  assign n2691 = ~n2687 & n2690;
  assign n2692 = n903 & ~n2691;
  assign n2693 = ~n2685 & ~n2692;
  assign n2694 = n2678 & n2693;
  assign n2695 = n2664 & n2694;
  assign n2696 = ~n2393 & n2688;
  assign n2697 = n950 & ~n2696;
  assign n2698 = ~n2451 & n2686;
  assign n2699 = n868 & ~n2698;
  assign n2700 = n2641 & ~n2699;
  assign n2701 = ~n2697 & n2700;
  assign n2702 = n903 & ~n2701;
  assign n2703 = n868 & n2342;
  assign n2704 = n950 & n2292;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = n1035 & ~n2705;
  assign n2707 = ~n2508 & n2667;
  assign n2708 = n731 & ~n2707;
  assign n2709 = n744 & n2317;
  assign n2710 = ~n2666 & ~n2709;
  assign n2711 = ~n2708 & n2710;
  assign n2712 = n865 & ~n2711;
  assign n2713 = ~n2706 & ~n2712;
  assign n2714 = ~Pi15 & ~n2654;
  assign n2715 = ~n2432 & n2637;
  assign n2716 = n868 & ~n2715;
  assign n2717 = ~n2369 & n2637;
  assign n2718 = n950 & ~n2717;
  assign n2719 = n2641 & ~n2718;
  assign n2720 = ~n2716 & n2719;
  assign n2721 = n994 & ~n2720;
  assign n2722 = n2714 & ~n2721;
  assign n2723 = n2713 & n2722;
  assign n2724 = ~n2495 & n2671;
  assign n2725 = n868 & ~n2724;
  assign n2726 = ~n2487 & n2673;
  assign n2727 = n950 & ~n2726;
  assign n2728 = n2641 & ~n2727;
  assign n2729 = ~n2725 & n2728;
  assign n2730 = n869 & ~n2729;
  assign n2731 = ~n2377 & n2647;
  assign n2732 = n950 & ~n2731;
  assign n2733 = ~n2465 & n2649;
  assign n2734 = n868 & ~n2733;
  assign n2735 = n2641 & ~n2734;
  assign n2736 = ~n2732 & n2735;
  assign n2737 = n955 & ~n2736;
  assign n2738 = ~n2444 & n2637;
  assign n2739 = n868 & ~n2738;
  assign n2740 = ~n2409 & n2637;
  assign n2741 = n950 & ~n2740;
  assign n2742 = n2641 & ~n2741;
  assign n2743 = ~n2739 & n2742;
  assign n2744 = n924 & ~n2743;
  assign n2745 = ~n2737 & ~n2744;
  assign n2746 = ~n2730 & n2745;
  assign n2747 = n2723 & n2746;
  assign n2748 = ~n2702 & n2747;
  assign n2749 = ~n2695 & ~n2748;
  assign n2750 = ~n2646 & ~n2749;
  assign n2751 = n2636 & ~n2750;
  assign n2752 = ~n2028 & ~n2302;
  assign n2753 = ~n2433 & n2752;
  assign n2754 = n868 & ~n2753;
  assign n2755 = ~n2370 & n2752;
  assign n2756 = n950 & ~n2755;
  assign n2757 = n2641 & ~n2756;
  assign n2758 = ~n2754 & n2757;
  assign n2759 = n994 & ~n2758;
  assign n2760 = ~n2321 & n2752;
  assign n2761 = ~n2318 & n2760;
  assign n2762 = n744 & ~n2761;
  assign n2763 = ~n2512 & n2752;
  assign n2764 = ~n2509 & n2763;
  assign n2765 = n731 & ~n2764;
  assign n2766 = ~n2762 & ~n2765;
  assign n2767 = n865 & ~n2766;
  assign n2768 = ~n2759 & ~n2767;
  assign n2769 = ~n2499 & n2752;
  assign n2770 = ~n2496 & n2769;
  assign n2771 = n868 & ~n2770;
  assign n2772 = ~n2485 & n2752;
  assign n2773 = ~n2488 & n2772;
  assign n2774 = n950 & ~n2773;
  assign n2775 = n2641 & ~n2774;
  assign n2776 = ~n2771 & n2775;
  assign n2777 = n869 & ~n2776;
  assign n2778 = n2768 & ~n2777;
  assign n2779 = ~n2398 & n2752;
  assign n2780 = ~n2394 & n2779;
  assign n2781 = n950 & ~n2780;
  assign n2782 = ~n2457 & n2752;
  assign n2783 = ~n2452 & n2782;
  assign n2784 = n868 & ~n2783;
  assign n2785 = n2641 & ~n2784;
  assign n2786 = ~n2781 & n2785;
  assign n2787 = n903 & ~n2786;
  assign n2788 = ~n2445 & n2752;
  assign n2789 = n868 & ~n2788;
  assign n2790 = ~n2410 & n2752;
  assign n2791 = n950 & ~n2790;
  assign n2792 = n2641 & ~n2791;
  assign n2793 = ~n2789 & n2792;
  assign n2794 = n924 & ~n2793;
  assign n2795 = ~n2470 & n2752;
  assign n2796 = ~n2466 & n2795;
  assign n2797 = n868 & ~n2796;
  assign n2798 = ~n2384 & n2752;
  assign n2799 = ~n2378 & n2798;
  assign n2800 = n950 & ~n2799;
  assign n2801 = n2641 & ~n2800;
  assign n2802 = ~n2797 & n2801;
  assign n2803 = n955 & ~n2802;
  assign n2804 = n2714 & ~n2803;
  assign n2805 = ~n2794 & n2804;
  assign n2806 = ~n2787 & n2805;
  assign n2807 = ~n2348 & n2752;
  assign n2808 = ~n2343 & n2807;
  assign n2809 = n868 & ~n2808;
  assign n2810 = ~n2301 & n2752;
  assign n2811 = ~n2293 & n2810;
  assign n2812 = n950 & ~n2811;
  assign n2813 = n2641 & ~n2812;
  assign n2814 = ~n2809 & n2813;
  assign n2815 = n1035 & ~n2814;
  assign n2816 = n2806 & ~n2815;
  assign n2817 = n2778 & n2816;
  assign n2818 = ~n2542 & n2752;
  assign n2819 = n950 & ~n2818;
  assign n2820 = ~n2578 & n2752;
  assign n2821 = n868 & ~n2820;
  assign n2822 = n2641 & ~n2821;
  assign n2823 = ~n2819 & n2822;
  assign n2824 = n994 & ~n2823;
  assign n2825 = n868 & ~n2769;
  assign n2826 = n950 & ~n2772;
  assign n2827 = n2641 & ~n2826;
  assign n2828 = ~n2825 & n2827;
  assign n2829 = n869 & ~n2828;
  assign n2830 = n744 & ~n2760;
  assign n2831 = n731 & ~n2763;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n865 & ~n2832;
  assign n2834 = ~n2829 & ~n2833;
  assign n2835 = n2655 & n2834;
  assign n2836 = ~n2566 & n2752;
  assign n2837 = n868 & ~n2836;
  assign n2838 = ~n2550 & n2752;
  assign n2839 = n950 & ~n2838;
  assign n2840 = n2641 & ~n2839;
  assign n2841 = ~n2837 & n2840;
  assign n2842 = n924 & ~n2841;
  assign n2843 = n950 & ~n2779;
  assign n2844 = n868 & ~n2782;
  assign n2845 = n2641 & ~n2844;
  assign n2846 = ~n2843 & n2845;
  assign n2847 = n903 & ~n2846;
  assign n2848 = n868 & ~n2807;
  assign n2849 = n950 & ~n2810;
  assign n2850 = n2641 & ~n2849;
  assign n2851 = ~n2848 & n2850;
  assign n2852 = n1035 & ~n2851;
  assign n2853 = n950 & ~n2798;
  assign n2854 = n868 & ~n2795;
  assign n2855 = n2641 & ~n2854;
  assign n2856 = ~n2853 & n2855;
  assign n2857 = n955 & ~n2856;
  assign n2858 = ~n2852 & ~n2857;
  assign n2859 = ~n2847 & n2858;
  assign n2860 = ~n2842 & n2859;
  assign n2861 = n2835 & n2860;
  assign n2862 = ~n2824 & n2861;
  assign n2863 = ~n2817 & ~n2862;
  assign n2864 = ~n569 & n2863;
  assign n2865 = ~n2751 & ~n2864;
  assign n2866 = ~n2634 & n2865;
  assign n2867 = ~Ni10 & ~n2866;
  assign n2868 = n1625 & ~n2724;
  assign n2869 = n1643 & ~n2726;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = n1610 & ~n2870;
  assign n2872 = n1610 & n1814;
  assign n2873 = ~n2707 & n2872;
  assign n2874 = ~n2871 & ~n2873;
  assign n2875 = n1643 & ~n2673;
  assign n2876 = n1814 & ~n2667;
  assign n2877 = n1625 & ~n2671;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = ~n2875 & n2878;
  assign n2880 = n1178 & ~n2879;
  assign n2881 = ~Pi15 & n2342;
  assign n2882 = n2642 & ~n2881;
  assign n2883 = n1625 & ~n2882;
  assign n2884 = n1814 & ~n2665;
  assign n2885 = ~Pi15 & n2292;
  assign n2886 = n2638 & ~n2885;
  assign n2887 = n1643 & ~n2886;
  assign n2888 = ~n2884 & ~n2887;
  assign n2889 = ~n2883 & n2888;
  assign n2890 = Pi16 & ~n2889;
  assign n2891 = n1878 & n2317;
  assign n2892 = Pi17 & n2017;
  assign n2893 = ~n2891 & n2892;
  assign n2894 = ~n2890 & n2893;
  assign n2895 = ~n2880 & n2894;
  assign n2896 = n2874 & n2895;
  assign n2897 = n1611 & ~n2696;
  assign n2898 = n1643 & ~n2717;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = n1636 & ~n2698;
  assign n2901 = n1625 & ~n2715;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = n2899 & n2902;
  assign n2904 = n2017 & n2903;
  assign n2905 = n1610 & ~n2904;
  assign n2906 = n1625 & ~n2679;
  assign n2907 = n1611 & ~n2647;
  assign n2908 = n1636 & ~n2649;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = n1643 & ~n2681;
  assign n2911 = n2017 & ~n2910;
  assign n2912 = n2909 & n2911;
  assign n2913 = ~n2906 & n2912;
  assign n2914 = n1769 & ~n2913;
  assign n2915 = n1611 & ~n2688;
  assign n2916 = n1643 & ~n2658;
  assign n2917 = n2017 & ~n2916;
  assign n2918 = n1625 & ~n2656;
  assign n2919 = n1636 & ~n2686;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n2917 & n2920;
  assign n2922 = ~n2915 & n2921;
  assign n2923 = n1178 & ~n2922;
  assign n2924 = n1636 & ~n2733;
  assign n2925 = n1611 & ~n2731;
  assign n2926 = n2017 & ~n2925;
  assign n2927 = n1643 & ~n2740;
  assign n2928 = n1625 & ~n2738;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2926 & n2929;
  assign n2931 = ~n2924 & n2930;
  assign n2932 = n1672 & ~n2931;
  assign n2933 = ~Pi17 & ~n2932;
  assign n2934 = ~n2923 & n2933;
  assign n2935 = ~n2914 & n2934;
  assign n2936 = ~n2905 & n2935;
  assign n2937 = n2636 & ~n2936;
  assign n2938 = ~n2896 & n2937;
  assign n2939 = n1814 & ~n2763;
  assign n2940 = n1643 & ~n2772;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n1625 & ~n2769;
  assign n2943 = n2017 & ~n2942;
  assign n2944 = n2941 & n2943;
  assign n2945 = n1178 & ~n2944;
  assign n2946 = n1643 & ~n2773;
  assign n2947 = n1625 & ~n2770;
  assign n2948 = n2017 & ~n2947;
  assign n2949 = ~n2946 & n2948;
  assign n2950 = n1610 & ~n2949;
  assign n2951 = ~n2764 & n2872;
  assign n2952 = n1878 & ~n2761;
  assign n2953 = Pi17 & ~n2952;
  assign n2954 = ~n2951 & n2953;
  assign n2955 = n1625 & ~n2808;
  assign n2956 = n1643 & ~n2811;
  assign n2957 = n2017 & ~n2956;
  assign n2958 = ~n2955 & n2957;
  assign n2959 = n1672 & ~n2958;
  assign n2960 = n1814 & ~n2760;
  assign n2961 = n1625 & ~n2807;
  assign n2962 = n1643 & ~n2810;
  assign n2963 = n2017 & ~n2962;
  assign n2964 = ~n2961 & n2963;
  assign n2965 = ~n2960 & n2964;
  assign n2966 = n1769 & ~n2965;
  assign n2967 = ~n2959 & ~n2966;
  assign n2968 = n2954 & n2967;
  assign n2969 = ~n2950 & n2968;
  assign n2970 = ~n2945 & n2969;
  assign n2971 = n1611 & ~n2779;
  assign n2972 = n1625 & ~n2820;
  assign n2973 = n2017 & ~n2972;
  assign n2974 = n1643 & ~n2818;
  assign n2975 = n1636 & ~n2782;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = n2973 & n2976;
  assign n2978 = ~n2971 & n2977;
  assign n2979 = n1178 & ~n2978;
  assign n2980 = n1643 & ~n2790;
  assign n2981 = n1611 & ~n2799;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = n1636 & ~n2796;
  assign n2984 = n1625 & ~n2788;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = n2982 & n2985;
  assign n2987 = n2017 & n2986;
  assign n2988 = n1672 & ~n2987;
  assign n2989 = n1643 & ~n2838;
  assign n2990 = n1625 & ~n2836;
  assign n2991 = n1636 & ~n2795;
  assign n2992 = n1611 & ~n2798;
  assign n2993 = n2017 & ~n2992;
  assign n2994 = ~n2991 & n2993;
  assign n2995 = ~n2990 & n2994;
  assign n2996 = ~n2989 & n2995;
  assign n2997 = n1769 & ~n2996;
  assign n2998 = ~n2988 & ~n2997;
  assign n2999 = n1636 & ~n2783;
  assign n3000 = n1625 & ~n2753;
  assign n3001 = n2017 & ~n3000;
  assign n3002 = n1611 & ~n2780;
  assign n3003 = n1643 & ~n2755;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = n3001 & n3004;
  assign n3006 = ~n2999 & n3005;
  assign n3007 = n1610 & ~n3006;
  assign n3008 = ~Pi17 & ~n3007;
  assign n3009 = n2998 & n3008;
  assign n3010 = ~n2979 & n3009;
  assign n3011 = ~n569 & ~n3010;
  assign n3012 = ~n2970 & n3011;
  assign n3013 = n1625 & ~n2351;
  assign n3014 = n1643 & ~n2307;
  assign n3015 = n2326 & ~n3014;
  assign n3016 = ~n3013 & n3015;
  assign n3017 = n1672 & ~n3016;
  assign n3018 = n1625 & ~n2503;
  assign n3019 = n1643 & ~n2491;
  assign n3020 = n2517 & ~n3019;
  assign n3021 = ~n3018 & n3020;
  assign n3022 = n1610 & ~n3021;
  assign n3023 = n1643 & ~n2624;
  assign n3024 = n1625 & ~n2615;
  assign n3025 = n2622 & ~n3024;
  assign n3026 = ~n3023 & n3025;
  assign n3027 = n1178 & ~n3026;
  assign n3028 = n1643 & ~n2599;
  assign n3029 = n1625 & ~n2607;
  assign n3030 = n2605 & ~n3029;
  assign n3031 = ~n3028 & n3030;
  assign n3032 = n1769 & ~n3031;
  assign n3033 = ~n3027 & ~n3032;
  assign n3034 = ~n3022 & n3033;
  assign n3035 = ~n3017 & n3034;
  assign n3036 = Pi17 & n3035;
  assign n3037 = n1625 & ~n2435;
  assign n3038 = n1643 & ~n2372;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = n1636 & ~n2461;
  assign n3041 = n1611 & ~n2401;
  assign n3042 = ~n3040 & ~n3041;
  assign n3043 = n3039 & n3042;
  assign n3044 = n2017 & n3043;
  assign n3045 = n1610 & ~n3044;
  assign n3046 = n1643 & ~n2544;
  assign n3047 = n1636 & ~n2571;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n1625 & ~n2580;
  assign n3050 = n1611 & ~n2530;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n3048 & n3051;
  assign n3053 = n2017 & n3052;
  assign n3054 = n1178 & ~n3053;
  assign n3055 = ~n3045 & ~n3054;
  assign n3056 = n1636 & ~n2473;
  assign n3057 = n1611 & ~n2387;
  assign n3058 = n1625 & ~n2447;
  assign n3059 = n2017 & ~n3058;
  assign n3060 = n1643 & ~n2413;
  assign n3061 = n3059 & ~n3060;
  assign n3062 = ~n3057 & n3061;
  assign n3063 = ~n3056 & n3062;
  assign n3064 = n1672 & ~n3063;
  assign n3065 = n1625 & ~n2568;
  assign n3066 = n1636 & ~n2559;
  assign n3067 = n2017 & ~n3066;
  assign n3068 = n1611 & ~n2533;
  assign n3069 = n1643 & ~n2553;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n3067 & n3070;
  assign n3072 = ~n3065 & n3071;
  assign n3073 = n1769 & ~n3072;
  assign n3074 = ~Pi17 & ~n3073;
  assign n3075 = ~n3064 & n3074;
  assign n3076 = n3055 & n3075;
  assign n3077 = n570 & ~n3076;
  assign n3078 = ~n3036 & n3077;
  assign n3079 = ~n3012 & ~n3078;
  assign n3080 = ~n2938 & n3079;
  assign n3081 = Ni10 & ~n3080;
  assign n3082 = ~n2867 & ~n3081;
  assign n3083 = n580 & ~n3082;
  assign n3084 = ~n2281 & ~n3083;
  assign n1007_1 = n2280 | ~n3084;
  assign n3086 = P__cmxcl_1 & ~n775;
  assign n3087 = ~n671 & ~n679;
  assign n3088 = Ni32 & Ni31;
  assign n3089 = ~n727 & ~n3088;
  assign n3090 = ~Pi21 & ~n3089;
  assign n3091 = ~Ni45 & n870;
  assign n3092 = ~n706 & ~n3088;
  assign n3093 = ~n3091 & n3092;
  assign n3094 = ~n727 & n3093;
  assign n3095 = n2000 & ~n3094;
  assign n3096 = ~Pi27 & Ni30;
  assign n3097 = n716 & ~n3096;
  assign n3098 = ~n3095 & ~n3097;
  assign n3099 = ~n3090 & n3098;
  assign n3100 = ~Ni32 & ~n3091;
  assign n3101 = n2000 & ~n3100;
  assign n3102 = ~Pi26 & n716;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n677 & ~n3103;
  assign n3105 = n3099 & ~n3104;
  assign n3106 = ~Ni47 & ~n874;
  assign n3107 = ~Ni45 & ~n3106;
  assign n3108 = ~Ni47 & n873;
  assign n3109 = n870 & ~n3108;
  assign n3110 = n3107 & n3109;
  assign n3111 = Pi27 & Ni32;
  assign n3112 = Ni32 & ~n855;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3110 & n3113;
  assign n3115 = ~Pi26 & Ni32;
  assign n3116 = n3114 & ~n3115;
  assign n3117 = n864 & ~n3116;
  assign n3118 = n3105 & ~n3117;
  assign n3119 = Ni11 & ~n3118;
  assign n3120 = ~n3087 & ~n3119;
  assign n3121 = ~Ni33 & Ni30;
  assign n3122 = ~Ni31 & n3121;
  assign n3123 = n716 & ~n3122;
  assign n3124 = ~n790 & n3093;
  assign n3125 = n3101 & ~n3124;
  assign n3126 = ~n3123 & ~n3125;
  assign n3127 = n3092 & ~n3110;
  assign n3128 = ~n790 & n3127;
  assign n3129 = n864 & ~n3128;
  assign n3130 = n3126 & ~n3129;
  assign n3131 = ~n716 & ~n3101;
  assign n3132 = n864 & n3110;
  assign n3133 = Ni32 & n864;
  assign n3134 = ~n3132 & ~n3133;
  assign n3135 = n3131 & n3134;
  assign n3136 = ~n691 & ~n3135;
  assign n3137 = n3130 & ~n3136;
  assign n3138 = ~n3120 & ~n3137;
  assign n3139 = Pi27 & n3094;
  assign n3140 = n3101 & ~n3139;
  assign n3141 = Pi27 & n855;
  assign n3142 = n716 & ~n3141;
  assign n3143 = ~n3140 & ~n3142;
  assign n3144 = n3133 & ~n3141;
  assign n3145 = ~n3132 & ~n3144;
  assign n3146 = n3143 & n3145;
  assign n3147 = ~n691 & n3146;
  assign n3148 = n2000 & ~n3093;
  assign n3149 = n3092 & ~n3148;
  assign n3150 = n726 & n769;
  assign n3151 = n3149 & ~n3150;
  assign n3152 = ~n3132 & n3151;
  assign n3153 = n678 & ~n3152;
  assign n3154 = n678 & ~n691;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3147 & ~n3155;
  assign n3157 = n2000 & ~n3124;
  assign n3158 = ~n3129 & ~n3157;
  assign n3159 = Pi26 & ~Pi24;
  assign n3160 = ~n3158 & n3159;
  assign n3161 = Ni32 & n3141;
  assign n3162 = n3127 & ~n3161;
  assign n3163 = n864 & ~n3162;
  assign n3164 = n3149 & ~n3163;
  assign n3165 = ~n3161 & n3164;
  assign n3166 = n790 & n3159;
  assign n3167 = n3165 & ~n3166;
  assign n3168 = ~Pi22 & n3161;
  assign n3169 = ~n3148 & ~n3168;
  assign n3170 = Pi21 & n3169;
  assign n3171 = ~n3163 & n3170;
  assign n3172 = ~n3167 & ~n3171;
  assign n3173 = ~n3160 & ~n3172;
  assign n3174 = Pi23 & ~n3173;
  assign n3175 = ~n604 & n3101;
  assign n3176 = Pi26 & n716;
  assign n3177 = n3099 & ~n3176;
  assign n3178 = ~n3175 & n3177;
  assign n3179 = Pi26 & Ni32;
  assign n3180 = n3114 & ~n3179;
  assign n3181 = n864 & ~n3180;
  assign n3182 = n3178 & ~n3181;
  assign n3183 = ~n691 & ~n3182;
  assign n3184 = ~n3174 & ~n3183;
  assign n3185 = n2635 & ~n3184;
  assign n3186 = ~n3156 & ~n3185;
  assign n3187 = n670 & ~n3186;
  assign n3188 = Ni41 & ~n3107;
  assign n3189 = ~Ni32 & n3188;
  assign n3190 = ~Ni38 & ~n3107;
  assign n3191 = ~Ni47 & Ni43;
  assign n3192 = ~Ni45 & ~n3108;
  assign n3193 = ~n3191 & n3192;
  assign n3194 = ~n3190 & n3193;
  assign n3195 = Ni36 & n3193;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = n870 & ~n3196;
  assign n3198 = ~n706 & ~n3197;
  assign n3199 = ~n18 & ~n3198;
  assign n3200 = ~n700 & ~n3199;
  assign n3201 = ~n3189 & ~n3200;
  assign n3202 = ~n706 & n3188;
  assign n3203 = ~n2018 & ~n3110;
  assign n3204 = ~n3196 & ~n3203;
  assign n3205 = ~n706 & ~n3204;
  assign n3206 = ~n3202 & ~n3205;
  assign n3207 = ~n3201 & ~n3206;
  assign n3208 = ~n691 & n1030;
  assign n3209 = ~n3207 & n3208;
  assign n3210 = ~n691 & ~n3131;
  assign n3211 = n3126 & ~n3210;
  assign n3212 = Ni32 & ~n3122;
  assign n3213 = n3188 & ~n3212;
  assign n3214 = n3211 & n3213;
  assign n3215 = n908 & n3190;
  assign n3216 = ~Ni47 & n2333;
  assign n3217 = ~n2029 & n3216;
  assign n3218 = n891 & n3190;
  assign n3219 = n3193 & ~n3218;
  assign n3220 = ~n3217 & n3219;
  assign n3221 = ~Ni40 & n3219;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~n3215 & ~n3222;
  assign n3224 = n870 & n3223;
  assign n3225 = ~n706 & ~n3224;
  assign n3226 = ~n18 & ~n3225;
  assign n3227 = ~n3203 & n3223;
  assign n3228 = ~n706 & ~n3227;
  assign n3229 = ~n790 & ~n3088;
  assign n3230 = n3228 & n3229;
  assign n3231 = ~n3226 & n3230;
  assign n3232 = n691 & n949;
  assign n3233 = ~n3231 & n3232;
  assign n3234 = n938 & n3190;
  assign n3235 = n3193 & ~n3234;
  assign n3236 = ~n2334 & n3216;
  assign n3237 = n3235 & ~n3236;
  assign n3238 = ~Ni40 & n3235;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3215 & ~n3239;
  assign n3241 = n870 & n3240;
  assign n3242 = ~n706 & ~n3241;
  assign n3243 = ~n18 & ~n3242;
  assign n3244 = ~n3203 & n3240;
  assign n3245 = ~n706 & ~n3244;
  assign n3246 = n3229 & n3245;
  assign n3247 = ~n3243 & n3246;
  assign n3248 = n691 & n867;
  assign n3249 = ~n3247 & n3248;
  assign n3250 = n3211 & ~n3249;
  assign n3251 = ~n3233 & n3250;
  assign n3252 = ~n3214 & ~n3251;
  assign n3253 = ~n700 & ~n3226;
  assign n3254 = ~n3189 & ~n3253;
  assign n3255 = ~n3202 & ~n3228;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = ~n691 & n949;
  assign n3258 = ~n3256 & n3257;
  assign n3259 = ~n700 & ~n3243;
  assign n3260 = ~n3189 & ~n3259;
  assign n3261 = ~n3202 & ~n3245;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = ~n691 & n867;
  assign n3264 = ~n3262 & n3263;
  assign n3265 = ~n3258 & ~n3264;
  assign n3266 = ~n3252 & n3265;
  assign n3267 = n738 & ~n3266;
  assign n3268 = n870 & n3237;
  assign n3269 = ~n706 & ~n3268;
  assign n3270 = ~n18 & ~n3269;
  assign n3271 = ~n3203 & n3237;
  assign n3272 = ~n706 & ~n3271;
  assign n3273 = n3229 & n3272;
  assign n3274 = ~n3270 & n3273;
  assign n3275 = n3248 & ~n3274;
  assign n3276 = n870 & n3220;
  assign n3277 = ~n706 & ~n3276;
  assign n3278 = ~n18 & ~n3277;
  assign n3279 = ~n3203 & n3220;
  assign n3280 = ~n706 & ~n3279;
  assign n3281 = n3229 & n3280;
  assign n3282 = ~n3278 & n3281;
  assign n3283 = n3232 & ~n3282;
  assign n3284 = ~n3275 & ~n3283;
  assign n3285 = n3211 & n3284;
  assign n3286 = ~n3214 & ~n3285;
  assign n3287 = ~n700 & ~n3270;
  assign n3288 = ~n3189 & ~n3287;
  assign n3289 = ~n3202 & ~n3272;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = n3263 & ~n3290;
  assign n3292 = ~n700 & ~n3278;
  assign n3293 = ~n3189 & ~n3292;
  assign n3294 = ~n3202 & ~n3280;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = n3257 & ~n3295;
  assign n3297 = ~n3291 & ~n3296;
  assign n3298 = ~n3286 & n3297;
  assign n3299 = n923 & ~n3298;
  assign n3300 = ~n3267 & ~n3299;
  assign n3301 = n822 & n3190;
  assign n3302 = Ni40 & n3219;
  assign n3303 = ~n3220 & ~n3302;
  assign n3304 = ~n3301 & ~n3303;
  assign n3305 = n870 & n3304;
  assign n3306 = ~n706 & ~n3305;
  assign n3307 = ~n18 & ~n3306;
  assign n3308 = ~n3203 & n3304;
  assign n3309 = ~n706 & ~n3308;
  assign n3310 = n3229 & n3309;
  assign n3311 = ~n3307 & n3310;
  assign n3312 = n3232 & ~n3311;
  assign n3313 = Ni40 & n3235;
  assign n3314 = ~n3237 & ~n3313;
  assign n3315 = ~n3301 & ~n3314;
  assign n3316 = n870 & n3315;
  assign n3317 = ~n706 & ~n3316;
  assign n3318 = ~n18 & ~n3317;
  assign n3319 = ~n3203 & n3315;
  assign n3320 = ~n706 & ~n3319;
  assign n3321 = n3229 & n3320;
  assign n3322 = ~n3318 & n3321;
  assign n3323 = n3248 & ~n3322;
  assign n3324 = n3211 & ~n3323;
  assign n3325 = ~n3312 & n3324;
  assign n3326 = ~n3213 & ~n3325;
  assign n3327 = ~n700 & ~n3318;
  assign n3328 = ~n3189 & ~n3327;
  assign n3329 = ~n3202 & ~n3320;
  assign n3330 = ~n3328 & ~n3329;
  assign n3331 = n3263 & ~n3330;
  assign n3332 = ~n700 & ~n3307;
  assign n3333 = ~n3189 & ~n3332;
  assign n3334 = ~n3202 & ~n3309;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = n3257 & ~n3335;
  assign n3337 = ~n3331 & ~n3336;
  assign n3338 = n3211 & n3337;
  assign n3339 = ~n3326 & n3338;
  assign n3340 = n736 & ~n3339;
  assign n3341 = n730 & ~n3211;
  assign n3342 = n3213 & ~n3341;
  assign n3343 = n3205 & n3229;
  assign n3344 = ~n3199 & n3343;
  assign n3345 = n691 & n1030;
  assign n3346 = ~n3344 & n3345;
  assign n3347 = ~n3341 & ~n3346;
  assign n3348 = ~n3342 & ~n3347;
  assign n3349 = ~n3340 & ~n3348;
  assign n3350 = n3300 & n3349;
  assign n3351 = ~n3209 & n3350;
  assign n3352 = n1610 & ~n3351;
  assign n3353 = n870 & n3194;
  assign n3354 = ~n706 & ~n3353;
  assign n3355 = ~n18 & ~n3354;
  assign n3356 = ~n700 & ~n3355;
  assign n3357 = ~n3189 & ~n3356;
  assign n3358 = n3194 & ~n3203;
  assign n3359 = ~n706 & ~n3358;
  assign n3360 = ~n3202 & ~n3359;
  assign n3361 = ~n3357 & ~n3360;
  assign n3362 = n3208 & ~n3361;
  assign n3363 = n816 & n3190;
  assign n3364 = ~Ni32 & n3363;
  assign n3365 = n3293 & ~n3364;
  assign n3366 = ~n706 & n3363;
  assign n3367 = n3294 & ~n3366;
  assign n3368 = ~n3365 & ~n3367;
  assign n3369 = n3257 & ~n3368;
  assign n3370 = n3288 & ~n3364;
  assign n3371 = n3289 & ~n3366;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3263 & ~n3372;
  assign n3374 = n3278 & ~n3366;
  assign n3375 = ~n3202 & n3374;
  assign n3376 = n3229 & ~n3375;
  assign n3377 = ~n3367 & n3376;
  assign n3378 = n3232 & ~n3377;
  assign n3379 = ~n3373 & ~n3378;
  assign n3380 = ~n3269 & ~n3366;
  assign n3381 = ~n18 & n3380;
  assign n3382 = ~n3202 & n3381;
  assign n3383 = n3229 & ~n3382;
  assign n3384 = ~n3371 & n3383;
  assign n3385 = n3248 & ~n3384;
  assign n3386 = n3379 & ~n3385;
  assign n3387 = n3211 & n3386;
  assign n3388 = ~n3369 & n3387;
  assign n3389 = n923 & ~n3388;
  assign n3390 = ~n822 & n3190;
  assign n3391 = ~n3222 & ~n3390;
  assign n3392 = n870 & n3391;
  assign n3393 = ~n706 & ~n3392;
  assign n3394 = ~n18 & ~n3393;
  assign n3395 = ~n700 & ~n3394;
  assign n3396 = ~n3189 & ~n3395;
  assign n3397 = ~n3203 & n3391;
  assign n3398 = ~n706 & ~n3397;
  assign n3399 = ~n3202 & ~n3398;
  assign n3400 = ~n3396 & ~n3399;
  assign n3401 = n3257 & ~n3400;
  assign n3402 = n3229 & n3398;
  assign n3403 = ~n3394 & n3402;
  assign n3404 = n3232 & ~n3403;
  assign n3405 = ~n3239 & ~n3390;
  assign n3406 = n870 & n3405;
  assign n3407 = ~n706 & ~n3406;
  assign n3408 = ~n18 & ~n3407;
  assign n3409 = ~n3203 & n3405;
  assign n3410 = ~n706 & ~n3409;
  assign n3411 = n3229 & n3410;
  assign n3412 = ~n3408 & n3411;
  assign n3413 = n3248 & ~n3412;
  assign n3414 = n3211 & ~n3413;
  assign n3415 = ~n3404 & n3414;
  assign n3416 = ~n3214 & ~n3415;
  assign n3417 = ~n700 & ~n3408;
  assign n3418 = ~n3189 & ~n3417;
  assign n3419 = ~n3202 & ~n3410;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = n3263 & ~n3420;
  assign n3422 = ~n3416 & ~n3421;
  assign n3423 = ~n3401 & n3422;
  assign n3424 = n738 & ~n3423;
  assign n3425 = ~n3389 & ~n3424;
  assign n3426 = n3229 & n3359;
  assign n3427 = ~n3355 & n3426;
  assign n3428 = n3345 & ~n3427;
  assign n3429 = ~n3341 & ~n3428;
  assign n3430 = ~n3342 & ~n3429;
  assign n3431 = ~n908 & n3190;
  assign n3432 = ~n3303 & ~n3431;
  assign n3433 = n870 & n3432;
  assign n3434 = ~n706 & ~n3433;
  assign n3435 = ~n18 & ~n3434;
  assign n3436 = ~Ni32 & ~n3435;
  assign n3437 = ~n3203 & n3432;
  assign n3438 = n3436 & ~n3437;
  assign n3439 = n3257 & ~n3438;
  assign n3440 = ~n3189 & n3439;
  assign n3441 = ~n706 & ~n3435;
  assign n3442 = n3229 & n3441;
  assign n3443 = ~n3437 & n3442;
  assign n3444 = n3232 & ~n3443;
  assign n3445 = ~n3314 & ~n3431;
  assign n3446 = n870 & n3445;
  assign n3447 = ~n706 & ~n3446;
  assign n3448 = ~n18 & ~n3447;
  assign n3449 = ~n3203 & n3445;
  assign n3450 = ~n706 & ~n3449;
  assign n3451 = n3229 & n3450;
  assign n3452 = ~n3448 & n3451;
  assign n3453 = n3248 & ~n3452;
  assign n3454 = n3211 & ~n3453;
  assign n3455 = ~n3444 & n3454;
  assign n3456 = ~n3214 & ~n3455;
  assign n3457 = ~n700 & ~n3448;
  assign n3458 = ~n3189 & ~n3457;
  assign n3459 = ~n3202 & ~n3450;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = n3263 & ~n3460;
  assign n3462 = ~n3456 & ~n3461;
  assign n3463 = ~n3440 & n3462;
  assign n3464 = n736 & ~n3463;
  assign n3465 = ~n3430 & ~n3464;
  assign n3466 = n3425 & n3465;
  assign n3467 = ~n3362 & n3466;
  assign n3468 = n1178 & ~n3467;
  assign n3469 = n3309 & n3332;
  assign n3470 = n3257 & ~n3469;
  assign n3471 = n3320 & n3327;
  assign n3472 = n3263 & ~n3471;
  assign n3473 = n3325 & ~n3472;
  assign n3474 = ~n3470 & n3473;
  assign n3475 = n736 & ~n3474;
  assign n3476 = n3245 & n3259;
  assign n3477 = n3263 & ~n3476;
  assign n3478 = n3228 & n3253;
  assign n3479 = n3257 & ~n3478;
  assign n3480 = n3251 & ~n3479;
  assign n3481 = ~n3477 & n3480;
  assign n3482 = n738 & ~n3481;
  assign n3483 = n3347 & ~n3482;
  assign n3484 = n3200 & n3205;
  assign n3485 = n3208 & ~n3484;
  assign n3486 = n3280 & n3292;
  assign n3487 = n3257 & ~n3486;
  assign n3488 = n3272 & n3287;
  assign n3489 = n3263 & ~n3488;
  assign n3490 = ~n3487 & ~n3489;
  assign n3491 = n3285 & n3490;
  assign n3492 = n923 & ~n3491;
  assign n3493 = ~n3485 & ~n3492;
  assign n3494 = n3483 & n3493;
  assign n3495 = ~n3475 & n3494;
  assign n3496 = n1672 & ~n3495;
  assign n3497 = n3450 & n3457;
  assign n3498 = n3263 & ~n3497;
  assign n3499 = ~n3439 & ~n3498;
  assign n3500 = n3455 & n3499;
  assign n3501 = n736 & ~n3500;
  assign n3502 = n3395 & n3398;
  assign n3503 = n3257 & ~n3502;
  assign n3504 = n3410 & n3417;
  assign n3505 = n3263 & ~n3504;
  assign n3506 = n3415 & ~n3505;
  assign n3507 = ~n3503 & n3506;
  assign n3508 = n738 & ~n3507;
  assign n3509 = n3429 & ~n3508;
  assign n3510 = n3356 & n3359;
  assign n3511 = n3208 & ~n3510;
  assign n3512 = n3229 & n3366;
  assign n3513 = ~n3284 & ~n3512;
  assign n3514 = ~n3364 & n3487;
  assign n3515 = ~n3287 & ~n3364;
  assign n3516 = ~n3272 & ~n3366;
  assign n3517 = ~n3515 & ~n3516;
  assign n3518 = n3263 & ~n3517;
  assign n3519 = ~n3514 & ~n3518;
  assign n3520 = n3211 & n3519;
  assign n3521 = ~n3513 & n3520;
  assign n3522 = n923 & ~n3521;
  assign n3523 = ~n3511 & ~n3522;
  assign n3524 = n3509 & n3523;
  assign n3525 = ~n3501 & n3524;
  assign n3526 = n1769 & ~n3525;
  assign n3527 = ~n3496 & ~n3526;
  assign n3528 = ~n3468 & n3527;
  assign n3529 = ~n3352 & n3528;
  assign n3530 = n570 & ~n3529;
  assign n3531 = ~n3187 & ~n3530;
  assign n3532 = ~n3138 & n3531;
  assign n3533 = n694 & ~n3532;
  assign n3534 = Ni12 & n2635;
  assign n3535 = Ni33 & n870;
  assign n3536 = ~n3110 & ~n3535;
  assign n3537 = ~n3196 & ~n3536;
  assign n3538 = ~n706 & ~n3537;
  assign n3539 = n3200 & n3538;
  assign n3540 = ~n604 & n1030;
  assign n3541 = ~n3539 & n3540;
  assign n3542 = n730 & ~n3178;
  assign n3543 = ~n736 & ~n3542;
  assign n3544 = n3304 & ~n3536;
  assign n3545 = ~n706 & ~n3544;
  assign n3546 = n3332 & n3545;
  assign n3547 = ~n604 & n949;
  assign n3548 = ~n3546 & n3547;
  assign n3549 = n3315 & ~n3536;
  assign n3550 = ~n706 & ~n3549;
  assign n3551 = n3327 & n3550;
  assign n3552 = ~n604 & n867;
  assign n3553 = ~n3551 & n3552;
  assign n3554 = ~n3112 & ~n3549;
  assign n3555 = ~n3318 & n3554;
  assign n3556 = n604 & n867;
  assign n3557 = ~n3555 & n3556;
  assign n3558 = ~n3112 & ~n3544;
  assign n3559 = ~n3307 & n3558;
  assign n3560 = n604 & n949;
  assign n3561 = ~n3559 & n3560;
  assign n3562 = ~n3557 & ~n3561;
  assign n3563 = ~n3553 & n3562;
  assign n3564 = n3178 & n3563;
  assign n3565 = ~n3548 & n3564;
  assign n3566 = ~n3543 & ~n3565;
  assign n3567 = n3240 & ~n3536;
  assign n3568 = ~n706 & ~n3567;
  assign n3569 = n3259 & n3568;
  assign n3570 = n3552 & ~n3569;
  assign n3571 = n3223 & ~n3536;
  assign n3572 = ~n706 & ~n3571;
  assign n3573 = n3089 & n3572;
  assign n3574 = ~n3226 & n3573;
  assign n3575 = n3560 & ~n3574;
  assign n3576 = n3089 & n3568;
  assign n3577 = ~n3243 & n3576;
  assign n3578 = n3556 & ~n3577;
  assign n3579 = ~n3575 & ~n3578;
  assign n3580 = n3253 & n3572;
  assign n3581 = n3547 & ~n3580;
  assign n3582 = n3178 & ~n3581;
  assign n3583 = n3579 & n3582;
  assign n3584 = ~n3570 & n3583;
  assign n3585 = n738 & ~n3584;
  assign n3586 = n3237 & ~n3536;
  assign n3587 = ~n3270 & ~n3586;
  assign n3588 = ~Ni32 & n3587;
  assign n3589 = n3552 & ~n3588;
  assign n3590 = n3220 & ~n3536;
  assign n3591 = ~n3278 & ~n3590;
  assign n3592 = ~Ni32 & n3591;
  assign n3593 = n3547 & ~n3592;
  assign n3594 = ~n3589 & ~n3593;
  assign n3595 = ~n3112 & n3591;
  assign n3596 = n3560 & ~n3595;
  assign n3597 = ~n3112 & n3587;
  assign n3598 = n3556 & ~n3597;
  assign n3599 = ~n3596 & ~n3598;
  assign n3600 = n3178 & n3599;
  assign n3601 = n3594 & n3600;
  assign n3602 = n923 & ~n3601;
  assign n3603 = ~n3112 & ~n3537;
  assign n3604 = ~n3199 & n3603;
  assign n3605 = n604 & n1030;
  assign n3606 = ~n3604 & n3605;
  assign n3607 = ~n3602 & ~n3606;
  assign n3608 = ~n3585 & n3607;
  assign n3609 = ~n3566 & n3608;
  assign n3610 = ~n3541 & n3609;
  assign n3611 = n1672 & ~n3610;
  assign n3612 = n3199 & ~n3202;
  assign n3613 = ~n3112 & n3188;
  assign n3614 = ~n3603 & ~n3613;
  assign n3615 = ~n3612 & ~n3614;
  assign n3616 = n3605 & ~n3615;
  assign n3617 = ~n3542 & ~n3616;
  assign n3618 = ~n3202 & ~n3538;
  assign n3619 = ~n3201 & ~n3618;
  assign n3620 = n3540 & ~n3619;
  assign n3621 = ~n706 & ~n3590;
  assign n3622 = ~n3202 & ~n3621;
  assign n3623 = ~n3293 & ~n3622;
  assign n3624 = n3547 & ~n3623;
  assign n3625 = ~n706 & ~n3586;
  assign n3626 = ~n3202 & ~n3625;
  assign n3627 = ~n3288 & ~n3626;
  assign n3628 = n3552 & ~n3627;
  assign n3629 = ~n3624 & ~n3628;
  assign n3630 = n3089 & n3202;
  assign n3631 = n3613 & n3625;
  assign n3632 = ~n3596 & n3631;
  assign n3633 = ~n3630 & ~n3632;
  assign n3634 = ~n3599 & n3633;
  assign n3635 = n3178 & ~n3634;
  assign n3636 = n3629 & n3635;
  assign n3637 = n923 & ~n3636;
  assign n3638 = ~n3620 & ~n3637;
  assign n3639 = ~n3202 & ~n3568;
  assign n3640 = ~n3260 & ~n3639;
  assign n3641 = n3552 & ~n3640;
  assign n3642 = ~n3202 & ~n3572;
  assign n3643 = ~n3254 & ~n3642;
  assign n3644 = n3547 & ~n3643;
  assign n3645 = ~n3579 & ~n3630;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = n3178 & n3646;
  assign n3648 = ~n3641 & n3647;
  assign n3649 = n738 & ~n3648;
  assign n3650 = ~n3202 & n3318;
  assign n3651 = ~n3554 & ~n3613;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = n3556 & ~n3652;
  assign n3654 = ~n3202 & n3307;
  assign n3655 = ~n3558 & ~n3613;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = n3560 & ~n3656;
  assign n3658 = ~n3653 & ~n3657;
  assign n3659 = ~n3202 & ~n3550;
  assign n3660 = ~n3328 & ~n3659;
  assign n3661 = n3552 & ~n3660;
  assign n3662 = ~n3202 & ~n3545;
  assign n3663 = ~n3333 & ~n3662;
  assign n3664 = n3547 & ~n3663;
  assign n3665 = ~n3661 & ~n3664;
  assign n3666 = n3658 & n3665;
  assign n3667 = n3178 & n3666;
  assign n3668 = n736 & ~n3667;
  assign n3669 = ~n3649 & ~n3668;
  assign n3670 = n3638 & n3669;
  assign n3671 = n3617 & n3670;
  assign n3672 = n1610 & ~n3671;
  assign n3673 = ~n738 & ~n3542;
  assign n3674 = n3405 & ~n3536;
  assign n3675 = ~n706 & ~n3674;
  assign n3676 = ~n3202 & ~n3675;
  assign n3677 = ~n3418 & ~n3676;
  assign n3678 = n3552 & ~n3677;
  assign n3679 = n3391 & ~n3536;
  assign n3680 = ~n706 & ~n3679;
  assign n3681 = ~n3202 & ~n3680;
  assign n3682 = ~n3396 & ~n3681;
  assign n3683 = n3547 & ~n3682;
  assign n3684 = n3178 & ~n3683;
  assign n3685 = ~n3678 & n3684;
  assign n3686 = ~n3673 & ~n3685;
  assign n3687 = ~n3366 & ~n3621;
  assign n3688 = n3089 & ~n3374;
  assign n3689 = ~n3687 & n3688;
  assign n3690 = n923 & ~n3689;
  assign n3691 = n3432 & ~n3536;
  assign n3692 = n3089 & n3441;
  assign n3693 = ~n3691 & n3692;
  assign n3694 = n736 & ~n3693;
  assign n3695 = ~n3690 & ~n3694;
  assign n3696 = n3560 & ~n3695;
  assign n3697 = n3089 & n3680;
  assign n3698 = ~n3394 & n3697;
  assign n3699 = n3560 & ~n3698;
  assign n3700 = n3089 & n3675;
  assign n3701 = ~n3408 & n3700;
  assign n3702 = n3556 & ~n3701;
  assign n3703 = ~n3699 & ~n3702;
  assign n3704 = ~n3673 & ~n3703;
  assign n3705 = n3194 & ~n3536;
  assign n3706 = ~n706 & ~n3705;
  assign n3707 = n3089 & n3706;
  assign n3708 = ~n3355 & n3707;
  assign n3709 = n3605 & ~n3708;
  assign n3710 = ~n3366 & ~n3625;
  assign n3711 = n3089 & ~n3381;
  assign n3712 = ~n3710 & n3711;
  assign n3713 = n923 & ~n3712;
  assign n3714 = n3445 & ~n3536;
  assign n3715 = ~n706 & ~n3714;
  assign n3716 = n3089 & n3715;
  assign n3717 = ~n3448 & n3716;
  assign n3718 = n736 & ~n3717;
  assign n3719 = ~n3713 & ~n3718;
  assign n3720 = n3556 & ~n3719;
  assign n3721 = ~n3709 & ~n3720;
  assign n3722 = ~n3704 & n3721;
  assign n3723 = ~n3696 & n3722;
  assign n3724 = ~n3630 & ~n3723;
  assign n3725 = ~n3202 & ~n3706;
  assign n3726 = ~n3357 & ~n3725;
  assign n3727 = n3540 & ~n3726;
  assign n3728 = n3436 & ~n3691;
  assign n3729 = n3547 & ~n3728;
  assign n3730 = ~n3189 & n3729;
  assign n3731 = ~n3202 & ~n3715;
  assign n3732 = ~n3458 & ~n3731;
  assign n3733 = n3552 & ~n3732;
  assign n3734 = n3178 & ~n3733;
  assign n3735 = ~n3730 & n3734;
  assign n3736 = n736 & ~n3735;
  assign n3737 = ~n3727 & ~n3736;
  assign n3738 = ~n3366 & n3622;
  assign n3739 = ~n3365 & ~n3738;
  assign n3740 = n3547 & ~n3739;
  assign n3741 = ~n3366 & n3626;
  assign n3742 = ~n3370 & ~n3741;
  assign n3743 = n3552 & ~n3742;
  assign n3744 = n3178 & ~n3743;
  assign n3745 = ~n3740 & n3744;
  assign n3746 = n923 & ~n3745;
  assign n3747 = n3737 & ~n3746;
  assign n3748 = ~n3724 & n3747;
  assign n3749 = ~n3686 & n3748;
  assign n3750 = n1178 & ~n3749;
  assign n3751 = n3356 & n3706;
  assign n3752 = n3540 & ~n3751;
  assign n3753 = ~n3515 & ~n3710;
  assign n3754 = n3552 & ~n3753;
  assign n3755 = ~n3292 & ~n3364;
  assign n3756 = ~n3687 & ~n3755;
  assign n3757 = n3547 & ~n3756;
  assign n3758 = n3178 & ~n3757;
  assign n3759 = ~n3754 & n3758;
  assign n3760 = n923 & ~n3759;
  assign n3761 = ~n3752 & ~n3760;
  assign n3762 = n3457 & n3715;
  assign n3763 = n3552 & ~n3762;
  assign n3764 = n3178 & ~n3729;
  assign n3765 = ~n3763 & n3764;
  assign n3766 = n736 & ~n3765;
  assign n3767 = n3417 & n3675;
  assign n3768 = n3552 & ~n3767;
  assign n3769 = n3395 & n3680;
  assign n3770 = n3547 & ~n3769;
  assign n3771 = n3178 & ~n3770;
  assign n3772 = ~n3768 & n3771;
  assign n3773 = ~n3673 & ~n3772;
  assign n3774 = ~n3766 & ~n3773;
  assign n3775 = n3723 & n3774;
  assign n3776 = n3761 & n3775;
  assign n3777 = n1769 & ~n3776;
  assign n3778 = ~n3750 & ~n3777;
  assign n3779 = ~n3672 & n3778;
  assign n3780 = ~n3611 & n3779;
  assign n3781 = n3534 & ~n3780;
  assign n3782 = n1625 & ~n3742;
  assign n3783 = n1636 & ~n3677;
  assign n3784 = n1643 & ~n3739;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = n1611 & ~n3682;
  assign n3787 = n3131 & ~n3786;
  assign n3788 = n3785 & n3787;
  assign n3789 = ~n3782 & n3788;
  assign n3790 = n1178 & ~n3789;
  assign n3791 = n1643 & ~n3756;
  assign n3792 = n1625 & ~n3753;
  assign n3793 = n3131 & ~n3792;
  assign n3794 = n1636 & ~n3767;
  assign n3795 = n1611 & ~n3769;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = n3793 & n3796;
  assign n3798 = ~n3791 & n3797;
  assign n3799 = n1769 & ~n3798;
  assign n3800 = n1611 & ~n3643;
  assign n3801 = n1636 & ~n3640;
  assign n3802 = n1643 & ~n3623;
  assign n3803 = n1625 & ~n3627;
  assign n3804 = n3131 & ~n3803;
  assign n3805 = ~n3802 & n3804;
  assign n3806 = ~n3801 & n3805;
  assign n3807 = ~n3800 & n3806;
  assign n3808 = n1610 & ~n3807;
  assign n3809 = ~n3799 & ~n3808;
  assign n3810 = n1636 & ~n3569;
  assign n3811 = n1611 & ~n3580;
  assign n3812 = n1625 & ~n3588;
  assign n3813 = n1643 & ~n3592;
  assign n3814 = n3131 & ~n3813;
  assign n3815 = ~n3812 & n3814;
  assign n3816 = ~n3811 & n3815;
  assign n3817 = ~n3810 & n3816;
  assign n3818 = n1672 & ~n3817;
  assign n3819 = ~Pi17 & ~n3818;
  assign n3820 = n3809 & n3819;
  assign n3821 = ~n3790 & n3820;
  assign n3822 = n1625 & ~n3660;
  assign n3823 = n1643 & ~n3663;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n1610 & ~n3824;
  assign n3826 = n1625 & ~n3551;
  assign n3827 = n1643 & ~n3546;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = n1672 & ~n3828;
  assign n3830 = n1878 & ~n3539;
  assign n3831 = Pi17 & n3131;
  assign n3832 = ~n3830 & n3831;
  assign n3833 = ~n3829 & n3832;
  assign n3834 = n2872 & ~n3619;
  assign n3835 = n1643 & ~n3728;
  assign n3836 = n1625 & ~n3762;
  assign n3837 = n1814 & ~n3751;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n3835 & n3838;
  assign n3840 = n1769 & ~n3839;
  assign n3841 = ~n3834 & ~n3840;
  assign n3842 = n1814 & ~n3726;
  assign n3843 = ~n3189 & n3835;
  assign n3844 = n1625 & ~n3732;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~n3842 & n3845;
  assign n3847 = n1178 & ~n3846;
  assign n3848 = n3841 & ~n3847;
  assign n3849 = n3833 & n3848;
  assign n3850 = ~n3825 & n3849;
  assign n3851 = ~n3821 & ~n3850;
  assign n3852 = Ni13 & Ni12;
  assign n3853 = n3851 & n3852;
  assign n3854 = ~Ni12 & ~n678;
  assign n3855 = n3851 & n3854;
  assign n3856 = ~n1769 & n3189;
  assign n3857 = Pi20 & ~n3220;
  assign n3858 = ~Pi20 & ~n3237;
  assign n3859 = ~n3363 & ~n3858;
  assign n3860 = n870 & n3859;
  assign n3861 = ~n3857 & n3860;
  assign n3862 = ~Ni32 & ~n3861;
  assign n3863 = n1624 & ~n3862;
  assign n3864 = ~Pi20 & n3406;
  assign n3865 = Pi20 & n3392;
  assign n3866 = ~Ni32 & ~n3865;
  assign n3867 = ~n3864 & n3866;
  assign n3868 = n1814 & ~n3867;
  assign n3869 = ~n3863 & ~n3868;
  assign n3870 = ~n3856 & ~n3869;
  assign n3871 = ~Pi20 & ~n3242;
  assign n3872 = Pi20 & ~n3225;
  assign n3873 = ~n700 & ~n3872;
  assign n3874 = ~n3871 & n3873;
  assign n3875 = n1878 & ~n3874;
  assign n3876 = ~Pi16 & n3189;
  assign n3877 = n1624 & ~n3876;
  assign n3878 = ~Pi15 & n3877;
  assign n3879 = ~Pi20 & ~n3269;
  assign n3880 = Pi20 & ~n3277;
  assign n3881 = ~n700 & ~n3880;
  assign n3882 = ~n3879 & n3881;
  assign n3883 = n3878 & ~n3882;
  assign n3884 = ~Pi20 & ~n3240;
  assign n3885 = ~n3188 & ~n3884;
  assign n3886 = Pi20 & ~n3223;
  assign n3887 = n870 & ~n3886;
  assign n3888 = n3885 & n3887;
  assign n3889 = ~Ni32 & ~n3888;
  assign n3890 = n2872 & ~n3889;
  assign n3891 = ~n3883 & ~n3890;
  assign n3892 = ~n3875 & n3891;
  assign n3893 = ~Pi17 & n3892;
  assign n3894 = ~n3870 & n3893;
  assign n3895 = n3131 & n3894;
  assign n3896 = ~Pi20 & n3446;
  assign n3897 = Pi20 & n3433;
  assign n3898 = ~Ni32 & ~n3897;
  assign n3899 = ~n3896 & n3898;
  assign n3900 = n1624 & ~n3899;
  assign n3901 = ~n3856 & n3900;
  assign n3902 = ~Pi20 & ~n3317;
  assign n3903 = Pi20 & ~n3306;
  assign n3904 = ~n700 & ~n3903;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = n3878 & ~n3905;
  assign n3907 = ~n3901 & ~n3906;
  assign n3908 = ~Ni32 & ~n3353;
  assign n3909 = ~n3856 & ~n3908;
  assign n3910 = n1610 & n3197;
  assign n3911 = ~n3189 & n3910;
  assign n3912 = ~n3909 & ~n3911;
  assign n3913 = n1814 & ~n3912;
  assign n3914 = ~Ni32 & ~n3197;
  assign n3915 = n1878 & ~n3914;
  assign n3916 = ~n3913 & ~n3915;
  assign n3917 = n3907 & n3916;
  assign n3918 = n3831 & n3917;
  assign n3919 = n679 & ~n3918;
  assign n3920 = ~n3895 & n3919;
  assign n3921 = ~n3855 & ~n3920;
  assign n3922 = Pi27 & n867;
  assign n3923 = ~n3712 & n3922;
  assign n3924 = Pi27 & n949;
  assign n3925 = ~n3689 & n3924;
  assign n3926 = ~n3923 & ~n3925;
  assign n3927 = ~n3630 & ~n3926;
  assign n3928 = ~Pi27 & n949;
  assign n3929 = ~n3739 & n3928;
  assign n3930 = ~Pi27 & n867;
  assign n3931 = ~n3742 & n3930;
  assign n3932 = ~n3929 & ~n3931;
  assign n3933 = ~n3927 & n3932;
  assign n3934 = n994 & ~n3933;
  assign n3935 = ~n3717 & n3922;
  assign n3936 = ~n3693 & n3924;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~n3630 & ~n3937;
  assign n3939 = ~n3732 & n3930;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = n869 & ~n3940;
  assign n3942 = ~Pi27 & n2205;
  assign n3943 = ~n3726 & n3942;
  assign n3944 = Pi27 & n1528;
  assign n3945 = Pi27 & n2205;
  assign n3946 = ~n3630 & n3945;
  assign n3947 = ~n3944 & ~n3946;
  assign n3948 = ~n3708 & ~n3947;
  assign n3949 = ~Pi27 & n1528;
  assign n3950 = ~n3751 & n3949;
  assign n3951 = ~n3948 & ~n3950;
  assign n3952 = ~n3943 & n3951;
  assign n3953 = n3143 & n3952;
  assign n3954 = n736 & ~n3876;
  assign n3955 = n3928 & n3954;
  assign n3956 = ~n3728 & n3955;
  assign n3957 = Pi15 & ~n3956;
  assign n3958 = n3953 & n3957;
  assign n3959 = ~n3941 & n3958;
  assign n3960 = ~n3762 & n3930;
  assign n3961 = n3937 & ~n3960;
  assign n3962 = n1035 & ~n3961;
  assign n3963 = ~n3769 & n3928;
  assign n3964 = ~n3701 & n3922;
  assign n3965 = ~n3698 & n3924;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3767 & n3930;
  assign n3968 = n3966 & ~n3967;
  assign n3969 = ~n3963 & n3968;
  assign n3970 = n955 & ~n3969;
  assign n3971 = ~n3756 & n3928;
  assign n3972 = ~n3753 & n3930;
  assign n3973 = n3926 & ~n3972;
  assign n3974 = ~n3971 & n3973;
  assign n3975 = n924 & ~n3974;
  assign n3976 = ~n3970 & ~n3975;
  assign n3977 = ~n3630 & ~n3966;
  assign n3978 = ~n3677 & n3930;
  assign n3979 = ~n3682 & n3928;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = ~n3977 & n3980;
  assign n3982 = n903 & ~n3981;
  assign n3983 = n3976 & ~n3982;
  assign n3984 = ~n3962 & n3983;
  assign n3985 = n3959 & n3984;
  assign n3986 = ~n3934 & n3985;
  assign n3987 = ~n3640 & n3930;
  assign n3988 = ~n3577 & n3922;
  assign n3989 = ~n3574 & n3924;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3630 & ~n3990;
  assign n3992 = ~n3643 & n3928;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~n3987 & n3993;
  assign n3995 = n903 & ~n3994;
  assign n3996 = ~n3559 & n3924;
  assign n3997 = ~n3546 & n3928;
  assign n3998 = ~n3551 & n3930;
  assign n3999 = ~n3555 & n3922;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = ~n3997 & n4000;
  assign n4002 = ~n3996 & n4001;
  assign n4003 = n1035 & ~n4002;
  assign n4004 = ~n3995 & ~n4003;
  assign n4005 = ~n3597 & n3922;
  assign n4006 = ~n3595 & n3924;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = ~n3588 & n3930;
  assign n4009 = ~n3592 & n3928;
  assign n4010 = ~n4008 & ~n4009;
  assign n4011 = n4007 & n4010;
  assign n4012 = n924 & ~n4011;
  assign n4013 = ~n3630 & ~n4007;
  assign n4014 = ~n3627 & n3930;
  assign n4015 = ~n3623 & n3928;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n4013 & n4016;
  assign n4018 = n994 & ~n4017;
  assign n4019 = ~n3604 & n3944;
  assign n4020 = ~n3539 & n3949;
  assign n4021 = ~Pi15 & ~n4020;
  assign n4022 = ~n3619 & n3942;
  assign n4023 = ~n3615 & n3945;
  assign n4024 = n3143 & ~n4023;
  assign n4025 = ~n4022 & n4024;
  assign n4026 = n4021 & n4025;
  assign n4027 = ~n4019 & n4026;
  assign n4028 = ~n4018 & n4027;
  assign n4029 = ~n4012 & n4028;
  assign n4030 = ~n3569 & n3930;
  assign n4031 = ~n3580 & n3928;
  assign n4032 = n3990 & ~n4031;
  assign n4033 = ~n4030 & n4032;
  assign n4034 = n955 & ~n4033;
  assign n4035 = ~n3663 & n3928;
  assign n4036 = ~n3656 & n3924;
  assign n4037 = ~n3652 & n3922;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~n3660 & n3930;
  assign n4040 = n4038 & ~n4039;
  assign n4041 = ~n4035 & n4040;
  assign n4042 = n869 & ~n4041;
  assign n4043 = ~n4034 & ~n4042;
  assign n4044 = n4029 & n4043;
  assign n4045 = n4004 & n4044;
  assign n4046 = Ni12 & n678;
  assign n4047 = ~n4045 & n4046;
  assign n4048 = ~n3986 & n4047;
  assign n4049 = n3921 & ~n4048;
  assign n4050 = ~n3853 & n4049;
  assign n4051 = ~n3781 & n4050;
  assign n4052 = ~Ni11 & ~n4051;
  assign n4053 = n677 & n1030;
  assign n4054 = ~n3604 & n4053;
  assign n4055 = n730 & ~n3105;
  assign n4056 = ~n923 & ~n4055;
  assign n4057 = n677 & n949;
  assign n4058 = ~n3595 & n4057;
  assign n4059 = n677 & n867;
  assign n4060 = ~n3597 & n4059;
  assign n4061 = ~n4058 & ~n4060;
  assign n4062 = ~n677 & n867;
  assign n4063 = ~n3588 & n4062;
  assign n4064 = n4061 & ~n4063;
  assign n4065 = ~n677 & n949;
  assign n4066 = ~n3592 & n4065;
  assign n4067 = n3105 & ~n4066;
  assign n4068 = n4064 & n4067;
  assign n4069 = ~n4056 & ~n4068;
  assign n4070 = ~n4054 & ~n4069;
  assign n4071 = ~n3555 & n4059;
  assign n4072 = ~n3559 & n4057;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = ~n3551 & n4062;
  assign n4075 = ~n3546 & n4065;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = n3105 & n4076;
  assign n4078 = n4073 & n4077;
  assign n4079 = n736 & ~n4078;
  assign n4080 = ~n3577 & n4059;
  assign n4081 = ~n3574 & n4057;
  assign n4082 = n3105 & ~n4081;
  assign n4083 = ~n4080 & n4082;
  assign n4084 = ~n3580 & n4065;
  assign n4085 = ~n3569 & n4062;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = n4083 & n4086;
  assign n4088 = n738 & ~n4087;
  assign n4089 = ~n677 & n1030;
  assign n4090 = ~n3539 & n4089;
  assign n4091 = ~n4088 & ~n4090;
  assign n4092 = ~n4079 & n4091;
  assign n4093 = n4070 & n4092;
  assign n4094 = n1672 & ~n4093;
  assign n4095 = ~n3693 & n4057;
  assign n4096 = ~n3717 & n4059;
  assign n4097 = n3105 & ~n4096;
  assign n4098 = ~n4095 & n4097;
  assign n4099 = n3105 & n3630;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = ~n3728 & n4065;
  assign n4102 = ~n3189 & n4101;
  assign n4103 = ~n3732 & n4062;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4100 & n4104;
  assign n4106 = n736 & ~n4105;
  assign n4107 = ~n3742 & n4062;
  assign n4108 = ~n3689 & n4057;
  assign n4109 = ~n3712 & n4059;
  assign n4110 = n3105 & ~n4109;
  assign n4111 = ~n4108 & n4110;
  assign n4112 = ~n4099 & ~n4111;
  assign n4113 = ~n3739 & n4065;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = ~n4107 & n4114;
  assign n4116 = n923 & ~n4115;
  assign n4117 = ~n3682 & n4065;
  assign n4118 = ~n3677 & n4062;
  assign n4119 = ~n3698 & n4057;
  assign n4120 = n3105 & ~n4119;
  assign n4121 = ~n4099 & ~n4120;
  assign n4122 = ~n4118 & ~n4121;
  assign n4123 = ~n4117 & n4122;
  assign n4124 = n738 & ~n4123;
  assign n4125 = ~n3708 & n4053;
  assign n4126 = n738 & n4059;
  assign n4127 = ~n3701 & n4126;
  assign n4128 = ~n4125 & ~n4127;
  assign n4129 = ~n3630 & ~n4128;
  assign n4130 = ~n4124 & ~n4129;
  assign n4131 = ~n4116 & n4130;
  assign n4132 = ~n3726 & n4089;
  assign n4133 = ~n4055 & ~n4132;
  assign n4134 = n4131 & n4133;
  assign n4135 = ~n4106 & n4134;
  assign n4136 = n1178 & ~n4135;
  assign n4137 = ~n3762 & n4062;
  assign n4138 = ~n4101 & ~n4137;
  assign n4139 = n4098 & n4138;
  assign n4140 = n736 & ~n4139;
  assign n4141 = ~n3756 & n4065;
  assign n4142 = ~n3753 & n4062;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = n4111 & n4143;
  assign n4145 = n923 & ~n4144;
  assign n4146 = ~n3769 & n4065;
  assign n4147 = ~n3767 & n4062;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = n4120 & n4148;
  assign n4150 = n738 & ~n4149;
  assign n4151 = ~n4145 & ~n4150;
  assign n4152 = ~n4140 & n4151;
  assign n4153 = ~n3751 & n4089;
  assign n4154 = n4128 & ~n4153;
  assign n4155 = n4152 & n4154;
  assign n4156 = ~n4055 & n4155;
  assign n4157 = n1769 & ~n4156;
  assign n4158 = ~n3660 & n4062;
  assign n4159 = ~n3663 & n4065;
  assign n4160 = ~n3652 & n4059;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = ~n3656 & n4057;
  assign n4163 = n3105 & ~n4162;
  assign n4164 = n4161 & n4163;
  assign n4165 = ~n4158 & n4164;
  assign n4166 = n736 & ~n4165;
  assign n4167 = ~n4083 & ~n4099;
  assign n4168 = ~n3643 & n4065;
  assign n4169 = ~n3640 & n4062;
  assign n4170 = ~n4168 & ~n4169;
  assign n4171 = ~n4167 & n4170;
  assign n4172 = n738 & ~n4171;
  assign n4173 = ~n3615 & n4053;
  assign n4174 = ~n3619 & n4089;
  assign n4175 = ~n4173 & ~n4174;
  assign n4176 = ~n3631 & n4060;
  assign n4177 = ~n4058 & ~n4176;
  assign n4178 = ~n3630 & ~n4177;
  assign n4179 = ~n3627 & n4062;
  assign n4180 = ~n3623 & n4065;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = n3105 & n4181;
  assign n4183 = ~n4178 & n4182;
  assign n4184 = ~n4056 & ~n4183;
  assign n4185 = n4175 & ~n4184;
  assign n4186 = ~n4172 & n4185;
  assign n4187 = ~n4166 & n4186;
  assign n4188 = n1610 & ~n4187;
  assign n4189 = ~n4157 & ~n4188;
  assign n4190 = ~n4136 & n4189;
  assign n4191 = ~n4094 & n4190;
  assign n4192 = n680 & ~n4191;
  assign n4193 = Ni11 & ~n679;
  assign n4194 = n3851 & n4193;
  assign n4195 = ~n4192 & ~n4194;
  assign n4196 = Ni10 & n4195;
  assign n4197 = ~n4052 & n4196;
  assign n4198 = n2388 & ~n3874;
  assign n4199 = n2462 & ~n3889;
  assign n4200 = n1031 & ~n3914;
  assign n4201 = ~n3876 & n4200;
  assign n4202 = n3131 & ~n4201;
  assign n4203 = ~Pi15 & n4202;
  assign n4204 = ~n4199 & n4203;
  assign n4205 = ~n4198 & n4204;
  assign n4206 = n865 & ~n3876;
  assign n4207 = n923 & ~n3882;
  assign n4208 = n736 & ~n3905;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = n4206 & ~n4209;
  assign n4211 = n4205 & ~n4210;
  assign n4212 = n923 & ~n3862;
  assign n4213 = n738 & ~n3867;
  assign n4214 = n730 & ~n3908;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = n736 & ~n3899;
  assign n4217 = n4215 & ~n4216;
  assign n4218 = ~n4212 & n4217;
  assign n4219 = n4206 & ~n4218;
  assign n4220 = Pi15 & n3131;
  assign n4221 = ~n4219 & n4220;
  assign n4222 = ~n4211 & ~n4221;
  assign n4223 = ~Pi25 & ~n3134;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~Ni10 & n4224;
  assign n4226 = ~n3852 & ~n4193;
  assign n4227 = ~Ni10 & n4226;
  assign n4228 = ~n4225 & ~n4227;
  assign n4229 = n3854 & ~n4224;
  assign n4230 = ~Pi25 & n867;
  assign n4231 = ~n3372 & n4230;
  assign n4232 = ~Pi25 & n949;
  assign n4233 = ~n3368 & n4232;
  assign n4234 = n865 & ~n3862;
  assign n4235 = ~n3189 & n4234;
  assign n4236 = ~n4233 & ~n4235;
  assign n4237 = ~n4231 & n4236;
  assign n4238 = n994 & ~n4237;
  assign n4239 = Pi15 & ~n4238;
  assign n4240 = n869 & n4230;
  assign n4241 = ~n3460 & n4240;
  assign n4242 = ~n3486 & n4232;
  assign n4243 = ~n3364 & n4242;
  assign n4244 = ~n3517 & n4230;
  assign n4245 = ~n4234 & ~n4244;
  assign n4246 = ~n4243 & n4245;
  assign n4247 = n924 & ~n4246;
  assign n4248 = ~n4241 & ~n4247;
  assign n4249 = n955 & n4232;
  assign n4250 = ~n3502 & n4249;
  assign n4251 = n4248 & ~n4250;
  assign n4252 = n4239 & n4251;
  assign n4253 = ~n3438 & n4232;
  assign n4254 = ~n3876 & n4253;
  assign n4255 = ~n3899 & n4206;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = n736 & ~n4256;
  assign n4258 = n1035 & n4230;
  assign n4259 = ~n3497 & n4258;
  assign n4260 = ~n4257 & ~n4259;
  assign n4261 = ~n3400 & n4232;
  assign n4262 = ~n3420 & n4230;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = n903 & ~n4263;
  assign n4265 = n955 & n4230;
  assign n4266 = ~n3504 & n4265;
  assign n4267 = n4206 & ~n4215;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n1814 & ~n3510;
  assign n4270 = n2159 & n4269;
  assign n4271 = n2205 & ~n3361;
  assign n4272 = n3131 & ~n4271;
  assign n4273 = ~n4270 & n4272;
  assign n4274 = n4268 & n4273;
  assign n4275 = ~n4264 & n4274;
  assign n4276 = n4260 & n4275;
  assign n4277 = n4252 & n4276;
  assign n4278 = n1035 & ~n3469;
  assign n4279 = n955 & ~n3478;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = n869 & ~n3335;
  assign n4282 = n994 & ~n3295;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = n4280 & n4283;
  assign n4285 = n4232 & ~n4284;
  assign n4286 = ~n3262 & n4230;
  assign n4287 = ~n3256 & n4232;
  assign n4288 = ~n4286 & ~n4287;
  assign n4289 = n903 & ~n4288;
  assign n4290 = ~n3471 & n4258;
  assign n4291 = ~n3476 & n4265;
  assign n4292 = n865 & ~n3882;
  assign n4293 = ~n4242 & ~n4292;
  assign n4294 = n924 & ~n4293;
  assign n4295 = n924 & n4230;
  assign n4296 = ~n3488 & n4295;
  assign n4297 = n2205 & ~n3207;
  assign n4298 = n1814 & ~n3484;
  assign n4299 = n2159 & n4298;
  assign n4300 = ~n4297 & ~n4299;
  assign n4301 = ~n4296 & n4300;
  assign n4302 = ~n4294 & n4301;
  assign n4303 = ~n4291 & n4302;
  assign n4304 = ~n4290 & n4303;
  assign n4305 = ~n4289 & n4304;
  assign n4306 = ~n3330 & n4240;
  assign n4307 = n4206 & n4208;
  assign n4308 = n994 & n4230;
  assign n4309 = ~n3290 & n4308;
  assign n4310 = n994 & n4292;
  assign n4311 = ~n3189 & n4310;
  assign n4312 = ~n4309 & ~n4311;
  assign n4313 = ~n4307 & n4312;
  assign n4314 = ~n4306 & n4313;
  assign n4315 = n4205 & n4314;
  assign n4316 = n4305 & n4315;
  assign n4317 = ~n4285 & n4316;
  assign n4318 = n679 & ~n4317;
  assign n4319 = ~n4277 & n4318;
  assign n4320 = ~n4229 & ~n4319;
  assign n4321 = ~n604 & n865;
  assign n4322 = ~n4218 & n4321;
  assign n4323 = ~n3189 & n4322;
  assign n4324 = n604 & n868;
  assign n4325 = ~n3112 & ~n3446;
  assign n4326 = n4324 & ~n4325;
  assign n4327 = n2282 & ~n3180;
  assign n4328 = n3178 & ~n4327;
  assign n4329 = n604 & n950;
  assign n4330 = ~n3112 & ~n3433;
  assign n4331 = n4329 & ~n4330;
  assign n4332 = n4328 & ~n4331;
  assign n4333 = ~n4326 & n4332;
  assign n4334 = n736 & ~n4333;
  assign n4335 = n3089 & ~n3380;
  assign n4336 = n4324 & ~n4335;
  assign n4337 = ~n3112 & ~n3276;
  assign n4338 = n4329 & ~n4337;
  assign n4339 = n4328 & ~n4338;
  assign n4340 = ~n3112 & n3363;
  assign n4341 = n4328 & n4340;
  assign n4342 = ~n4339 & ~n4341;
  assign n4343 = ~n4336 & ~n4342;
  assign n4344 = n923 & ~n4343;
  assign n4345 = ~n3112 & ~n3406;
  assign n4346 = n4324 & ~n4345;
  assign n4347 = n4328 & ~n4346;
  assign n4348 = n738 & ~n4347;
  assign n4349 = ~n3112 & ~n3392;
  assign n4350 = n738 & n4329;
  assign n4351 = ~n4349 & n4350;
  assign n4352 = ~n4348 & ~n4351;
  assign n4353 = ~n4344 & n4352;
  assign n4354 = ~n4334 & n4353;
  assign n4355 = n3630 & n4328;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n730 & ~n4328;
  assign n4358 = ~n3112 & ~n3353;
  assign n4359 = n604 & n1031;
  assign n4360 = ~n4358 & n4359;
  assign n4361 = ~n3630 & n4360;
  assign n4362 = ~n4357 & ~n4361;
  assign n4363 = ~n4356 & n4362;
  assign n4364 = ~n4323 & n4363;
  assign n4365 = n1178 & ~n4364;
  assign n4366 = ~n3112 & ~n3268;
  assign n4367 = n4324 & ~n4366;
  assign n4368 = n4339 & ~n4367;
  assign n4369 = ~n4355 & ~n4368;
  assign n4370 = ~n3882 & n4321;
  assign n4371 = ~n3189 & n4370;
  assign n4372 = ~n4369 & ~n4371;
  assign n4373 = n923 & ~n4372;
  assign n4374 = ~n604 & n4200;
  assign n4375 = ~n3189 & n4374;
  assign n4376 = ~n4357 & ~n4375;
  assign n4377 = ~n4373 & n4376;
  assign n4378 = ~n3112 & ~n3305;
  assign n4379 = n4329 & ~n4378;
  assign n4380 = ~n3112 & ~n3316;
  assign n4381 = n4324 & ~n4380;
  assign n4382 = n4328 & ~n4381;
  assign n4383 = ~n4379 & n4382;
  assign n4384 = ~n4355 & ~n4383;
  assign n4385 = ~n3905 & n4321;
  assign n4386 = ~n3189 & n4385;
  assign n4387 = ~n4384 & ~n4386;
  assign n4388 = n736 & ~n4387;
  assign n4389 = ~n3112 & ~n3241;
  assign n4390 = n4324 & ~n4389;
  assign n4391 = n4328 & ~n4390;
  assign n4392 = ~n4355 & ~n4391;
  assign n4393 = ~n3889 & n4321;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = n738 & ~n4394;
  assign n4396 = ~n3112 & ~n3197;
  assign n4397 = n4359 & ~n4396;
  assign n4398 = ~n3112 & ~n3224;
  assign n4399 = n4350 & ~n4398;
  assign n4400 = ~n4397 & ~n4399;
  assign n4401 = ~n3630 & ~n4400;
  assign n4402 = ~n4395 & ~n4401;
  assign n4403 = ~n4388 & n4402;
  assign n4404 = n4377 & n4403;
  assign n4405 = n1610 & ~n4404;
  assign n4406 = ~n4365 & ~n4405;
  assign n4407 = n4383 & ~n4385;
  assign n4408 = n736 & ~n4407;
  assign n4409 = ~n3874 & n4321;
  assign n4410 = n4391 & ~n4409;
  assign n4411 = n738 & ~n4410;
  assign n4412 = n4400 & ~n4411;
  assign n4413 = n4368 & ~n4370;
  assign n4414 = n923 & ~n4413;
  assign n4415 = ~n4374 & ~n4414;
  assign n4416 = n4412 & n4415;
  assign n4417 = ~n4408 & n4416;
  assign n4418 = n1672 & ~n4417;
  assign n4419 = Pi16 & n4357;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = ~n4322 & n4354;
  assign n4422 = ~n4360 & n4421;
  assign n4423 = n1769 & ~n4422;
  assign n4424 = ~Ni14 & ~n4423;
  assign n4425 = n4420 & n4424;
  assign n4426 = n4406 & n4425;
  assign n4427 = ~Ni13 & Ni12;
  assign n4428 = ~Pi27 & n4200;
  assign n4429 = ~Pi27 & n865;
  assign n4430 = ~n4209 & n4429;
  assign n4431 = ~n4428 & ~n4430;
  assign n4432 = ~n3189 & ~n4431;
  assign n4433 = Pi25 & n3143;
  assign n4434 = ~n3146 & ~n4433;
  assign n4435 = Pi27 & n950;
  assign n4436 = ~n4337 & n4435;
  assign n4437 = Pi27 & n868;
  assign n4438 = ~n4366 & n4437;
  assign n4439 = ~n4436 & ~n4438;
  assign n4440 = ~n4434 & n4439;
  assign n4441 = n923 & ~n4440;
  assign n4442 = ~n4380 & n4437;
  assign n4443 = ~n4378 & n4435;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4434 & n4444;
  assign n4446 = n736 & ~n4445;
  assign n4447 = ~n4398 & n4435;
  assign n4448 = ~n4389 & n4437;
  assign n4449 = ~n4434 & ~n4448;
  assign n4450 = ~n4447 & n4449;
  assign n4451 = n738 & ~n4450;
  assign n4452 = ~n4446 & ~n4451;
  assign n4453 = ~n4441 & n4452;
  assign n4454 = n3630 & ~n4434;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = n738 & n4429;
  assign n4457 = ~n3889 & n4456;
  assign n4458 = n730 & n4434;
  assign n4459 = Pi27 & n1031;
  assign n4460 = ~n4396 & n4459;
  assign n4461 = ~n4458 & ~n4460;
  assign n4462 = n3630 & ~n4458;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = ~n4457 & ~n4463;
  assign n4465 = ~n4455 & n4464;
  assign n4466 = ~n4432 & n4465;
  assign n4467 = n1610 & ~n4466;
  assign n4468 = ~n4218 & n4429;
  assign n4469 = ~n4349 & n4435;
  assign n4470 = ~n4345 & n4437;
  assign n4471 = ~n4434 & ~n4470;
  assign n4472 = ~n4469 & n4471;
  assign n4473 = n738 & ~n4472;
  assign n4474 = ~n4330 & n4435;
  assign n4475 = ~n4325 & n4437;
  assign n4476 = ~n4434 & ~n4475;
  assign n4477 = ~n4474 & n4476;
  assign n4478 = n736 & ~n4477;
  assign n4479 = ~n4335 & n4437;
  assign n4480 = ~n4340 & n4436;
  assign n4481 = ~n4434 & ~n4480;
  assign n4482 = ~n4479 & n4481;
  assign n4483 = n923 & ~n4482;
  assign n4484 = ~n4478 & ~n4483;
  assign n4485 = ~n4473 & n4484;
  assign n4486 = ~n4358 & n4459;
  assign n4487 = ~n4458 & ~n4486;
  assign n4488 = n4485 & n4487;
  assign n4489 = ~n4468 & n4488;
  assign n4490 = n1769 & ~n4489;
  assign n4491 = ~n3874 & n4456;
  assign n4492 = n4461 & ~n4491;
  assign n4493 = n4453 & n4492;
  assign n4494 = n4431 & n4493;
  assign n4495 = n1672 & ~n4494;
  assign n4496 = Ni14 & ~n4495;
  assign n4497 = ~n4490 & n4496;
  assign n4498 = n3613 & ~n4458;
  assign n4499 = ~n4487 & ~n4498;
  assign n4500 = ~n4454 & ~n4485;
  assign n4501 = ~n3189 & n4468;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = ~n4499 & n4502;
  assign n4504 = n1178 & ~n4503;
  assign n4505 = n4497 & ~n4504;
  assign n4506 = ~n4467 & n4505;
  assign n4507 = n4427 & ~n4506;
  assign n4508 = ~n4426 & n4507;
  assign n4509 = n4320 & ~n4508;
  assign n4510 = ~Ni11 & ~n4509;
  assign n4511 = ~Pi25 & n3117;
  assign n4512 = n3105 & ~n4511;
  assign n4513 = n730 & ~n4512;
  assign n4514 = ~n677 & n865;
  assign n4515 = ~n4209 & n4514;
  assign n4516 = ~n677 & n1031;
  assign n4517 = ~n3914 & n4516;
  assign n4518 = ~n4515 & ~n4517;
  assign n4519 = ~n3189 & ~n4518;
  assign n4520 = n677 & n868;
  assign n4521 = ~n4366 & n4520;
  assign n4522 = n677 & n950;
  assign n4523 = ~n4337 & n4522;
  assign n4524 = n4512 & ~n4523;
  assign n4525 = ~n4521 & n4524;
  assign n4526 = n923 & ~n4525;
  assign n4527 = ~n4378 & n4522;
  assign n4528 = ~n4380 & n4520;
  assign n4529 = n4512 & ~n4528;
  assign n4530 = ~n4527 & n4529;
  assign n4531 = n736 & ~n4530;
  assign n4532 = ~n4526 & ~n4531;
  assign n4533 = n3630 & n4512;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = n677 & n1031;
  assign n4536 = ~n4396 & n4535;
  assign n4537 = ~n4389 & n4520;
  assign n4538 = ~n4398 & n4522;
  assign n4539 = n4512 & ~n4538;
  assign n4540 = ~n4537 & n4539;
  assign n4541 = n738 & ~n4540;
  assign n4542 = ~n4536 & ~n4541;
  assign n4543 = ~n3630 & ~n4542;
  assign n4544 = n738 & ~n4512;
  assign n4545 = n738 & n4514;
  assign n4546 = ~n3889 & n4545;
  assign n4547 = ~n4544 & ~n4546;
  assign n4548 = n1610 & n4547;
  assign n4549 = ~n4543 & n4548;
  assign n4550 = ~n4534 & n4549;
  assign n4551 = ~n4519 & n4550;
  assign n4552 = ~Pi16 & n3630;
  assign n4553 = n4512 & n4552;
  assign n4554 = ~n4325 & n4520;
  assign n4555 = ~n4330 & n4522;
  assign n4556 = n4512 & ~n4555;
  assign n4557 = ~n4554 & n4556;
  assign n4558 = n736 & ~n4557;
  assign n4559 = ~n4349 & n4522;
  assign n4560 = ~n4345 & n4520;
  assign n4561 = n4512 & ~n4560;
  assign n4562 = ~n4559 & n4561;
  assign n4563 = n738 & ~n4562;
  assign n4564 = ~n4335 & n4520;
  assign n4565 = n4340 & n4512;
  assign n4566 = ~n4524 & ~n4565;
  assign n4567 = ~n4564 & ~n4566;
  assign n4568 = n923 & ~n4567;
  assign n4569 = ~n4563 & ~n4568;
  assign n4570 = ~n4558 & n4569;
  assign n4571 = ~n4553 & ~n4570;
  assign n4572 = ~n677 & n4219;
  assign n4573 = n4535 & ~n4552;
  assign n4574 = ~n4358 & n4573;
  assign n4575 = Pi15 & ~n4574;
  assign n4576 = ~n4572 & n4575;
  assign n4577 = ~n4571 & n4576;
  assign n4578 = ~n4551 & ~n4577;
  assign n4579 = ~n4513 & ~n4578;
  assign n4580 = n1672 & ~n4513;
  assign n4581 = n4542 & n4580;
  assign n4582 = ~n3874 & n4545;
  assign n4583 = n4532 & ~n4582;
  assign n4584 = n4518 & n4583;
  assign n4585 = n4581 & n4584;
  assign n4586 = n680 & ~n4585;
  assign n4587 = ~n4579 & n4586;
  assign n4588 = ~n4510 & ~n4587;
  assign n4589 = ~n4228 & n4588;
  assign n4590 = n579 & ~n4589;
  assign n4591 = ~n4197 & n4590;
  assign n4592 = ~n686 & ~n693;
  assign n4593 = ~n3135 & n3854;
  assign n4594 = n1643 & ~n3438;
  assign n4595 = n3131 & ~n4594;
  assign n4596 = ~n3101 & n3189;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = n1814 & ~n3361;
  assign n4599 = n1625 & ~n3460;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = ~n4597 & n4600;
  assign n4602 = n1178 & ~n4601;
  assign n4603 = n1643 & ~n3335;
  assign n4604 = n1625 & ~n3330;
  assign n4605 = n3131 & ~n4604;
  assign n4606 = ~n4603 & n4605;
  assign n4607 = n1610 & ~n4606;
  assign n4608 = ~n4602 & ~n4607;
  assign n4609 = n1625 & ~n3471;
  assign n4610 = n1643 & ~n3469;
  assign n4611 = ~n4298 & ~n4610;
  assign n4612 = n3131 & n4611;
  assign n4613 = ~n4609 & n4612;
  assign n4614 = n1672 & ~n4613;
  assign n4615 = n1625 & ~n3497;
  assign n4616 = ~n4269 & ~n4615;
  assign n4617 = n4595 & n4616;
  assign n4618 = n1769 & ~n4617;
  assign n4619 = n2872 & ~n3207;
  assign n4620 = Pi17 & ~n4619;
  assign n4621 = ~n4618 & n4620;
  assign n4622 = ~n4614 & n4621;
  assign n4623 = n4608 & n4622;
  assign n4624 = n1636 & ~n3420;
  assign n4625 = n1625 & ~n3372;
  assign n4626 = n3131 & ~n4625;
  assign n4627 = n1611 & ~n3400;
  assign n4628 = n1643 & ~n3368;
  assign n4629 = ~n4627 & ~n4628;
  assign n4630 = n4626 & n4629;
  assign n4631 = ~n4624 & n4630;
  assign n4632 = n1178 & ~n4631;
  assign n4633 = n1643 & ~n3295;
  assign n4634 = n1625 & ~n3290;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = n1611 & ~n3256;
  assign n4637 = n1636 & ~n3262;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = n4635 & n4638;
  assign n4640 = n3131 & n4639;
  assign n4641 = n1610 & ~n4640;
  assign n4642 = n1611 & ~n3502;
  assign n4643 = n1643 & ~n3486;
  assign n4644 = n3131 & ~n4643;
  assign n4645 = ~n3101 & n3364;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = n1625 & ~n3517;
  assign n4648 = n1636 & ~n3504;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4646 & n4649;
  assign n4651 = ~n4642 & n4650;
  assign n4652 = n1769 & ~n4651;
  assign n4653 = ~n4641 & ~n4652;
  assign n4654 = n1636 & ~n3476;
  assign n4655 = n1611 & ~n3478;
  assign n4656 = n1625 & ~n3488;
  assign n4657 = n4644 & ~n4656;
  assign n4658 = ~n4655 & n4657;
  assign n4659 = ~n4654 & n4658;
  assign n4660 = n1672 & ~n4659;
  assign n4661 = ~Pi17 & ~n4660;
  assign n4662 = n4653 & n4661;
  assign n4663 = ~n4632 & n4662;
  assign n4664 = n679 & ~n4663;
  assign n4665 = ~n4623 & n4664;
  assign n4666 = ~n4593 & ~n4665;
  assign n4667 = ~Ni11 & ~n4666;
  assign n4668 = ~n3135 & ~n4226;
  assign n4669 = n2635 & ~n3182;
  assign n4670 = n678 & ~n3146;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = Ni12 & ~n4671;
  assign n4673 = ~n4668 & ~n4672;
  assign n4674 = Ni11 & n3135;
  assign n4675 = ~n680 & ~n4674;
  assign n4676 = ~n4673 & n4675;
  assign n4677 = n679 & n3119;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = ~n4667 & n4678;
  assign n4680 = n4592 & ~n4679;
  assign n4681 = Ni8 & n686;
  assign n4682 = Ni10 & n4681;
  assign n4683 = Pi24 & n1528;
  assign n4684 = Pi24 & n2205;
  assign n4685 = ~n3213 & n4684;
  assign n4686 = ~n4683 & ~n4685;
  assign n4687 = ~n3427 & ~n4686;
  assign n4688 = ~Pi24 & ~n4273;
  assign n4689 = n3126 & ~n4688;
  assign n4690 = ~n4687 & n4689;
  assign n4691 = ~Pi24 & n867;
  assign n4692 = ~n3420 & n4691;
  assign n4693 = Pi24 & n867;
  assign n4694 = ~n3412 & n4693;
  assign n4695 = Pi24 & n949;
  assign n4696 = ~n3403 & n4695;
  assign n4697 = ~n4694 & ~n4696;
  assign n4698 = ~n3213 & ~n4697;
  assign n4699 = ~Pi24 & n949;
  assign n4700 = ~n3400 & n4699;
  assign n4701 = ~n4698 & ~n4700;
  assign n4702 = ~n4692 & n4701;
  assign n4703 = n903 & ~n4702;
  assign n4704 = n4690 & ~n4703;
  assign n4705 = ~n3438 & n4699;
  assign n4706 = ~n3452 & n4693;
  assign n4707 = ~n3443 & n4695;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n3497 & n4691;
  assign n4710 = n4708 & ~n4709;
  assign n4711 = ~n4705 & n4710;
  assign n4712 = n1035 & ~n4711;
  assign n4713 = ~n3377 & n4695;
  assign n4714 = ~n3384 & n4693;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = ~n3372 & n4691;
  assign n4717 = ~n3368 & n4699;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = n4715 & n4718;
  assign n4720 = n994 & ~n4719;
  assign n4721 = ~n3504 & n4691;
  assign n4722 = ~n3502 & n4699;
  assign n4723 = n4697 & ~n4722;
  assign n4724 = ~n4721 & n4723;
  assign n4725 = n955 & ~n4724;
  assign n4726 = ~n4720 & ~n4725;
  assign n4727 = ~n4712 & n4726;
  assign n4728 = ~n3189 & n4705;
  assign n4729 = ~n3460 & n4691;
  assign n4730 = ~n3213 & ~n4708;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~n4728 & n4731;
  assign n4733 = n869 & ~n4732;
  assign n4734 = ~n3517 & n4691;
  assign n4735 = ~n3486 & n4699;
  assign n4736 = ~n3364 & n4735;
  assign n4737 = ~n3282 & n4695;
  assign n4738 = ~n3274 & n4693;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = ~n3512 & ~n4739;
  assign n4741 = ~n4736 & ~n4740;
  assign n4742 = ~n4734 & n4741;
  assign n4743 = n924 & ~n4742;
  assign n4744 = ~n4733 & ~n4743;
  assign n4745 = n4727 & n4744;
  assign n4746 = n4704 & n4745;
  assign n4747 = n1381 & ~n4746;
  assign n4748 = n670 & ~n4671;
  assign n4749 = n3087 & ~n3135;
  assign n4750 = ~Pi24 & ~n4677;
  assign n4751 = ~n4749 & n4750;
  assign n4752 = ~n4748 & n4751;
  assign n4753 = ~Pi26 & n3165;
  assign n4754 = ~n3123 & n3158;
  assign n4755 = Pi26 & n4754;
  assign n4756 = n2635 & ~n4755;
  assign n4757 = ~n4753 & n4756;
  assign n4758 = ~n3153 & ~n4757;
  assign n4759 = n670 & ~n4758;
  assign n4760 = ~Pi26 & n4754;
  assign n4761 = Pi26 & n3165;
  assign n4762 = n680 & ~n4761;
  assign n4763 = ~n4760 & n4762;
  assign n4764 = Pi24 & ~n4763;
  assign n4765 = ~n4759 & n4764;
  assign n4766 = ~n4752 & ~n4765;
  assign n4767 = n3087 & ~n3130;
  assign n4768 = ~n3247 & n4693;
  assign n4769 = ~n3231 & n4695;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = ~n3476 & n4691;
  assign n4772 = n4770 & ~n4771;
  assign n4773 = n955 & ~n4772;
  assign n4774 = ~n3213 & ~n4739;
  assign n4775 = ~n3290 & n4691;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n994 & ~n4776;
  assign n4778 = ~n4773 & ~n4777;
  assign n4779 = ~n3322 & n4693;
  assign n4780 = ~n3311 & n4695;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = ~n3471 & n4691;
  assign n4783 = n4781 & ~n4782;
  assign n4784 = n1035 & ~n4783;
  assign n4785 = n4778 & ~n4784;
  assign n4786 = n949 & ~n4280;
  assign n4787 = n3131 & n4300;
  assign n4788 = ~n4786 & n4787;
  assign n4789 = ~Pi24 & ~n4788;
  assign n4790 = ~n4283 & n4699;
  assign n4791 = ~n3488 & n4691;
  assign n4792 = ~n4735 & n4739;
  assign n4793 = ~n4791 & n4792;
  assign n4794 = n924 & ~n4793;
  assign n4795 = ~n3344 & ~n4686;
  assign n4796 = n3126 & ~n4795;
  assign n4797 = ~n4794 & n4796;
  assign n4798 = ~n4790 & n4797;
  assign n4799 = ~n4789 & n4798;
  assign n4800 = ~n3256 & n4699;
  assign n4801 = ~n3262 & n4691;
  assign n4802 = ~n3213 & ~n4770;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = ~n4800 & n4803;
  assign n4805 = n903 & ~n4804;
  assign n4806 = ~n3213 & ~n4781;
  assign n4807 = ~n3330 & n4691;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = n869 & ~n4808;
  assign n4810 = ~n4805 & ~n4809;
  assign n4811 = n4799 & n4810;
  assign n4812 = n4785 & n4811;
  assign n4813 = n1190 & ~n4812;
  assign n4814 = ~n4767 & ~n4813;
  assign n4815 = ~n4766 & n4814;
  assign n4816 = ~n4747 & n4815;
  assign n4817 = n4682 & ~n4816;
  assign n4818 = ~n4680 & ~n4817;
  assign n4819 = ~Ni10 & n4681;
  assign n4820 = ~n637 & ~n3135;
  assign n4821 = n3130 & ~n4820;
  assign n4822 = ~n3120 & ~n4821;
  assign n4823 = ~n637 & n3146;
  assign n4824 = ~n637 & n678;
  assign n4825 = ~n3153 & ~n4824;
  assign n4826 = ~n4823 & ~n4825;
  assign n4827 = ~n637 & n4669;
  assign n4828 = ~Pi23 & n2635;
  assign n4829 = ~n3173 & n4828;
  assign n4830 = ~n4827 & ~n4829;
  assign n4831 = ~n4826 & n4830;
  assign n4832 = n670 & ~n4831;
  assign n4833 = ~n637 & n949;
  assign n4834 = ~n3438 & n4833;
  assign n4835 = ~n3189 & n4834;
  assign n4836 = ~n637 & ~n3131;
  assign n4837 = n3126 & ~n4836;
  assign n4838 = n3213 & n4837;
  assign n4839 = n637 & n949;
  assign n4840 = ~n3443 & n4839;
  assign n4841 = n637 & n867;
  assign n4842 = ~n3452 & n4841;
  assign n4843 = n4837 & ~n4842;
  assign n4844 = ~n4840 & n4843;
  assign n4845 = ~n4838 & ~n4844;
  assign n4846 = ~n637 & n867;
  assign n4847 = ~n3460 & n4846;
  assign n4848 = ~n4845 & ~n4847;
  assign n4849 = ~n4835 & n4848;
  assign n4850 = n736 & ~n4849;
  assign n4851 = ~n3372 & n4846;
  assign n4852 = ~n3377 & n4839;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~n3368 & n4833;
  assign n4855 = ~n3384 & n4841;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = n4837 & n4856;
  assign n4858 = n4853 & n4857;
  assign n4859 = n923 & ~n4858;
  assign n4860 = n730 & ~n4837;
  assign n4861 = n637 & n1030;
  assign n4862 = ~n3427 & n4861;
  assign n4863 = ~n4860 & ~n4862;
  assign n4864 = n3213 & ~n4860;
  assign n4865 = ~n4863 & ~n4864;
  assign n4866 = ~n4859 & ~n4865;
  assign n4867 = ~n3400 & n4833;
  assign n4868 = ~n3412 & n4841;
  assign n4869 = ~n3403 & n4839;
  assign n4870 = n4837 & ~n4869;
  assign n4871 = ~n4868 & n4870;
  assign n4872 = ~n4838 & ~n4871;
  assign n4873 = ~n3420 & n4846;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n4867 & n4874;
  assign n4876 = n738 & ~n4875;
  assign n4877 = ~n637 & n1030;
  assign n4878 = ~n3361 & n4877;
  assign n4879 = ~n4876 & ~n4878;
  assign n4880 = n4866 & n4879;
  assign n4881 = ~n4850 & n4880;
  assign n4882 = n1178 & ~n4881;
  assign n4883 = ~n3207 & n4877;
  assign n4884 = ~n3330 & n4846;
  assign n4885 = ~n3311 & n4839;
  assign n4886 = ~n3322 & n4841;
  assign n4887 = n4837 & ~n4886;
  assign n4888 = ~n4885 & n4887;
  assign n4889 = ~n4838 & ~n4888;
  assign n4890 = ~n3335 & n4833;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~n4884 & n4891;
  assign n4893 = n736 & ~n4892;
  assign n4894 = ~n3256 & n4833;
  assign n4895 = ~n3231 & n4839;
  assign n4896 = ~n3247 & n4841;
  assign n4897 = n4837 & ~n4896;
  assign n4898 = ~n4895 & n4897;
  assign n4899 = ~n4838 & ~n4898;
  assign n4900 = ~n3262 & n4846;
  assign n4901 = ~n4899 & ~n4900;
  assign n4902 = ~n4894 & n4901;
  assign n4903 = n738 & ~n4902;
  assign n4904 = ~n3282 & n4839;
  assign n4905 = ~n3274 & n4841;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = n4837 & n4906;
  assign n4908 = ~n4838 & ~n4907;
  assign n4909 = ~n3290 & n4846;
  assign n4910 = ~n3295 & n4833;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4908 & n4911;
  assign n4913 = n923 & ~n4912;
  assign n4914 = ~n3344 & n4861;
  assign n4915 = ~n4860 & ~n4914;
  assign n4916 = ~n4864 & ~n4915;
  assign n4917 = ~n4913 & ~n4916;
  assign n4918 = ~n4903 & n4917;
  assign n4919 = ~n4893 & n4918;
  assign n4920 = ~n4883 & n4919;
  assign n4921 = n1610 & ~n4920;
  assign n4922 = ~n3471 & n4846;
  assign n4923 = ~n3469 & n4833;
  assign n4924 = n4888 & ~n4923;
  assign n4925 = ~n4922 & n4924;
  assign n4926 = n736 & ~n4925;
  assign n4927 = ~n3486 & n4833;
  assign n4928 = ~n3488 & n4846;
  assign n4929 = n4907 & ~n4928;
  assign n4930 = ~n4927 & n4929;
  assign n4931 = n923 & ~n4930;
  assign n4932 = n4915 & ~n4931;
  assign n4933 = ~n3478 & n4833;
  assign n4934 = ~n3476 & n4846;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = n4898 & n4935;
  assign n4937 = n738 & ~n4936;
  assign n4938 = ~n3484 & n4877;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = n4932 & n4939;
  assign n4941 = ~n4926 & n4940;
  assign n4942 = n1672 & ~n4941;
  assign n4943 = ~n3497 & n4846;
  assign n4944 = ~n4834 & ~n4943;
  assign n4945 = n4844 & n4944;
  assign n4946 = n736 & ~n4945;
  assign n4947 = ~n3512 & ~n4906;
  assign n4948 = ~n3517 & n4846;
  assign n4949 = ~n3364 & n4927;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = n4837 & n4950;
  assign n4952 = ~n4947 & n4951;
  assign n4953 = n923 & ~n4952;
  assign n4954 = n4863 & ~n4953;
  assign n4955 = ~n3502 & n4833;
  assign n4956 = ~n3504 & n4846;
  assign n4957 = ~n4955 & ~n4956;
  assign n4958 = n4871 & n4957;
  assign n4959 = n738 & ~n4958;
  assign n4960 = ~n3510 & n4877;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = n4954 & n4961;
  assign n4963 = ~n4946 & n4962;
  assign n4964 = n1769 & ~n4963;
  assign n4965 = ~n4942 & ~n4964;
  assign n4966 = ~n4921 & n4965;
  assign n4967 = ~n4882 & n4966;
  assign n4968 = n570 & ~n4967;
  assign n4969 = ~n4832 & ~n4968;
  assign n4970 = ~n4822 & n4969;
  assign n4971 = n4819 & ~n4970;
  assign n4972 = n4818 & ~n4971;
  assign n4973 = ~n4591 & n4972;
  assign n4974 = ~n3533 & n4973;
  assign n4975 = n3086 & ~n4974;
  assign n4976 = ~n582 & ~n3135;
  assign n4977 = ~n4667 & ~n4976;
  assign n4978 = ~n579 & n776;
  assign n4979 = ~n4977 & n4978;
  assign n4980 = Ni32 & ~P__cmxcl_1;
  assign n4981 = n580 & n775;
  assign n4982 = ~Ni11 & ~Ni10;
  assign n4983 = ~n4320 & n4982;
  assign n4984 = ~Ni11 & Ni10;
  assign n4985 = ~n3921 & n4984;
  assign n4986 = Ni10 & ~n3851;
  assign n4987 = ~n582 & ~n4986;
  assign n4988 = ~n4225 & n4987;
  assign n4989 = ~n4985 & ~n4988;
  assign n4990 = ~n4983 & n4989;
  assign n4991 = n4981 & ~n4990;
  assign n4992 = ~n4980 & ~n4991;
  assign n4993 = ~n4979 & n4992;
  assign n1012 = n4975 | ~n4993;
  assign n4995 = ~Ni32 & ~Ni30;
  assign n4996 = n864 & n876;
  assign n4997 = P__cmxcl_1 & ~n4996;
  assign n4998 = n4995 & n4997;
  assign n1017_1 = Ni31 | n4998;
  assign n5000 = n872 & ~n875;
  assign n5001 = n1195 & n5000;
  assign n5002 = ~Ni30 & ~n5001;
  assign n5003 = n3854 & ~n5002;
  assign n5004 = P__cmxig_1 & ~n5000;
  assign n5005 = n880 & ~n2107;
  assign n5006 = ~Ni42 & n1054;
  assign n5007 = n5005 & ~n5006;
  assign n5008 = n816 & ~n5007;
  assign n5009 = ~Ni38 & ~n872;
  assign n5010 = n871 & ~n5009;
  assign n5011 = ~n2297 & ~n5007;
  assign n5012 = n5010 & ~n5011;
  assign n5013 = ~n5008 & n5012;
  assign n5014 = ~n5004 & n5013;
  assign n5015 = ~Ni30 & ~n5014;
  assign n5016 = n1643 & ~n5015;
  assign n5017 = n816 & ~n5005;
  assign n5018 = ~Ni30 & n5017;
  assign n5019 = Ni30 & ~n864;
  assign n5020 = ~n1814 & ~n5019;
  assign n5021 = Ni38 & ~n5005;
  assign n5022 = n5010 & ~n5021;
  assign n5023 = ~n5004 & n5022;
  assign n5024 = ~Ni30 & ~n5023;
  assign n5025 = ~n5020 & ~n5024;
  assign n5026 = ~n5018 & n5025;
  assign n5027 = ~Ni42 & n1037;
  assign n5028 = n5005 & ~n5027;
  assign n5029 = n816 & ~n5028;
  assign n5030 = ~Ni30 & n5029;
  assign n5031 = ~n2344 & ~n5028;
  assign n5032 = n5010 & ~n5031;
  assign n5033 = ~n5004 & n5032;
  assign n5034 = ~Ni30 & ~n5033;
  assign n5035 = n1625 & ~n5034;
  assign n5036 = ~n5030 & n5035;
  assign n5037 = ~n5026 & ~n5036;
  assign n5038 = ~n5016 & n5037;
  assign n5039 = n1610 & ~n5038;
  assign n5040 = n816 & ~n880;
  assign n5041 = ~Ni30 & n5040;
  assign n5042 = Ni38 & ~n880;
  assign n5043 = n5010 & ~n5042;
  assign n5044 = ~n5004 & n5043;
  assign n5045 = ~Ni30 & ~n5044;
  assign n5046 = ~n5020 & ~n5045;
  assign n5047 = ~n5041 & n5046;
  assign n5048 = n880 & ~n5027;
  assign n5049 = n816 & ~n5048;
  assign n5050 = ~Ni30 & n5049;
  assign n5051 = ~n2344 & ~n5048;
  assign n5052 = n5010 & ~n5051;
  assign n5053 = ~n5004 & n5052;
  assign n5054 = ~Ni30 & ~n5053;
  assign n5055 = n1625 & ~n5054;
  assign n5056 = ~n5050 & n5055;
  assign n5057 = n880 & ~n5006;
  assign n5058 = n816 & ~n5057;
  assign n5059 = ~Ni30 & n5058;
  assign n5060 = ~n2297 & ~n5057;
  assign n5061 = n5010 & ~n5060;
  assign n5062 = ~n5004 & n5061;
  assign n5063 = ~Ni30 & ~n5062;
  assign n5064 = n1643 & ~n5063;
  assign n5065 = ~n5059 & n5064;
  assign n5066 = ~n5056 & ~n5065;
  assign n5067 = ~n5047 & n5066;
  assign n5068 = n1672 & ~n5067;
  assign n5069 = ~n5046 & ~n5055;
  assign n5070 = ~n5064 & n5069;
  assign n5071 = n1769 & ~n5070;
  assign n5072 = ~n5004 & n5012;
  assign n5073 = ~Ni30 & ~n5072;
  assign n5074 = n1643 & ~n5073;
  assign n5075 = ~n5025 & ~n5035;
  assign n5076 = ~n5074 & n5075;
  assign n5077 = n1178 & ~n5076;
  assign n5078 = ~n5071 & ~n5077;
  assign n5079 = ~n5068 & n5078;
  assign n5080 = ~n5039 & n5079;
  assign n5081 = Pi17 & n5080;
  assign n5082 = ~Ni42 & n957;
  assign n5083 = n880 & ~n5082;
  assign n5084 = n816 & ~n5083;
  assign n5085 = ~Ni30 & n5084;
  assign n5086 = ~n2453 & ~n5083;
  assign n5087 = n5010 & ~n5086;
  assign n5088 = ~n5004 & n5087;
  assign n5089 = ~Ni30 & ~n5088;
  assign n5090 = n1636 & ~n5089;
  assign n5091 = ~n5085 & n5090;
  assign n5092 = ~Ni32 & n816;
  assign n5093 = n870 & n5092;
  assign n5094 = ~n5010 & ~n5093;
  assign n5095 = n880 & ~n1005;
  assign n5096 = ~Ni38 & ~n891;
  assign n5097 = ~n816 & n5096;
  assign n5098 = ~n5095 & ~n5097;
  assign n5099 = ~n5094 & ~n5098;
  assign n5100 = ~n5004 & n5099;
  assign n5101 = ~Ni30 & ~n5100;
  assign n5102 = n1625 & ~n5101;
  assign n5103 = Ni44 & n2333;
  assign n5104 = n880 & ~n5103;
  assign n5105 = ~Ni38 & ~n938;
  assign n5106 = ~n816 & n5105;
  assign n5107 = ~n5104 & ~n5106;
  assign n5108 = ~n5094 & ~n5107;
  assign n5109 = ~n5004 & n5108;
  assign n5110 = ~Ni30 & ~n5109;
  assign n5111 = n1643 & ~n5110;
  assign n5112 = ~n5102 & ~n5111;
  assign n5113 = n973 & n2333;
  assign n5114 = n880 & ~n5113;
  assign n5115 = n816 & ~n5114;
  assign n5116 = ~n2380 & ~n5114;
  assign n5117 = n5010 & ~n5116;
  assign n5118 = ~n5115 & n5117;
  assign n5119 = ~n5004 & n5118;
  assign n5120 = ~Ni30 & ~n5119;
  assign n5121 = ~n1611 & ~n5019;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = n5112 & ~n5122;
  assign n5124 = ~n5091 & n5123;
  assign n5125 = n1672 & ~n5124;
  assign n5126 = n5005 & ~n5113;
  assign n5127 = ~n2380 & ~n5126;
  assign n5128 = n5010 & ~n5127;
  assign n5129 = ~n5004 & n5128;
  assign n5130 = ~Ni30 & ~n5129;
  assign n5131 = n816 & ~n5126;
  assign n5132 = ~Ni30 & n5131;
  assign n5133 = ~n5130 & ~n5132;
  assign n5134 = n1611 & n5133;
  assign n5135 = n5005 & ~n5103;
  assign n5136 = ~n5106 & ~n5135;
  assign n5137 = ~n5094 & ~n5136;
  assign n5138 = ~n5004 & n5137;
  assign n5139 = ~Ni30 & ~n5138;
  assign n5140 = n1643 & ~n5139;
  assign n5141 = ~n1005 & n5005;
  assign n5142 = ~n5097 & ~n5141;
  assign n5143 = ~n5094 & ~n5142;
  assign n5144 = ~n5004 & n5143;
  assign n5145 = ~Ni30 & ~n5144;
  assign n5146 = n1625 & ~n5145;
  assign n5147 = ~n5140 & ~n5146;
  assign n5148 = ~n2107 & n5083;
  assign n5149 = n816 & ~n5148;
  assign n5150 = ~Ni30 & n5149;
  assign n5151 = ~n2453 & ~n5148;
  assign n5152 = n5010 & ~n5151;
  assign n5153 = ~n5004 & n5152;
  assign n5154 = ~Ni30 & ~n5153;
  assign n5155 = ~n5150 & ~n5154;
  assign n5156 = ~n1636 & ~n5019;
  assign n5157 = n5155 & ~n5156;
  assign n5158 = n5147 & ~n5157;
  assign n5159 = ~n5134 & n5158;
  assign n5160 = n1610 & ~n5159;
  assign n5161 = n1636 & ~n5154;
  assign n5162 = ~n5096 & ~n5141;
  assign n5163 = n5010 & ~n5162;
  assign n5164 = ~n5004 & n5163;
  assign n5165 = ~Ni30 & ~n5164;
  assign n5166 = n1625 & ~n5165;
  assign n5167 = ~n5105 & ~n5135;
  assign n5168 = n5010 & ~n5167;
  assign n5169 = ~n5004 & n5168;
  assign n5170 = ~Ni30 & ~n5169;
  assign n5171 = n1643 & ~n5170;
  assign n5172 = ~n5166 & ~n5171;
  assign n5173 = ~n5121 & ~n5130;
  assign n5174 = n5172 & ~n5173;
  assign n5175 = ~n5161 & n5174;
  assign n5176 = n1178 & ~n5175;
  assign n5177 = ~n5160 & ~n5176;
  assign n5178 = ~n5125 & n5177;
  assign n5179 = ~n5095 & ~n5096;
  assign n5180 = n5010 & ~n5179;
  assign n5181 = ~n5004 & n5180;
  assign n5182 = ~Ni30 & ~n5181;
  assign n5183 = n1625 & ~n5182;
  assign n5184 = ~n5004 & n5117;
  assign n5185 = ~Ni30 & ~n5184;
  assign n5186 = n1611 & ~n5185;
  assign n5187 = ~n5104 & ~n5105;
  assign n5188 = n5010 & ~n5187;
  assign n5189 = ~n5004 & n5188;
  assign n5190 = ~Ni30 & ~n5189;
  assign n5191 = ~n1643 & ~n5019;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = ~n5186 & ~n5192;
  assign n5194 = ~n5090 & n5193;
  assign n5195 = ~n5183 & n5194;
  assign n5196 = n1769 & ~n5195;
  assign n5197 = ~Pi17 & ~n5196;
  assign n5198 = n5178 & n5197;
  assign n5199 = n679 & ~n5198;
  assign n5200 = ~n5081 & n5199;
  assign n5201 = ~n5003 & ~n5200;
  assign n5202 = ~Ni11 & ~n5201;
  assign n5203 = ~n582 & ~n5002;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = n4978 & ~n5204;
  assign n5206 = ~n865 & ~n5002;
  assign n5207 = ~Ni30 & ~n5022;
  assign n5208 = Pi16 & n5043;
  assign n5209 = n5207 & ~n5208;
  assign n5210 = n1031 & ~n5209;
  assign n5211 = ~Pi20 & n5087;
  assign n5212 = ~Pi20 & ~Ni30;
  assign n5213 = ~Ni30 & ~n5117;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = ~n5211 & ~n5214;
  assign n5216 = n955 & ~n5215;
  assign n5217 = ~n5152 & n5212;
  assign n5218 = Pi20 & ~Ni30;
  assign n5219 = ~n5128 & n5218;
  assign n5220 = ~n5217 & ~n5219;
  assign n5221 = n903 & n5220;
  assign n5222 = ~n5052 & n5212;
  assign n5223 = ~n5061 & n5218;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = n1035 & n5224;
  assign n5226 = ~n5221 & ~n5225;
  assign n5227 = ~n5032 & n5212;
  assign n5228 = ~n5012 & n5218;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = n869 & n5229;
  assign n5231 = ~n5168 & n5218;
  assign n5232 = ~n5163 & n5212;
  assign n5233 = ~n5231 & ~n5232;
  assign n5234 = n994 & n5233;
  assign n5235 = ~n5188 & n5218;
  assign n5236 = ~n5180 & n5212;
  assign n5237 = ~n5235 & ~n5236;
  assign n5238 = n924 & n5237;
  assign n5239 = ~n5234 & ~n5238;
  assign n5240 = ~n5230 & n5239;
  assign n5241 = n5226 & n5240;
  assign n5242 = ~n5216 & n5241;
  assign n5243 = n865 & ~n5242;
  assign n5244 = Pi15 & ~n5243;
  assign n5245 = ~n5210 & n5244;
  assign n5246 = ~n5040 & n5208;
  assign n5247 = ~n5018 & ~n5207;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n1031 & ~n5248;
  assign n5250 = ~n5084 & n5211;
  assign n5251 = ~Ni30 & ~n5118;
  assign n5252 = ~n5212 & ~n5251;
  assign n5253 = ~n5250 & ~n5252;
  assign n5254 = n955 & ~n5253;
  assign n5255 = ~n5029 & n5032;
  assign n5256 = n5212 & ~n5255;
  assign n5257 = ~n5013 & n5218;
  assign n5258 = ~n5256 & ~n5257;
  assign n5259 = n869 & n5258;
  assign n5260 = ~n5143 & n5212;
  assign n5261 = ~n5137 & n5218;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = n994 & n5262;
  assign n5264 = ~n5259 & ~n5263;
  assign n5265 = ~n5149 & n5152;
  assign n5266 = n5212 & ~n5265;
  assign n5267 = n5128 & ~n5131;
  assign n5268 = n5218 & ~n5267;
  assign n5269 = ~n5266 & ~n5268;
  assign n5270 = n903 & n5269;
  assign n5271 = ~n5049 & n5052;
  assign n5272 = n5212 & ~n5271;
  assign n5273 = ~n5058 & n5061;
  assign n5274 = n5218 & ~n5273;
  assign n5275 = ~n5272 & ~n5274;
  assign n5276 = n1035 & n5275;
  assign n5277 = ~n5270 & ~n5276;
  assign n5278 = ~n5099 & n5212;
  assign n5279 = ~n5108 & n5218;
  assign n5280 = ~n5278 & ~n5279;
  assign n5281 = n924 & n5280;
  assign n5282 = n5277 & ~n5281;
  assign n5283 = n5264 & n5282;
  assign n5284 = ~n5254 & n5283;
  assign n5285 = n865 & ~n5284;
  assign n5286 = ~Pi15 & ~n5285;
  assign n5287 = ~n5249 & n5286;
  assign n5288 = ~n5245 & ~n5287;
  assign n5289 = ~n5206 & ~n5288;
  assign n5290 = n3854 & ~n5289;
  assign n5291 = n903 & n5155;
  assign n5292 = n1035 & ~n5054;
  assign n5293 = ~n5050 & n5292;
  assign n5294 = ~n5291 & ~n5293;
  assign n5295 = n4230 & ~n5294;
  assign n5296 = n4265 & ~n5089;
  assign n5297 = ~n5085 & n5296;
  assign n5298 = n994 & n4232;
  assign n5299 = ~n5139 & n5298;
  assign n5300 = ~n5297 & ~n5299;
  assign n5301 = n1528 & ~n5045;
  assign n5302 = ~n5041 & n5301;
  assign n5303 = n2205 & ~n5024;
  assign n5304 = ~n5018 & n5303;
  assign n5305 = ~n5302 & ~n5304;
  assign n5306 = n4308 & ~n5145;
  assign n5307 = n5305 & ~n5306;
  assign n5308 = n5300 & n5307;
  assign n5309 = n1035 & ~n5063;
  assign n5310 = ~n5059 & n5309;
  assign n5311 = n924 & ~n5110;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = n955 & ~n5120;
  assign n5314 = n903 & ~n5130;
  assign n5315 = ~n5132 & n5314;
  assign n5316 = ~n5313 & ~n5315;
  assign n5317 = n869 & ~n5015;
  assign n5318 = n5316 & ~n5317;
  assign n5319 = n5312 & n5318;
  assign n5320 = n4232 & ~n5319;
  assign n5321 = n4240 & ~n5034;
  assign n5322 = ~n5030 & n5321;
  assign n5323 = ~n4295 & ~n5019;
  assign n5324 = ~n5101 & ~n5323;
  assign n5325 = ~n5322 & ~n5324;
  assign n5326 = ~n5320 & n5325;
  assign n5327 = n5308 & n5326;
  assign n5328 = ~n5295 & n5327;
  assign n5329 = n5287 & n5328;
  assign n5330 = n869 & ~n5073;
  assign n5331 = n955 & ~n5185;
  assign n5332 = n924 & ~n5190;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5330 & n5333;
  assign n5335 = n4232 & ~n5334;
  assign n5336 = n4230 & ~n5154;
  assign n5337 = n4232 & ~n5130;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = n903 & ~n5338;
  assign n5340 = n4230 & n5292;
  assign n5341 = ~n5182 & ~n5323;
  assign n5342 = ~n5340 & ~n5341;
  assign n5343 = n4308 & ~n5165;
  assign n5344 = n5342 & ~n5343;
  assign n5345 = ~n5301 & ~n5303;
  assign n5346 = ~n5170 & n5298;
  assign n5347 = n5345 & ~n5346;
  assign n5348 = ~n5296 & n5347;
  assign n5349 = ~n5321 & n5348;
  assign n5350 = n4232 & n5309;
  assign n5351 = n5349 & ~n5350;
  assign n5352 = n5344 & n5351;
  assign n5353 = ~n5339 & n5352;
  assign n5354 = n5245 & n5353;
  assign n5355 = ~n5335 & n5354;
  assign n5356 = n679 & ~n5355;
  assign n5357 = ~n5329 & n5356;
  assign n5358 = ~n5290 & ~n5357;
  assign n5359 = n4982 & ~n5358;
  assign n5360 = ~n652 & ~n3121;
  assign n5361 = ~n5267 & n5360;
  assign n5362 = P__cmxig_0 & ~n5000;
  assign n5363 = n5360 & n5362;
  assign n5364 = ~n5361 & ~n5363;
  assign n5365 = n3560 & n5364;
  assign n5366 = ~n5265 & n5360;
  assign n5367 = ~n5363 & ~n5366;
  assign n5368 = n3556 & n5367;
  assign n5369 = ~n5365 & ~n5368;
  assign n5370 = Ni30 & ~n769;
  assign n5371 = ~n652 & ~n5370;
  assign n5372 = Pi26 & Ni30;
  assign n5373 = n5371 & ~n5372;
  assign n5374 = ~n864 & ~n5373;
  assign n5375 = ~Ni30 & n5362;
  assign n5376 = ~Ni30 & ~n5152;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = n3552 & n5377;
  assign n5379 = ~n5150 & n5378;
  assign n5380 = n5128 & ~n5362;
  assign n5381 = ~Ni30 & ~n5380;
  assign n5382 = n3547 & ~n5381;
  assign n5383 = ~n5132 & n5382;
  assign n5384 = ~n5379 & ~n5383;
  assign n5385 = ~n5374 & n5384;
  assign n5386 = n5369 & n5385;
  assign n5387 = n738 & ~n5386;
  assign n5388 = n730 & n5374;
  assign n5389 = ~n736 & ~n5388;
  assign n5390 = ~n5255 & n5360;
  assign n5391 = ~n5363 & ~n5390;
  assign n5392 = n3556 & n5391;
  assign n5393 = n5013 & ~n5362;
  assign n5394 = ~Ni30 & ~n5393;
  assign n5395 = n3547 & ~n5394;
  assign n5396 = n5360 & ~n5393;
  assign n5397 = n3560 & ~n5396;
  assign n5398 = ~n5395 & ~n5397;
  assign n5399 = n5032 & ~n5362;
  assign n5400 = ~Ni30 & ~n5399;
  assign n5401 = n3552 & ~n5400;
  assign n5402 = ~n5030 & n5401;
  assign n5403 = n5398 & ~n5402;
  assign n5404 = ~n5392 & n5403;
  assign n5405 = ~n5374 & n5404;
  assign n5406 = ~n5389 & ~n5405;
  assign n5407 = ~n5207 & ~n5375;
  assign n5408 = n3540 & n5407;
  assign n5409 = ~n5018 & n5408;
  assign n5410 = n5143 & ~n5362;
  assign n5411 = n5360 & ~n5410;
  assign n5412 = n3556 & ~n5411;
  assign n5413 = n5137 & ~n5362;
  assign n5414 = n5360 & ~n5413;
  assign n5415 = n3560 & ~n5414;
  assign n5416 = ~Ni30 & ~n5410;
  assign n5417 = n3552 & ~n5416;
  assign n5418 = ~n5415 & ~n5417;
  assign n5419 = ~Ni30 & ~n5413;
  assign n5420 = n3547 & ~n5419;
  assign n5421 = ~n5374 & ~n5420;
  assign n5422 = n5418 & n5421;
  assign n5423 = ~n5412 & n5422;
  assign n5424 = n923 & ~n5423;
  assign n5425 = n5017 & n5360;
  assign n5426 = ~n5022 & n5360;
  assign n5427 = ~n5363 & ~n5426;
  assign n5428 = n3605 & n5427;
  assign n5429 = ~n5425 & n5428;
  assign n5430 = ~n5424 & ~n5429;
  assign n5431 = ~n5409 & n5430;
  assign n5432 = ~n5406 & n5431;
  assign n5433 = ~n5387 & n5432;
  assign n5434 = n1610 & ~n5433;
  assign n5435 = n5087 & ~n5362;
  assign n5436 = ~Ni30 & ~n5435;
  assign n5437 = n3552 & ~n5436;
  assign n5438 = ~n5213 & ~n5375;
  assign n5439 = n3547 & n5438;
  assign n5440 = ~n5437 & ~n5439;
  assign n5441 = n5360 & ~n5435;
  assign n5442 = n3556 & ~n5441;
  assign n5443 = ~n5117 & n5360;
  assign n5444 = ~n5363 & ~n5443;
  assign n5445 = n3560 & n5444;
  assign n5446 = ~n5442 & ~n5445;
  assign n5447 = n5440 & n5446;
  assign n5448 = ~n5374 & n5447;
  assign n5449 = n738 & ~n5448;
  assign n5450 = ~Ni30 & ~n5043;
  assign n5451 = ~n5375 & ~n5450;
  assign n5452 = n3540 & n5451;
  assign n5453 = ~n5061 & n5360;
  assign n5454 = ~n5363 & ~n5453;
  assign n5455 = n3560 & n5454;
  assign n5456 = ~n5374 & ~n5455;
  assign n5457 = n5052 & ~n5362;
  assign n5458 = ~Ni30 & ~n5457;
  assign n5459 = n3552 & ~n5458;
  assign n5460 = ~n5052 & n5360;
  assign n5461 = ~n5363 & ~n5460;
  assign n5462 = n3556 & n5461;
  assign n5463 = ~n5459 & ~n5462;
  assign n5464 = n5061 & ~n5362;
  assign n5465 = ~Ni30 & ~n5464;
  assign n5466 = n3547 & ~n5465;
  assign n5467 = n5463 & ~n5466;
  assign n5468 = n5456 & n5467;
  assign n5469 = n736 & ~n5468;
  assign n5470 = ~n5043 & n5360;
  assign n5471 = ~n5363 & ~n5470;
  assign n5472 = n3605 & n5471;
  assign n5473 = ~n923 & ~n5388;
  assign n5474 = n5188 & ~n5362;
  assign n5475 = ~Ni30 & ~n5474;
  assign n5476 = n3547 & ~n5475;
  assign n5477 = ~n5180 & n5360;
  assign n5478 = ~n5363 & ~n5477;
  assign n5479 = n3556 & n5478;
  assign n5480 = ~n5374 & ~n5479;
  assign n5481 = ~Ni30 & ~n5180;
  assign n5482 = ~n5375 & ~n5481;
  assign n5483 = n3552 & n5482;
  assign n5484 = ~n5188 & n5360;
  assign n5485 = ~n5363 & ~n5484;
  assign n5486 = n3560 & n5485;
  assign n5487 = ~n5483 & ~n5486;
  assign n5488 = n5480 & n5487;
  assign n5489 = ~n5476 & n5488;
  assign n5490 = ~n5473 & ~n5489;
  assign n5491 = ~n5472 & ~n5490;
  assign n5492 = ~n5469 & n5491;
  assign n5493 = ~n5452 & n5492;
  assign n5494 = ~n5449 & n5493;
  assign n5495 = n1769 & ~n5494;
  assign n5496 = ~n5374 & ~n5382;
  assign n5497 = ~n5152 & n5360;
  assign n5498 = ~n5363 & ~n5497;
  assign n5499 = n3556 & n5498;
  assign n5500 = n5496 & ~n5499;
  assign n5501 = ~n5128 & n5360;
  assign n5502 = ~n5363 & ~n5501;
  assign n5503 = n3560 & n5502;
  assign n5504 = ~n5378 & ~n5503;
  assign n5505 = n5500 & n5504;
  assign n5506 = n738 & ~n5505;
  assign n5507 = ~n5408 & ~n5506;
  assign n5508 = n5012 & ~n5362;
  assign n5509 = n5360 & ~n5508;
  assign n5510 = n3560 & ~n5509;
  assign n5511 = n5360 & ~n5399;
  assign n5512 = n3556 & ~n5511;
  assign n5513 = ~n5401 & ~n5512;
  assign n5514 = ~Ni30 & ~n5508;
  assign n5515 = n3547 & ~n5514;
  assign n5516 = ~n5374 & ~n5515;
  assign n5517 = n5513 & n5516;
  assign n5518 = ~n5510 & n5517;
  assign n5519 = ~n5389 & ~n5518;
  assign n5520 = ~Ni30 & ~n5163;
  assign n5521 = ~n5375 & ~n5520;
  assign n5522 = n3552 & n5521;
  assign n5523 = ~Ni30 & ~n5168;
  assign n5524 = ~n5375 & ~n5523;
  assign n5525 = n3547 & n5524;
  assign n5526 = ~n5522 & ~n5525;
  assign n5527 = ~n5168 & n5360;
  assign n5528 = ~n5363 & ~n5527;
  assign n5529 = n3560 & n5528;
  assign n5530 = ~n5163 & n5360;
  assign n5531 = ~n5363 & ~n5530;
  assign n5532 = n3556 & n5531;
  assign n5533 = ~n5529 & ~n5532;
  assign n5534 = n5526 & n5533;
  assign n5535 = ~n5374 & n5534;
  assign n5536 = n923 & ~n5535;
  assign n5537 = ~n5428 & ~n5536;
  assign n5538 = ~n5519 & n5537;
  assign n5539 = n5507 & n5538;
  assign n5540 = n1178 & ~n5539;
  assign n5541 = n5040 & n5360;
  assign n5542 = n5472 & ~n5541;
  assign n5543 = ~n5059 & n5466;
  assign n5544 = ~n5271 & n5360;
  assign n5545 = ~n5363 & ~n5544;
  assign n5546 = n3556 & n5545;
  assign n5547 = ~n5543 & ~n5546;
  assign n5548 = ~n5050 & n5459;
  assign n5549 = ~n5374 & ~n5548;
  assign n5550 = ~n5273 & n5360;
  assign n5551 = ~n5363 & ~n5550;
  assign n5552 = n3560 & n5551;
  assign n5553 = n5549 & ~n5552;
  assign n5554 = n5547 & n5553;
  assign n5555 = n736 & ~n5554;
  assign n5556 = ~n5118 & n5360;
  assign n5557 = ~n5363 & ~n5556;
  assign n5558 = n3560 & n5557;
  assign n5559 = n5084 & n5360;
  assign n5560 = n5442 & ~n5559;
  assign n5561 = ~n5251 & ~n5375;
  assign n5562 = n3547 & n5561;
  assign n5563 = ~n5560 & ~n5562;
  assign n5564 = ~n5085 & n5437;
  assign n5565 = ~n5374 & ~n5564;
  assign n5566 = n5563 & n5565;
  assign n5567 = ~n5558 & n5566;
  assign n5568 = n738 & ~n5567;
  assign n5569 = n5108 & ~n5362;
  assign n5570 = n5360 & ~n5569;
  assign n5571 = n3560 & ~n5570;
  assign n5572 = ~Ni30 & ~n5569;
  assign n5573 = n3547 & ~n5572;
  assign n5574 = n5099 & ~n5362;
  assign n5575 = ~Ni30 & ~n5574;
  assign n5576 = n3552 & ~n5575;
  assign n5577 = ~n5573 & ~n5576;
  assign n5578 = n5360 & ~n5574;
  assign n5579 = n3556 & ~n5578;
  assign n5580 = n5577 & ~n5579;
  assign n5581 = ~n5571 & n5580;
  assign n5582 = ~n5374 & n5581;
  assign n5583 = ~n5473 & ~n5582;
  assign n5584 = ~n5041 & n5451;
  assign n5585 = n3540 & n5584;
  assign n5586 = ~n5583 & ~n5585;
  assign n5587 = ~n5568 & n5586;
  assign n5588 = ~n5555 & n5587;
  assign n5589 = ~n5542 & n5588;
  assign n5590 = n1672 & ~n5589;
  assign n5591 = ~n5540 & ~n5590;
  assign n5592 = ~n5495 & n5591;
  assign n5593 = ~n5434 & n5592;
  assign n5594 = n3534 & ~n5593;
  assign n5595 = n1625 & ~n5400;
  assign n5596 = n1643 & ~n5514;
  assign n5597 = ~n5020 & n5407;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = ~n5595 & n5598;
  assign n5600 = n1178 & ~n5599;
  assign n5601 = n1625 & ~n5458;
  assign n5602 = ~n5050 & n5601;
  assign n5603 = ~n5191 & ~n5465;
  assign n5604 = ~n5059 & n5603;
  assign n5605 = ~n5602 & ~n5604;
  assign n5606 = n1672 & ~n5605;
  assign n5607 = ~n5600 & ~n5606;
  assign n5608 = n1814 & n5451;
  assign n5609 = ~n5601 & ~n5603;
  assign n5610 = ~n5608 & n5609;
  assign n5611 = n1769 & ~n5610;
  assign n5612 = n1878 & n5584;
  assign n5613 = ~n5018 & n5407;
  assign n5614 = n2872 & n5613;
  assign n5615 = Pi17 & ~n5614;
  assign n5616 = ~n5612 & n5615;
  assign n5617 = ~n5191 & ~n5394;
  assign n5618 = ~n5030 & n5595;
  assign n5619 = ~n5617 & ~n5618;
  assign n5620 = n1610 & ~n5619;
  assign n5621 = n5616 & ~n5620;
  assign n5622 = ~n5611 & n5621;
  assign n5623 = n5607 & n5622;
  assign n5624 = n1625 & n5521;
  assign n5625 = n1636 & n5377;
  assign n5626 = n1611 & ~n5381;
  assign n5627 = ~n5191 & n5524;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = ~n5625 & n5628;
  assign n5630 = ~n5624 & n5629;
  assign n5631 = n1178 & ~n5630;
  assign n5632 = ~n5132 & n5626;
  assign n5633 = ~n5191 & ~n5419;
  assign n5634 = n1625 & ~n5416;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = ~n5150 & n5625;
  assign n5637 = n5635 & ~n5636;
  assign n5638 = ~n5632 & n5637;
  assign n5639 = n1610 & ~n5638;
  assign n5640 = ~n5156 & ~n5436;
  assign n5641 = ~n5085 & n5640;
  assign n5642 = n1625 & ~n5575;
  assign n5643 = n1643 & ~n5572;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = n1611 & n5561;
  assign n5646 = n5644 & ~n5645;
  assign n5647 = ~n5641 & n5646;
  assign n5648 = n1672 & ~n5647;
  assign n5649 = n1643 & ~n5475;
  assign n5650 = n1625 & n5482;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = n1611 & n5438;
  assign n5653 = n5651 & ~n5652;
  assign n5654 = ~n5640 & n5653;
  assign n5655 = n1769 & ~n5654;
  assign n5656 = ~Pi17 & ~n5655;
  assign n5657 = ~n5648 & n5656;
  assign n5658 = ~n5639 & n5657;
  assign n5659 = ~n5631 & n5658;
  assign n5660 = ~n5623 & ~n5659;
  assign n5661 = n3854 & n5660;
  assign n5662 = n1769 & n5224;
  assign n5663 = n1178 & n5229;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = ~n5258 & n5664;
  assign n5666 = n1672 & n5275;
  assign n5667 = Pi17 & ~n5666;
  assign n5668 = n5665 & n5667;
  assign n5669 = n1178 & n5233;
  assign n5670 = n1672 & n5280;
  assign n5671 = n1769 & n5237;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = ~n5262 & n5672;
  assign n5674 = ~n5669 & n5673;
  assign n5675 = ~Pi17 & n5674;
  assign n5676 = n1624 & ~n5675;
  assign n5677 = ~n5668 & n5676;
  assign n5678 = n1672 & ~n5253;
  assign n5679 = n1769 & ~n5215;
  assign n5680 = n1178 & n5220;
  assign n5681 = ~n5269 & ~n5680;
  assign n5682 = ~n5679 & n5681;
  assign n5683 = ~n5678 & n5682;
  assign n5684 = ~Pi17 & n5683;
  assign n5685 = ~Pi15 & n5041;
  assign n5686 = Pi16 & ~n5685;
  assign n5687 = ~n5450 & n5686;
  assign n5688 = ~n1178 & n5018;
  assign n5689 = ~n5207 & ~n5688;
  assign n5690 = ~n5687 & ~n5689;
  assign n5691 = Pi17 & n5690;
  assign n5692 = n1814 & ~n5691;
  assign n5693 = ~n5684 & n5692;
  assign n5694 = ~n5677 & ~n5693;
  assign n5695 = ~n5019 & n5694;
  assign n5696 = n679 & ~n5695;
  assign n5697 = ~n5661 & ~n5696;
  assign n5698 = ~n3096 & n5360;
  assign n5699 = ~n864 & ~n5698;
  assign n5700 = n3930 & ~n5458;
  assign n5701 = ~n5050 & n5700;
  assign n5702 = n3922 & n5545;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = n3928 & ~n5465;
  assign n5705 = ~n5059 & n5704;
  assign n5706 = n3924 & n5551;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = n5703 & n5707;
  assign n5709 = n1035 & ~n5708;
  assign n5710 = n3942 & n5407;
  assign n5711 = ~n5018 & n5710;
  assign n5712 = ~n5709 & ~n5711;
  assign n5713 = n3928 & ~n5394;
  assign n5714 = n3930 & ~n5400;
  assign n5715 = ~n5030 & n5714;
  assign n5716 = n3924 & ~n5396;
  assign n5717 = ~n5715 & ~n5716;
  assign n5718 = n3922 & n5391;
  assign n5719 = n5717 & ~n5718;
  assign n5720 = ~n5713 & n5719;
  assign n5721 = n869 & ~n5720;
  assign n5722 = n3922 & ~n5578;
  assign n5723 = n3928 & ~n5572;
  assign n5724 = n3930 & ~n5575;
  assign n5725 = n3924 & ~n5570;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n5723 & n5726;
  assign n5728 = ~n5722 & n5727;
  assign n5729 = n924 & ~n5728;
  assign n5730 = n3944 & n5471;
  assign n5731 = ~n5541 & n5730;
  assign n5732 = ~n5729 & ~n5731;
  assign n5733 = ~n5721 & n5732;
  assign n5734 = n5712 & n5733;
  assign n5735 = n3930 & n5377;
  assign n5736 = ~n5150 & n5735;
  assign n5737 = n3924 & n5364;
  assign n5738 = n3922 & n5367;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = n3928 & ~n5381;
  assign n5741 = ~n5132 & n5740;
  assign n5742 = n5739 & ~n5741;
  assign n5743 = ~n5736 & n5742;
  assign n5744 = n903 & ~n5743;
  assign n5745 = n3924 & ~n5414;
  assign n5746 = n3928 & ~n5419;
  assign n5747 = n3930 & ~n5416;
  assign n5748 = n3922 & ~n5411;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = ~n5746 & n5749;
  assign n5751 = ~n5745 & n5750;
  assign n5752 = n994 & ~n5751;
  assign n5753 = n3949 & n5451;
  assign n5754 = ~Pi15 & ~n5753;
  assign n5755 = ~n5685 & ~n5754;
  assign n5756 = ~n5752 & ~n5755;
  assign n5757 = ~n5744 & n5756;
  assign n5758 = n3928 & n5561;
  assign n5759 = n3924 & n5557;
  assign n5760 = n3922 & ~n5441;
  assign n5761 = ~n5559 & n5760;
  assign n5762 = n3930 & ~n5436;
  assign n5763 = ~n5085 & n5762;
  assign n5764 = ~n5761 & ~n5763;
  assign n5765 = ~n5759 & n5764;
  assign n5766 = ~n5758 & n5765;
  assign n5767 = n955 & ~n5766;
  assign n5768 = n3945 & n5427;
  assign n5769 = ~n5425 & n5768;
  assign n5770 = ~n5767 & ~n5769;
  assign n5771 = n5757 & n5770;
  assign n5772 = n5734 & n5771;
  assign n5773 = n3924 & n5444;
  assign n5774 = n3928 & n5438;
  assign n5775 = ~n5760 & ~n5774;
  assign n5776 = ~n5773 & n5775;
  assign n5777 = ~n5762 & n5776;
  assign n5778 = n955 & ~n5777;
  assign n5779 = n3922 & ~n5511;
  assign n5780 = n3924 & ~n5509;
  assign n5781 = n3928 & ~n5514;
  assign n5782 = ~n5780 & ~n5781;
  assign n5783 = ~n5714 & n5782;
  assign n5784 = ~n5779 & n5783;
  assign n5785 = n869 & ~n5784;
  assign n5786 = n3924 & n5502;
  assign n5787 = n3922 & n5498;
  assign n5788 = ~n5735 & ~n5787;
  assign n5789 = ~n5740 & n5788;
  assign n5790 = ~n5786 & n5789;
  assign n5791 = n903 & ~n5790;
  assign n5792 = ~n5785 & ~n5791;
  assign n5793 = n3922 & n5461;
  assign n5794 = n3924 & n5454;
  assign n5795 = ~n5704 & ~n5794;
  assign n5796 = ~n5793 & n5795;
  assign n5797 = ~n5700 & n5796;
  assign n5798 = n1035 & ~n5797;
  assign n5799 = n3922 & n5478;
  assign n5800 = n3928 & ~n5475;
  assign n5801 = n3930 & n5482;
  assign n5802 = n3924 & n5485;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804 = ~n5800 & n5803;
  assign n5805 = ~n5799 & n5804;
  assign n5806 = n924 & ~n5805;
  assign n5807 = n3930 & n5521;
  assign n5808 = n3928 & n5524;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = n3922 & n5531;
  assign n5811 = n3924 & n5528;
  assign n5812 = ~n5810 & ~n5811;
  assign n5813 = n5809 & n5812;
  assign n5814 = n994 & ~n5813;
  assign n5815 = Pi15 & ~n5753;
  assign n5816 = ~n5768 & n5815;
  assign n5817 = ~n5710 & n5816;
  assign n5818 = ~n5730 & n5817;
  assign n5819 = ~n5814 & n5818;
  assign n5820 = ~n5806 & n5819;
  assign n5821 = ~n5798 & n5820;
  assign n5822 = n5792 & n5821;
  assign n5823 = ~n5778 & n5822;
  assign n5824 = ~n5772 & ~n5823;
  assign n5825 = ~n5699 & ~n5824;
  assign n5826 = n4046 & ~n5825;
  assign n5827 = n3852 & n5660;
  assign n5828 = ~n5826 & ~n5827;
  assign n5829 = n5697 & n5828;
  assign n5830 = ~n5594 & n5829;
  assign n5831 = ~Ni11 & ~n5830;
  assign n5832 = ~Pi26 & Ni30;
  assign n5833 = n5371 & ~n5832;
  assign n5834 = ~n864 & ~n5833;
  assign n5835 = n4062 & ~n5400;
  assign n5836 = ~n5030 & n5835;
  assign n5837 = n4059 & n5391;
  assign n5838 = ~n5836 & ~n5837;
  assign n5839 = n4057 & ~n5396;
  assign n5840 = n4065 & ~n5394;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = n5838 & n5841;
  assign n5843 = ~n5834 & n5842;
  assign n5844 = n736 & ~n5843;
  assign n5845 = n4065 & ~n5381;
  assign n5846 = ~n5132 & n5845;
  assign n5847 = n4059 & n5367;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = n4057 & n5364;
  assign n5850 = n4062 & n5377;
  assign n5851 = ~n5150 & n5850;
  assign n5852 = ~n5849 & ~n5851;
  assign n5853 = n5848 & n5852;
  assign n5854 = ~n5834 & n5853;
  assign n5855 = n738 & ~n5854;
  assign n5856 = n730 & n5834;
  assign n5857 = ~n923 & ~n5856;
  assign n5858 = n4062 & ~n5416;
  assign n5859 = n4059 & ~n5411;
  assign n5860 = n4065 & ~n5419;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = n4057 & ~n5414;
  assign n5863 = n5861 & ~n5862;
  assign n5864 = ~n5858 & n5863;
  assign n5865 = ~n5834 & n5864;
  assign n5866 = ~n5857 & ~n5865;
  assign n5867 = ~n5855 & ~n5866;
  assign n5868 = n4053 & n5427;
  assign n5869 = ~n5425 & n5868;
  assign n5870 = n4089 & n5613;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = n5867 & n5871;
  assign n5873 = ~n5844 & n5872;
  assign n5874 = n1610 & ~n5873;
  assign n5875 = n4059 & ~n5511;
  assign n5876 = n4057 & ~n5509;
  assign n5877 = n4065 & ~n5514;
  assign n5878 = ~n5834 & ~n5877;
  assign n5879 = ~n5876 & n5878;
  assign n5880 = ~n5875 & n5879;
  assign n5881 = ~n5835 & n5880;
  assign n5882 = n736 & ~n5881;
  assign n5883 = n4059 & n5498;
  assign n5884 = ~n5845 & ~n5883;
  assign n5885 = n4057 & n5502;
  assign n5886 = ~n5850 & ~n5885;
  assign n5887 = n5884 & n5886;
  assign n5888 = ~n5834 & n5887;
  assign n5889 = n738 & ~n5888;
  assign n5890 = n4059 & n5531;
  assign n5891 = ~n5834 & ~n5890;
  assign n5892 = n4062 & n5521;
  assign n5893 = n4057 & n5528;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = n4065 & n5524;
  assign n5896 = n5894 & ~n5895;
  assign n5897 = n5891 & n5896;
  assign n5898 = ~n5857 & ~n5897;
  assign n5899 = n4089 & n5407;
  assign n5900 = ~n5868 & ~n5899;
  assign n5901 = ~n5898 & n5900;
  assign n5902 = ~n5889 & n5901;
  assign n5903 = ~n5882 & n5902;
  assign n5904 = n1178 & ~n5903;
  assign n5905 = n4053 & n5471;
  assign n5906 = ~n5541 & n5905;
  assign n5907 = n4057 & n5551;
  assign n5908 = n4065 & ~n5465;
  assign n5909 = ~n5059 & n5908;
  assign n5910 = n4059 & n5545;
  assign n5911 = n4062 & ~n5458;
  assign n5912 = ~n5050 & n5911;
  assign n5913 = ~n5910 & ~n5912;
  assign n5914 = ~n5909 & n5913;
  assign n5915 = ~n5834 & n5914;
  assign n5916 = ~n5907 & n5915;
  assign n5917 = n736 & ~n5916;
  assign n5918 = n4065 & n5561;
  assign n5919 = n4062 & ~n5436;
  assign n5920 = ~n5085 & n5919;
  assign n5921 = ~n5918 & ~n5920;
  assign n5922 = n4057 & n5557;
  assign n5923 = n4059 & ~n5441;
  assign n5924 = ~n5559 & n5923;
  assign n5925 = ~n5922 & ~n5924;
  assign n5926 = n5921 & n5925;
  assign n5927 = ~n5834 & n5926;
  assign n5928 = n738 & ~n5927;
  assign n5929 = n4059 & ~n5578;
  assign n5930 = n4057 & ~n5570;
  assign n5931 = ~n5834 & ~n5930;
  assign n5932 = n4062 & ~n5575;
  assign n5933 = n4065 & ~n5572;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = n5931 & n5934;
  assign n5936 = ~n5929 & n5935;
  assign n5937 = ~n5857 & ~n5936;
  assign n5938 = n4089 & n5451;
  assign n5939 = ~n5041 & n5938;
  assign n5940 = ~n5937 & ~n5939;
  assign n5941 = ~n5928 & n5940;
  assign n5942 = ~n5917 & n5941;
  assign n5943 = ~n5906 & n5942;
  assign n5944 = n1672 & ~n5943;
  assign n5945 = n4057 & n5454;
  assign n5946 = n4059 & n5461;
  assign n5947 = ~n5911 & ~n5946;
  assign n5948 = ~n5908 & n5947;
  assign n5949 = ~n5834 & n5948;
  assign n5950 = ~n5945 & n5949;
  assign n5951 = n736 & ~n5950;
  assign n5952 = ~n5919 & ~n5923;
  assign n5953 = n4057 & n5444;
  assign n5954 = n4065 & n5438;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = n5952 & n5955;
  assign n5957 = ~n5834 & n5956;
  assign n5958 = n738 & ~n5957;
  assign n5959 = n4059 & n5478;
  assign n5960 = n4057 & n5485;
  assign n5961 = ~n5834 & ~n5960;
  assign n5962 = n4065 & ~n5475;
  assign n5963 = n4062 & n5482;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = n5961 & n5964;
  assign n5966 = ~n5959 & n5965;
  assign n5967 = ~n5857 & ~n5966;
  assign n5968 = ~n5905 & ~n5967;
  assign n5969 = ~n5938 & n5968;
  assign n5970 = ~n5958 & n5969;
  assign n5971 = ~n5951 & n5970;
  assign n5972 = n1769 & ~n5971;
  assign n5973 = ~n5944 & ~n5972;
  assign n5974 = ~n5904 & n5973;
  assign n5975 = ~n5874 & n5974;
  assign n5976 = n680 & ~n5975;
  assign n5977 = n4193 & n5660;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = Ni10 & n5978;
  assign n5980 = ~n5831 & n5979;
  assign n5981 = n4437 & ~n5544;
  assign n5982 = n4429 & n5275;
  assign n5983 = ~n5001 & n5698;
  assign n5984 = ~n865 & ~n5983;
  assign n5985 = n4435 & ~n5550;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = ~n5982 & n5986;
  assign n5988 = ~n5981 & n5987;
  assign n5989 = n736 & ~n5988;
  assign n5990 = Pi19 & n5984;
  assign n5991 = ~n738 & ~n5990;
  assign n5992 = n4435 & ~n5556;
  assign n5993 = n4429 & ~n5253;
  assign n5994 = ~n5087 & n5360;
  assign n5995 = n4437 & ~n5994;
  assign n5996 = ~n5559 & n5995;
  assign n5997 = ~n5993 & ~n5996;
  assign n5998 = ~n5992 & n5997;
  assign n5999 = ~n5984 & n5998;
  assign n6000 = ~n5991 & ~n5999;
  assign n6001 = n4429 & n5280;
  assign n6002 = ~n5108 & n5360;
  assign n6003 = n4435 & ~n6002;
  assign n6004 = ~n5099 & n5360;
  assign n6005 = n4437 & ~n6004;
  assign n6006 = ~n5984 & ~n6005;
  assign n6007 = ~n6003 & n6006;
  assign n6008 = ~n6001 & n6007;
  assign n6009 = n923 & ~n6008;
  assign n6010 = n4459 & ~n5470;
  assign n6011 = ~n5541 & n6010;
  assign n6012 = ~Pi27 & n1031;
  assign n6013 = ~n5450 & n6012;
  assign n6014 = ~n5041 & n6013;
  assign n6015 = ~n6011 & ~n6014;
  assign n6016 = ~n6009 & n6015;
  assign n6017 = ~n6000 & n6016;
  assign n6018 = ~n5989 & n6017;
  assign n6019 = n1672 & ~n6018;
  assign n6020 = n4429 & ~n5215;
  assign n6021 = n4435 & ~n5443;
  assign n6022 = ~n5984 & ~n5995;
  assign n6023 = ~n6021 & n6022;
  assign n6024 = ~n6020 & n6023;
  assign n6025 = ~n5991 & ~n6024;
  assign n6026 = n4429 & n5224;
  assign n6027 = n4437 & ~n5460;
  assign n6028 = n4435 & ~n5453;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = ~n5984 & n6029;
  assign n6031 = ~n6026 & n6030;
  assign n6032 = n736 & ~n6031;
  assign n6033 = n4437 & ~n5477;
  assign n6034 = n4435 & ~n5484;
  assign n6035 = ~n6033 & ~n6034;
  assign n6036 = n4429 & n5237;
  assign n6037 = n6035 & ~n6036;
  assign n6038 = ~n5984 & n6037;
  assign n6039 = n923 & ~n6038;
  assign n6040 = ~n6032 & ~n6039;
  assign n6041 = ~n6010 & ~n6013;
  assign n6042 = n6040 & n6041;
  assign n6043 = ~n6025 & n6042;
  assign n6044 = n1769 & ~n6043;
  assign n6045 = ~n5207 & n6012;
  assign n6046 = ~n5012 & n5360;
  assign n6047 = n4435 & ~n6046;
  assign n6048 = n4429 & n5229;
  assign n6049 = ~n5032 & n5360;
  assign n6050 = n4437 & ~n6049;
  assign n6051 = ~n5984 & ~n6050;
  assign n6052 = ~n6048 & n6051;
  assign n6053 = ~n6047 & n6052;
  assign n6054 = n736 & ~n6053;
  assign n6055 = n4429 & n5220;
  assign n6056 = n4435 & ~n5501;
  assign n6057 = n4437 & ~n5497;
  assign n6058 = ~n5984 & ~n6057;
  assign n6059 = ~n6056 & n6058;
  assign n6060 = ~n6055 & n6059;
  assign n6061 = ~n5991 & ~n6060;
  assign n6062 = n4459 & ~n5426;
  assign n6063 = n4435 & ~n5527;
  assign n6064 = n4437 & ~n5530;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = n4429 & n5233;
  assign n6067 = n6065 & ~n6066;
  assign n6068 = ~n5984 & n6067;
  assign n6069 = n923 & ~n6068;
  assign n6070 = ~n6062 & ~n6069;
  assign n6071 = ~n6061 & n6070;
  assign n6072 = ~n6054 & n6071;
  assign n6073 = ~n6045 & n6072;
  assign n6074 = n1178 & ~n6073;
  assign n6075 = ~n6044 & ~n6074;
  assign n6076 = ~n6019 & n6075;
  assign n6077 = ~n5013 & n5360;
  assign n6078 = n4435 & ~n6077;
  assign n6079 = n4429 & n5258;
  assign n6080 = n4437 & ~n5390;
  assign n6081 = ~n5984 & ~n6080;
  assign n6082 = ~n6079 & n6081;
  assign n6083 = ~n6078 & n6082;
  assign n6084 = n736 & ~n6083;
  assign n6085 = n4429 & n5269;
  assign n6086 = n4435 & ~n5361;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = n4437 & ~n5366;
  assign n6089 = ~n5984 & ~n6088;
  assign n6090 = n6087 & n6089;
  assign n6091 = ~n5991 & ~n6090;
  assign n6092 = n4429 & n5262;
  assign n6093 = ~n5137 & n5360;
  assign n6094 = n4435 & ~n6093;
  assign n6095 = ~n5143 & n5360;
  assign n6096 = n4437 & ~n6095;
  assign n6097 = ~n5984 & ~n6096;
  assign n6098 = ~n6094 & n6097;
  assign n6099 = ~n6092 & n6098;
  assign n6100 = n923 & ~n6099;
  assign n6101 = ~n6091 & ~n6100;
  assign n6102 = ~n5425 & n6062;
  assign n6103 = ~n5018 & n6045;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = n6101 & n6104;
  assign n6106 = ~n6084 & n6105;
  assign n6107 = n1610 & ~n6106;
  assign n6108 = Ni14 & ~n6107;
  assign n6109 = n6076 & n6108;
  assign n6110 = n4321 & ~n5253;
  assign n6111 = ~n5001 & n5373;
  assign n6112 = ~n865 & ~n6111;
  assign n6113 = n4324 & ~n5994;
  assign n6114 = ~n5559 & n6113;
  assign n6115 = ~n6112 & ~n6114;
  assign n6116 = ~n6110 & n6115;
  assign n6117 = n738 & ~n6116;
  assign n6118 = n4321 & n5275;
  assign n6119 = n4329 & ~n5550;
  assign n6120 = n4324 & ~n5544;
  assign n6121 = ~n6112 & ~n6120;
  assign n6122 = ~n6119 & n6121;
  assign n6123 = ~n6118 & n6122;
  assign n6124 = n736 & ~n6123;
  assign n6125 = n4350 & ~n5556;
  assign n6126 = ~n604 & n1031;
  assign n6127 = ~n5450 & n6126;
  assign n6128 = ~n5041 & n6127;
  assign n6129 = n923 & n4321;
  assign n6130 = n5280 & n6129;
  assign n6131 = ~n6128 & ~n6130;
  assign n6132 = ~n6125 & n6131;
  assign n6133 = ~n6124 & n6132;
  assign n6134 = n730 & n6112;
  assign n6135 = ~n923 & ~n6134;
  assign n6136 = n4329 & ~n6002;
  assign n6137 = n4324 & ~n6004;
  assign n6138 = ~n6112 & ~n6137;
  assign n6139 = ~n6136 & n6138;
  assign n6140 = ~n6135 & ~n6139;
  assign n6141 = n4359 & ~n5470;
  assign n6142 = ~n5541 & n6141;
  assign n6143 = ~n6140 & ~n6142;
  assign n6144 = n6133 & n6143;
  assign n6145 = ~n6117 & n6144;
  assign n6146 = n1672 & ~n6145;
  assign n6147 = n4321 & n5269;
  assign n6148 = n4324 & ~n5366;
  assign n6149 = ~n6112 & ~n6148;
  assign n6150 = ~n6147 & n6149;
  assign n6151 = n738 & ~n6150;
  assign n6152 = n4321 & n5258;
  assign n6153 = n4329 & ~n6077;
  assign n6154 = n4324 & ~n5390;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6112 & n6155;
  assign n6157 = ~n6152 & n6156;
  assign n6158 = n736 & ~n6157;
  assign n6159 = n4350 & ~n5361;
  assign n6160 = ~n5207 & n6126;
  assign n6161 = ~n5018 & n6160;
  assign n6162 = n4359 & ~n5426;
  assign n6163 = ~n5425 & n6162;
  assign n6164 = ~n6161 & ~n6163;
  assign n6165 = ~n6159 & n6164;
  assign n6166 = n4321 & n5262;
  assign n6167 = n4324 & ~n6095;
  assign n6168 = ~n6166 & ~n6167;
  assign n6169 = n4329 & ~n6093;
  assign n6170 = ~n6112 & ~n6169;
  assign n6171 = n6168 & n6170;
  assign n6172 = ~n6135 & ~n6171;
  assign n6173 = n6165 & ~n6172;
  assign n6174 = ~n6158 & n6173;
  assign n6175 = ~n6151 & n6174;
  assign n6176 = n1610 & ~n6175;
  assign n6177 = n4321 & ~n5215;
  assign n6178 = ~n6113 & ~n6177;
  assign n6179 = n738 & ~n6178;
  assign n6180 = n4329 & ~n5484;
  assign n6181 = n4324 & ~n5477;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = n923 & ~n6182;
  assign n6184 = ~n6127 & ~n6183;
  assign n6185 = n4350 & ~n5443;
  assign n6186 = n6184 & ~n6185;
  assign n6187 = n4321 & n5224;
  assign n6188 = n4329 & ~n5453;
  assign n6189 = n4324 & ~n5460;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~n6187 & n6190;
  assign n6192 = n736 & ~n6191;
  assign n6193 = n5237 & n6129;
  assign n6194 = ~n6112 & ~n6193;
  assign n6195 = ~n6141 & n6194;
  assign n6196 = ~n6192 & n6195;
  assign n6197 = n6186 & n6196;
  assign n6198 = ~n6179 & n6197;
  assign n6199 = n1769 & ~n6198;
  assign n6200 = n4324 & ~n5530;
  assign n6201 = n4329 & ~n5527;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = n923 & ~n6202;
  assign n6204 = n4321 & n5229;
  assign n6205 = n4329 & ~n6046;
  assign n6206 = n4324 & ~n6049;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = ~n6204 & n6207;
  assign n6209 = n736 & ~n6208;
  assign n6210 = n4321 & n5220;
  assign n6211 = n4329 & ~n5501;
  assign n6212 = n4324 & ~n5497;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = ~n6210 & n6213;
  assign n6215 = n738 & ~n6214;
  assign n6216 = ~n6112 & ~n6160;
  assign n6217 = ~n6162 & n6216;
  assign n6218 = n5233 & n6129;
  assign n6219 = n6217 & ~n6218;
  assign n6220 = ~n6215 & n6219;
  assign n6221 = ~n6209 & n6220;
  assign n6222 = ~n6203 & n6221;
  assign n6223 = n1178 & ~n6222;
  assign n6224 = ~n6199 & ~n6223;
  assign n6225 = ~n6176 & n6224;
  assign n6226 = ~n6146 & n6225;
  assign n6227 = ~Ni14 & n6226;
  assign n6228 = n671 & ~n6227;
  assign n6229 = ~n6109 & n6228;
  assign n6230 = n4522 & ~n5443;
  assign n6231 = n4520 & ~n5994;
  assign n6232 = n4514 & ~n5215;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = ~n6230 & n6233;
  assign n6235 = n738 & ~n6234;
  assign n6236 = n736 & n4514;
  assign n6237 = n5224 & n6236;
  assign n6238 = n4520 & ~n5460;
  assign n6239 = ~n5001 & n5833;
  assign n6240 = ~n865 & ~n6239;
  assign n6241 = n4522 & ~n5453;
  assign n6242 = ~n6240 & ~n6241;
  assign n6243 = ~n6238 & n6242;
  assign n6244 = n736 & ~n6243;
  assign n6245 = n4514 & n5237;
  assign n6246 = n4522 & ~n5484;
  assign n6247 = n4520 & ~n5477;
  assign n6248 = ~n6240 & ~n6247;
  assign n6249 = ~n6246 & n6248;
  assign n6250 = ~n6245 & n6249;
  assign n6251 = n923 & ~n6250;
  assign n6252 = n4535 & ~n5470;
  assign n6253 = n4516 & ~n5450;
  assign n6254 = Pi19 & n6240;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6252 & n6255;
  assign n6257 = ~n6251 & n6256;
  assign n6258 = ~n6244 & n6257;
  assign n6259 = ~n6237 & n6258;
  assign n6260 = ~n6235 & n6259;
  assign n6261 = n1769 & ~n6260;
  assign n6262 = n4514 & ~n5253;
  assign n6263 = n4522 & ~n5556;
  assign n6264 = ~n5559 & n6231;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = ~n6262 & n6265;
  assign n6267 = n738 & ~n6266;
  assign n6268 = n4522 & ~n6002;
  assign n6269 = n4520 & ~n6004;
  assign n6270 = n4514 & n5280;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = ~n6268 & n6271;
  assign n6273 = n923 & ~n6272;
  assign n6274 = ~n5541 & n6252;
  assign n6275 = ~n6240 & ~n6274;
  assign n6276 = ~n6273 & n6275;
  assign n6277 = ~n5041 & n6253;
  assign n6278 = n4522 & ~n5550;
  assign n6279 = n4520 & ~n5544;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = n736 & ~n6280;
  assign n6282 = n5275 & n6236;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~n6277 & n6283;
  assign n6285 = n6276 & n6284;
  assign n6286 = ~n6267 & n6285;
  assign n6287 = n1672 & ~n6286;
  assign n6288 = n4514 & n5220;
  assign n6289 = n4522 & ~n5501;
  assign n6290 = n4520 & ~n5497;
  assign n6291 = Pi19 & ~n6290;
  assign n6292 = ~n6289 & n6291;
  assign n6293 = ~n6288 & n6292;
  assign n6294 = n4514 & n5233;
  assign n6295 = n4520 & ~n5530;
  assign n6296 = n4522 & ~n5527;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = n923 & n6297;
  assign n6299 = ~n6294 & n6298;
  assign n6300 = ~n6293 & ~n6299;
  assign n6301 = n4514 & n5229;
  assign n6302 = n4522 & ~n6046;
  assign n6303 = n4520 & ~n6049;
  assign n6304 = ~n6302 & ~n6303;
  assign n6305 = ~n6301 & n6304;
  assign n6306 = ~Pi19 & ~n6305;
  assign n6307 = Pi17 & ~n6306;
  assign n6308 = n6300 & ~n6307;
  assign n6309 = n4516 & ~n5207;
  assign n6310 = n4535 & ~n5426;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n6308 & n6311;
  assign n6313 = ~n6240 & n6312;
  assign n6314 = n1178 & ~n6313;
  assign n6315 = n4520 & ~n5390;
  assign n6316 = n4522 & ~n6077;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~n6240 & n6317;
  assign n6319 = n736 & ~n6318;
  assign n6320 = n4520 & ~n5366;
  assign n6321 = n4522 & ~n5361;
  assign n6322 = ~n6240 & ~n6321;
  assign n6323 = ~n6320 & n6322;
  assign n6324 = n738 & ~n6323;
  assign n6325 = n4545 & n5269;
  assign n6326 = Pi17 & n6254;
  assign n6327 = ~n6325 & ~n6326;
  assign n6328 = ~n6324 & n6327;
  assign n6329 = n4522 & ~n6093;
  assign n6330 = n4514 & n5262;
  assign n6331 = n4520 & ~n6095;
  assign n6332 = ~n6240 & ~n6331;
  assign n6333 = ~n6330 & n6332;
  assign n6334 = ~n6329 & n6333;
  assign n6335 = n923 & ~n6334;
  assign n6336 = n5258 & n6236;
  assign n6337 = n4516 & n5247;
  assign n6338 = ~n5425 & n6310;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = ~n6336 & n6339;
  assign n6341 = ~n6335 & n6340;
  assign n6342 = n6328 & n6341;
  assign n6343 = ~n6319 & n6342;
  assign n6344 = n1610 & ~n6343;
  assign n6345 = ~n6314 & ~n6344;
  assign n6346 = ~n6287 & n6345;
  assign n6347 = ~n6261 & n6346;
  assign n6348 = n680 & ~n6347;
  assign n6349 = ~Ni10 & n5289;
  assign n6350 = ~n4227 & ~n6349;
  assign n6351 = ~n6348 & ~n6350;
  assign n6352 = ~n6229 & n6351;
  assign n6353 = ~n5980 & ~n6352;
  assign n6354 = ~n5359 & ~n6353;
  assign n6355 = n579 & ~n6354;
  assign n6356 = n680 & ~n6239;
  assign n6357 = ~n4226 & ~n5002;
  assign n6358 = ~Ni14 & ~n6111;
  assign n6359 = n4427 & n6358;
  assign n6360 = n4046 & ~n5983;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n6357 & n6361;
  assign n6363 = Ni11 & n5002;
  assign n6364 = ~n6362 & ~n6363;
  assign n6365 = ~n680 & n6364;
  assign n6366 = ~n6356 & ~n6365;
  assign n6367 = ~n5202 & n6366;
  assign n6368 = n4592 & ~n6367;
  assign n6369 = ~Pi27 & n854;
  assign n6370 = ~n652 & ~n6369;
  assign n6371 = Ni14 & ~n6370;
  assign n6372 = Ni14 & ~n5698;
  assign n6373 = ~n6358 & ~n6372;
  assign n6374 = ~Pi24 & ~n6373;
  assign n6375 = ~n652 & ~n854;
  assign n6376 = n604 & ~n652;
  assign n6377 = ~n6375 & ~n6376;
  assign n6378 = ~Ni14 & n6377;
  assign n6379 = ~n5001 & ~n6378;
  assign n6380 = ~n6374 & n6379;
  assign n6381 = ~n6371 & n6380;
  assign n6382 = n671 & ~n6381;
  assign n6383 = n4691 & ~n5089;
  assign n6384 = ~n5184 & n6375;
  assign n6385 = n4695 & ~n6384;
  assign n6386 = n4699 & ~n5185;
  assign n6387 = ~n5088 & n6375;
  assign n6388 = n4693 & ~n6387;
  assign n6389 = ~n6386 & ~n6388;
  assign n6390 = ~n6385 & n6389;
  assign n6391 = ~n6383 & n6390;
  assign n6392 = n955 & ~n6391;
  assign n6393 = ~Pi24 & ~n5345;
  assign n6394 = n4699 & ~n5170;
  assign n6395 = ~n5164 & n6375;
  assign n6396 = n4693 & ~n6395;
  assign n6397 = n4691 & ~n5165;
  assign n6398 = ~n5169 & n6375;
  assign n6399 = n4695 & ~n6398;
  assign n6400 = ~n6397 & ~n6399;
  assign n6401 = ~n6396 & n6400;
  assign n6402 = ~n6394 & n6401;
  assign n6403 = n994 & ~n6402;
  assign n6404 = ~n6393 & ~n6403;
  assign n6405 = ~n6392 & n6404;
  assign n6406 = ~n5309 & ~n5314;
  assign n6407 = n4699 & ~n6406;
  assign n6408 = ~n5153 & n6375;
  assign n6409 = n4693 & ~n6408;
  assign n6410 = n4691 & ~n5154;
  assign n6411 = ~n5129 & n6375;
  assign n6412 = n4695 & ~n6411;
  assign n6413 = ~n6410 & ~n6412;
  assign n6414 = ~n6409 & n6413;
  assign n6415 = n903 & ~n6414;
  assign n6416 = n4691 & ~n5182;
  assign n6417 = ~n5181 & n6375;
  assign n6418 = n4693 & ~n6417;
  assign n6419 = n4699 & ~n5190;
  assign n6420 = ~n5189 & n6375;
  assign n6421 = n4695 & ~n6420;
  assign n6422 = ~n6419 & ~n6421;
  assign n6423 = ~n6418 & n6422;
  assign n6424 = ~n6416 & n6423;
  assign n6425 = n924 & ~n6424;
  assign n6426 = ~n6415 & ~n6425;
  assign n6427 = ~n6407 & n6426;
  assign n6428 = ~n5053 & n6375;
  assign n6429 = n4693 & ~n6428;
  assign n6430 = n4691 & ~n5054;
  assign n6431 = ~n5062 & n6375;
  assign n6432 = n4695 & ~n6431;
  assign n6433 = ~n6430 & ~n6432;
  assign n6434 = ~n6429 & n6433;
  assign n6435 = n1035 & ~n6434;
  assign n6436 = ~n5033 & n6375;
  assign n6437 = n4693 & ~n6436;
  assign n6438 = ~n5072 & n6375;
  assign n6439 = n4695 & ~n6438;
  assign n6440 = n4699 & ~n5073;
  assign n6441 = n4691 & ~n5034;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n6439 & n6442;
  assign n6444 = ~n6437 & n6443;
  assign n6445 = n869 & ~n6444;
  assign n6446 = ~n864 & ~n6375;
  assign n6447 = ~Pi24 & n5019;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n5023 & n6375;
  assign n6450 = n4684 & ~n6449;
  assign n6451 = ~n5044 & n6375;
  assign n6452 = n4683 & ~n6451;
  assign n6453 = ~n6450 & ~n6452;
  assign n6454 = n6448 & n6453;
  assign n6455 = ~n6445 & n6454;
  assign n6456 = ~n6435 & n6455;
  assign n6457 = n6427 & n6456;
  assign n6458 = n6405 & n6457;
  assign n6459 = n1381 & ~n6458;
  assign n6460 = ~n678 & ~n4427;
  assign n6461 = n871 & n5000;
  assign n6462 = ~Ni12 & n5833;
  assign n6463 = ~n6461 & n6462;
  assign n6464 = Ni11 & ~n6463;
  assign n6465 = ~n6460 & ~n6464;
  assign n6466 = n6375 & ~n6461;
  assign n6467 = n864 & ~n6466;
  assign n6468 = Ni30 & n864;
  assign n6469 = ~n5001 & ~n6468;
  assign n6470 = ~Pi24 & ~n6469;
  assign n6471 = n6448 & ~n6470;
  assign n6472 = ~n6467 & n6471;
  assign n6473 = ~n6465 & ~n6472;
  assign n6474 = n4699 & ~n5139;
  assign n6475 = ~n5138 & n6375;
  assign n6476 = n4695 & ~n6475;
  assign n6477 = n4691 & ~n5145;
  assign n6478 = ~n5144 & n6375;
  assign n6479 = n4693 & ~n6478;
  assign n6480 = ~n6477 & ~n6479;
  assign n6481 = ~n6476 & n6480;
  assign n6482 = ~n6474 & n6481;
  assign n6483 = n994 & ~n6482;
  assign n6484 = ~n5030 & n6441;
  assign n6485 = ~n5014 & n6375;
  assign n6486 = n4695 & ~n6485;
  assign n6487 = n5029 & n6375;
  assign n6488 = n6437 & ~n6487;
  assign n6489 = ~n6486 & ~n6488;
  assign n6490 = ~n6484 & n6489;
  assign n6491 = n869 & ~n6490;
  assign n6492 = ~Pi24 & ~n5305;
  assign n6493 = n5040 & n6375;
  assign n6494 = n6452 & ~n6493;
  assign n6495 = ~n6492 & ~n6494;
  assign n6496 = n6448 & n6495;
  assign n6497 = ~n6491 & n6496;
  assign n6498 = ~n6483 & n6497;
  assign n6499 = n4699 & ~n5319;
  assign n6500 = n5017 & n6375;
  assign n6501 = n6450 & ~n6500;
  assign n6502 = n4691 & ~n5101;
  assign n6503 = ~n5109 & n6375;
  assign n6504 = n4695 & ~n6503;
  assign n6505 = ~n5100 & n6375;
  assign n6506 = n4693 & ~n6505;
  assign n6507 = ~n6504 & ~n6506;
  assign n6508 = ~n6502 & n6507;
  assign n6509 = n924 & ~n6508;
  assign n6510 = ~n6501 & ~n6509;
  assign n6511 = ~n6499 & n6510;
  assign n6512 = ~n5050 & n6430;
  assign n6513 = n5049 & n6375;
  assign n6514 = n6429 & ~n6513;
  assign n6515 = n5058 & n6375;
  assign n6516 = n6432 & ~n6515;
  assign n6517 = ~n6514 & ~n6516;
  assign n6518 = ~n6512 & n6517;
  assign n6519 = n1035 & ~n6518;
  assign n6520 = n5149 & n6375;
  assign n6521 = n6409 & ~n6520;
  assign n6522 = n4691 & n5155;
  assign n6523 = n5131 & n6375;
  assign n6524 = n6412 & ~n6523;
  assign n6525 = ~n6522 & ~n6524;
  assign n6526 = ~n6521 & n6525;
  assign n6527 = n903 & ~n6526;
  assign n6528 = ~n6519 & ~n6527;
  assign n6529 = ~n5119 & n6375;
  assign n6530 = n4695 & ~n6529;
  assign n6531 = n5084 & n6375;
  assign n6532 = n6388 & ~n6531;
  assign n6533 = ~n5085 & n6383;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = ~n6530 & n6534;
  assign n6536 = n955 & ~n6535;
  assign n6537 = n6528 & ~n6536;
  assign n6538 = n6511 & n6537;
  assign n6539 = n6498 & n6538;
  assign n6540 = n1190 & ~n6539;
  assign n6541 = ~n6473 & ~n6540;
  assign n6542 = ~n6459 & n6541;
  assign n6543 = ~n6382 & n6542;
  assign n6544 = n4682 & ~n6543;
  assign n6545 = n3208 & ~n5024;
  assign n6546 = ~n5018 & n6545;
  assign n6547 = n3257 & ~n5139;
  assign n6548 = n691 & n6375;
  assign n6549 = n5019 & ~n6548;
  assign n6550 = n3232 & ~n6475;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = n3248 & ~n6478;
  assign n6553 = n3263 & ~n5145;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n6551 & n6554;
  assign n6556 = ~n6547 & n6555;
  assign n6557 = n923 & ~n6556;
  assign n6558 = n730 & n6549;
  assign n6559 = ~n736 & ~n6558;
  assign n6560 = n3263 & ~n5034;
  assign n6561 = ~n6549 & ~n6560;
  assign n6562 = ~n5030 & ~n6561;
  assign n6563 = n3232 & ~n6485;
  assign n6564 = n3248 & ~n6436;
  assign n6565 = ~n6487 & n6564;
  assign n6566 = ~n6563 & ~n6565;
  assign n6567 = n3257 & ~n5015;
  assign n6568 = n6566 & ~n6567;
  assign n6569 = ~n6562 & n6568;
  assign n6570 = ~n6559 & ~n6569;
  assign n6571 = ~n6557 & ~n6570;
  assign n6572 = n3345 & ~n6449;
  assign n6573 = ~n6500 & n6572;
  assign n6574 = n3248 & ~n6408;
  assign n6575 = ~n6520 & n6574;
  assign n6576 = n3257 & ~n5130;
  assign n6577 = ~n6549 & ~n6576;
  assign n6578 = ~n5132 & ~n6577;
  assign n6579 = n3263 & n5155;
  assign n6580 = n3232 & ~n6411;
  assign n6581 = ~n6523 & n6580;
  assign n6582 = ~n6579 & ~n6581;
  assign n6583 = ~n6578 & n6582;
  assign n6584 = ~n6575 & n6583;
  assign n6585 = n738 & ~n6584;
  assign n6586 = ~n6573 & ~n6585;
  assign n6587 = n6571 & n6586;
  assign n6588 = ~n6546 & n6587;
  assign n6589 = n1610 & ~n6588;
  assign n6590 = n3232 & ~n6438;
  assign n6591 = n3257 & ~n5073;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = n6561 & n6592;
  assign n6594 = ~n6564 & n6593;
  assign n6595 = n736 & ~n6594;
  assign n6596 = ~n923 & ~n6558;
  assign n6597 = n3248 & ~n6395;
  assign n6598 = n3257 & ~n5170;
  assign n6599 = n3232 & ~n6398;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = n3263 & ~n5165;
  assign n6602 = n6600 & ~n6601;
  assign n6603 = ~n6597 & n6602;
  assign n6604 = ~n6549 & n6603;
  assign n6605 = ~n6596 & ~n6604;
  assign n6606 = ~n6545 & ~n6605;
  assign n6607 = n3263 & ~n5154;
  assign n6608 = ~n6574 & ~n6580;
  assign n6609 = n6577 & n6608;
  assign n6610 = ~n6607 & n6609;
  assign n6611 = n738 & ~n6610;
  assign n6612 = ~n6572 & ~n6611;
  assign n6613 = n6606 & n6612;
  assign n6614 = ~n6595 & n6613;
  assign n6615 = n1178 & ~n6614;
  assign n6616 = n3208 & ~n5045;
  assign n6617 = ~n5041 & n6616;
  assign n6618 = n3257 & ~n5120;
  assign n6619 = n3232 & ~n6529;
  assign n6620 = n3248 & ~n6387;
  assign n6621 = ~n6531 & n6620;
  assign n6622 = ~n6619 & ~n6621;
  assign n6623 = n3263 & ~n5089;
  assign n6624 = ~n6549 & ~n6623;
  assign n6625 = ~n5085 & ~n6624;
  assign n6626 = n6622 & ~n6625;
  assign n6627 = ~n6618 & n6626;
  assign n6628 = n738 & ~n6627;
  assign n6629 = n3248 & ~n6428;
  assign n6630 = ~n6513 & n6629;
  assign n6631 = n3263 & ~n5054;
  assign n6632 = ~n6549 & ~n6631;
  assign n6633 = ~n5050 & ~n6632;
  assign n6634 = n3257 & ~n5063;
  assign n6635 = ~n5059 & n6634;
  assign n6636 = n3232 & ~n6431;
  assign n6637 = ~n6515 & n6636;
  assign n6638 = ~n6635 & ~n6637;
  assign n6639 = ~n6633 & n6638;
  assign n6640 = ~n6630 & n6639;
  assign n6641 = n736 & ~n6640;
  assign n6642 = n3263 & ~n5101;
  assign n6643 = n3257 & ~n5110;
  assign n6644 = n3248 & ~n6505;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = n3232 & ~n6503;
  assign n6647 = n6645 & ~n6646;
  assign n6648 = ~n6642 & n6647;
  assign n6649 = ~n6549 & n6648;
  assign n6650 = ~n6596 & ~n6649;
  assign n6651 = n3345 & ~n6451;
  assign n6652 = ~n6493 & n6651;
  assign n6653 = ~n6650 & ~n6652;
  assign n6654 = ~n6641 & n6653;
  assign n6655 = ~n6628 & n6654;
  assign n6656 = ~n6617 & n6655;
  assign n6657 = n1672 & ~n6656;
  assign n6658 = ~n6629 & ~n6636;
  assign n6659 = n6632 & n6658;
  assign n6660 = ~n6634 & n6659;
  assign n6661 = n736 & ~n6660;
  assign n6662 = n3257 & ~n5185;
  assign n6663 = n3232 & ~n6384;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = ~n6620 & n6664;
  assign n6666 = n6624 & n6665;
  assign n6667 = n738 & ~n6666;
  assign n6668 = n3263 & ~n5182;
  assign n6669 = n3257 & ~n5190;
  assign n6670 = ~n6549 & ~n6669;
  assign n6671 = n3248 & ~n6417;
  assign n6672 = n3232 & ~n6420;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = n6670 & n6673;
  assign n6675 = ~n6668 & n6674;
  assign n6676 = ~n6596 & ~n6675;
  assign n6677 = ~n6616 & ~n6676;
  assign n6678 = ~n6667 & n6677;
  assign n6679 = ~n6651 & n6678;
  assign n6680 = ~n6661 & n6679;
  assign n6681 = n1769 & ~n6680;
  assign n6682 = ~n6657 & ~n6681;
  assign n6683 = ~n6615 & n6682;
  assign n6684 = ~n6589 & n6683;
  assign n6685 = n570 & ~n6684;
  assign n6686 = ~n691 & ~n6469;
  assign n6687 = ~n6549 & ~n6686;
  assign n6688 = ~n6467 & n6687;
  assign n6689 = n3087 & ~n6688;
  assign n6690 = Ni14 & n864;
  assign n6691 = ~n5983 & n6690;
  assign n6692 = ~Ni14 & ~n5373;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = ~n691 & ~n6693;
  assign n6695 = ~Ni14 & ~n864;
  assign n6696 = ~n5699 & ~n6358;
  assign n6697 = ~n6695 & ~n6696;
  assign n6698 = ~Pi23 & n6697;
  assign n6699 = ~Pi24 & n6370;
  assign n6700 = n6372 & ~n6699;
  assign n6701 = ~n6111 & ~n6379;
  assign n6702 = ~n6700 & ~n6701;
  assign n6703 = ~n6698 & n6702;
  assign n6704 = ~n6694 & n6703;
  assign n6705 = n670 & ~n6704;
  assign n6706 = ~n5001 & n6548;
  assign n6707 = n6356 & ~n6706;
  assign n6708 = ~n6705 & ~n6707;
  assign n6709 = ~n6689 & n6708;
  assign n6710 = ~n6685 & n6709;
  assign n6711 = n694 & ~n6710;
  assign n6712 = ~n6544 & ~n6711;
  assign n6713 = n637 & n6375;
  assign n6714 = n5019 & ~n6713;
  assign n6715 = n730 & n6714;
  assign n6716 = ~n923 & ~n6715;
  assign n6717 = n4846 & ~n5165;
  assign n6718 = n4839 & ~n6398;
  assign n6719 = n4833 & ~n5170;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = n4841 & ~n6395;
  assign n6722 = n6720 & ~n6721;
  assign n6723 = ~n6717 & n6722;
  assign n6724 = ~n6714 & n6723;
  assign n6725 = ~n6716 & ~n6724;
  assign n6726 = n4877 & ~n5024;
  assign n6727 = n4839 & ~n6411;
  assign n6728 = n4833 & ~n5130;
  assign n6729 = ~n6714 & ~n6728;
  assign n6730 = n4841 & ~n6408;
  assign n6731 = n4846 & ~n5154;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = n6729 & n6732;
  assign n6734 = ~n6727 & n6733;
  assign n6735 = n738 & ~n6734;
  assign n6736 = n4861 & ~n6449;
  assign n6737 = n4839 & ~n6438;
  assign n6738 = n4846 & ~n5034;
  assign n6739 = ~n6714 & ~n6738;
  assign n6740 = n4841 & ~n6436;
  assign n6741 = n4833 & ~n5073;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = n6739 & n6742;
  assign n6744 = ~n6737 & n6743;
  assign n6745 = n736 & ~n6744;
  assign n6746 = ~n6736 & ~n6745;
  assign n6747 = ~n6735 & n6746;
  assign n6748 = ~n6726 & n6747;
  assign n6749 = ~n6725 & n6748;
  assign n6750 = n1178 & ~n6749;
  assign n6751 = ~n736 & ~n6715;
  assign n6752 = n4846 & ~n5054;
  assign n6753 = ~n6714 & ~n6752;
  assign n6754 = n4839 & ~n6431;
  assign n6755 = n4841 & ~n6428;
  assign n6756 = ~n6754 & ~n6755;
  assign n6757 = n4833 & ~n5063;
  assign n6758 = n6756 & ~n6757;
  assign n6759 = n6753 & n6758;
  assign n6760 = ~n6751 & ~n6759;
  assign n6761 = n4846 & ~n5089;
  assign n6762 = ~n6714 & ~n6761;
  assign n6763 = n4839 & ~n6384;
  assign n6764 = n6762 & ~n6763;
  assign n6765 = n4841 & ~n6387;
  assign n6766 = n4833 & ~n5185;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = n6764 & n6767;
  assign n6769 = n738 & ~n6768;
  assign n6770 = n4877 & ~n5045;
  assign n6771 = n4861 & ~n6451;
  assign n6772 = n4846 & ~n5182;
  assign n6773 = n4833 & ~n5190;
  assign n6774 = n4841 & ~n6417;
  assign n6775 = ~n6773 & ~n6774;
  assign n6776 = n4839 & ~n6420;
  assign n6777 = ~n6714 & ~n6776;
  assign n6778 = n6775 & n6777;
  assign n6779 = ~n6772 & n6778;
  assign n6780 = n923 & ~n6779;
  assign n6781 = ~n6771 & ~n6780;
  assign n6782 = ~n6770 & n6781;
  assign n6783 = ~n6769 & n6782;
  assign n6784 = ~n6760 & n6783;
  assign n6785 = n1769 & ~n6784;
  assign n6786 = ~n5018 & n6726;
  assign n6787 = n4839 & ~n6485;
  assign n6788 = ~n5030 & ~n6739;
  assign n6789 = ~n6487 & n6740;
  assign n6790 = n4833 & ~n5015;
  assign n6791 = ~n6789 & ~n6790;
  assign n6792 = ~n6788 & n6791;
  assign n6793 = ~n6787 & n6792;
  assign n6794 = n736 & ~n6793;
  assign n6795 = ~n6520 & n6730;
  assign n6796 = n4846 & n5155;
  assign n6797 = ~n6795 & ~n6796;
  assign n6798 = ~n6523 & n6727;
  assign n6799 = n4833 & n5133;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = n6797 & n6800;
  assign n6802 = ~n6714 & n6801;
  assign n6803 = n738 & ~n6802;
  assign n6804 = n4846 & ~n5145;
  assign n6805 = n4833 & ~n5139;
  assign n6806 = n4839 & ~n6475;
  assign n6807 = ~n6714 & ~n6806;
  assign n6808 = n4841 & ~n6478;
  assign n6809 = n6807 & ~n6808;
  assign n6810 = ~n6805 & n6809;
  assign n6811 = ~n6804 & n6810;
  assign n6812 = ~n6716 & ~n6811;
  assign n6813 = ~n6500 & n6736;
  assign n6814 = ~n6812 & ~n6813;
  assign n6815 = ~n6803 & n6814;
  assign n6816 = ~n6794 & n6815;
  assign n6817 = ~n6786 & n6816;
  assign n6818 = n1610 & ~n6817;
  assign n6819 = ~n6493 & n6771;
  assign n6820 = ~n6513 & n6755;
  assign n6821 = ~n5050 & ~n6753;
  assign n6822 = ~n5059 & n6757;
  assign n6823 = ~n6515 & n6754;
  assign n6824 = ~n6822 & ~n6823;
  assign n6825 = ~n6821 & n6824;
  assign n6826 = ~n6820 & n6825;
  assign n6827 = n736 & ~n6826;
  assign n6828 = ~n6531 & n6765;
  assign n6829 = ~n5085 & ~n6762;
  assign n6830 = n4839 & ~n6529;
  assign n6831 = n4833 & ~n5120;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = ~n6829 & n6832;
  assign n6834 = ~n6828 & n6833;
  assign n6835 = n738 & ~n6834;
  assign n6836 = n4846 & ~n5101;
  assign n6837 = n4833 & ~n5110;
  assign n6838 = ~n6714 & ~n6837;
  assign n6839 = n4839 & ~n6503;
  assign n6840 = n4841 & ~n6505;
  assign n6841 = ~n6839 & ~n6840;
  assign n6842 = n6838 & n6841;
  assign n6843 = ~n6836 & n6842;
  assign n6844 = ~n6716 & ~n6843;
  assign n6845 = ~n5041 & n6770;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n6835 & n6846;
  assign n6848 = ~n6827 & n6847;
  assign n6849 = ~n6819 & n6848;
  assign n6850 = n1672 & ~n6849;
  assign n6851 = ~n6818 & ~n6850;
  assign n6852 = ~n6785 & n6851;
  assign n6853 = ~n6750 & n6852;
  assign n6854 = n570 & ~n6853;
  assign n6855 = ~n637 & ~n6469;
  assign n6856 = ~n6714 & ~n6855;
  assign n6857 = ~n6467 & n6856;
  assign n6858 = n3087 & ~n6857;
  assign n6859 = ~n637 & ~n6693;
  assign n6860 = Pi23 & n6697;
  assign n6861 = n6702 & ~n6860;
  assign n6862 = ~n6859 & n6861;
  assign n6863 = n670 & ~n6862;
  assign n6864 = ~n5001 & n6713;
  assign n6865 = n6356 & ~n6864;
  assign n6866 = ~n6863 & ~n6865;
  assign n6867 = ~n6858 & n6866;
  assign n6868 = ~n6854 & n6867;
  assign n6869 = n4819 & ~n6868;
  assign n6870 = n6712 & ~n6869;
  assign n6871 = ~n6368 & n6870;
  assign n6872 = ~n6355 & n6871;
  assign n6873 = n3086 & ~n6872;
  assign n6874 = ~n5205 & ~n6873;
  assign n6875 = Ni30 & ~P__cmxcl_1;
  assign n6876 = n4984 & ~n5697;
  assign n6877 = Ni10 & ~n5660;
  assign n6878 = ~n582 & ~n6877;
  assign n6879 = ~n6349 & n6878;
  assign n6880 = ~n6876 & ~n6879;
  assign n6881 = ~n5359 & n6880;
  assign n6882 = n4981 & ~n6881;
  assign n6883 = ~n6875 & ~n6882;
  assign n1022_1 = ~n6874 | ~n6883;
  assign n6885 = ~n571 & ~n580;
  assign n6886 = n18 & n659;
  assign n6887 = Ni36 & ~Ni32;
  assign n6888 = ~n873 & n877;
  assign n6889 = n6887 & ~n6888;
  assign n6890 = n750 & n3106;
  assign n6891 = Ni38 & n877;
  assign n6892 = ~n6890 & ~n6891;
  assign n6893 = n653 & n6892;
  assign n6894 = ~n6889 & ~n6893;
  assign n6895 = ~Ni45 & ~n874;
  assign n6896 = ~Ni38 & ~n6895;
  assign n6897 = ~n873 & ~n6896;
  assign n6898 = Ni38 & ~n928;
  assign n6899 = n6897 & ~n6898;
  assign n6900 = Ni36 & ~n928;
  assign n6901 = n6899 & ~n6900;
  assign n6902 = Ni32 & ~n6901;
  assign n6903 = n6894 & ~n6902;
  assign n6904 = n6886 & ~n6903;
  assign n6905 = n18 & n700;
  assign n6906 = n750 & n872;
  assign n6907 = n6905 & ~n6906;
  assign n6908 = Ni36 & n6905;
  assign n6909 = ~n6907 & ~n6908;
  assign n6910 = n18 & n870;
  assign n6911 = ~n1027_1 & n6910;
  assign n6912 = n18 & n703;
  assign n6913 = ~n1023 & n6912;
  assign n6914 = ~n6911 & ~n6913;
  assign n6915 = n6909 & n6914;
  assign n6916 = ~n6904 & n6915;
  assign n6917 = n1528 & ~n6916;
  assign n6918 = ~n1077_1 & n6912;
  assign n6919 = ~Ni32 & n822;
  assign n6920 = ~Ni41 & n6891;
  assign n6921 = ~n1053 & n6920;
  assign n6922 = ~n6890 & ~n6921;
  assign n6923 = n6919 & n6922;
  assign n6924 = ~Ni35 & ~Ni32;
  assign n6925 = ~Ni38 & ~n3106;
  assign n6926 = n891 & n6925;
  assign n6927 = ~n873 & ~n6926;
  assign n6928 = n878 & ~n1053;
  assign n6929 = ~n939 & ~n6928;
  assign n6930 = n6927 & ~n6929;
  assign n6931 = n6924 & ~n6930;
  assign n6932 = ~n6923 & ~n6931;
  assign n6933 = n1053 & n6887;
  assign n6934 = Ni41 & n6887;
  assign n6935 = ~n6889 & ~n6934;
  assign n6936 = ~n6933 & n6935;
  assign n6937 = n6932 & n6936;
  assign n6938 = Ni36 & Ni32;
  assign n6939 = n995 & ~n1053;
  assign n6940 = ~n873 & n6939;
  assign n6941 = n6938 & ~n6940;
  assign n6942 = ~Ni35 & Ni32;
  assign n6943 = n891 & n6896;
  assign n6944 = ~n939 & ~n6940;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = n6942 & ~n6945;
  assign n6947 = Ni35 & Ni32;
  assign n6948 = ~Ni36 & n6947;
  assign n6949 = Ni38 & ~n6939;
  assign n6950 = n6897 & ~n6949;
  assign n6951 = n6948 & ~n6950;
  assign n6952 = ~n6946 & ~n6951;
  assign n6953 = ~n6941 & n6952;
  assign n6954 = n6937 & n6953;
  assign n6955 = n6886 & ~n6954;
  assign n6956 = Ni35 & n6909;
  assign n6957 = ~Ni35 & ~n6907;
  assign n6958 = ~n890 & n6905;
  assign n6959 = n6957 & ~n6958;
  assign n6960 = ~n6956 & ~n6959;
  assign n6961 = ~n1086_1 & n6910;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = ~n6955 & n6962;
  assign n6964 = ~n6918 & n6963;
  assign n6965 = n949 & ~n6964;
  assign n6966 = n938 & n6925;
  assign n6967 = ~n873 & ~n6966;
  assign n6968 = n878 & ~n1036;
  assign n6969 = ~n926 & ~n6968;
  assign n6970 = n6967 & ~n6969;
  assign n6971 = n6924 & ~n6970;
  assign n6972 = n6935 & ~n6971;
  assign n6973 = n1036 & n6887;
  assign n6974 = ~n1036 & n6920;
  assign n6975 = ~n6890 & ~n6974;
  assign n6976 = n6919 & n6975;
  assign n6977 = ~n6973 & ~n6976;
  assign n6978 = n6972 & n6977;
  assign n6979 = n995 & ~n1036;
  assign n6980 = ~n873 & n6979;
  assign n6981 = n6938 & ~n6980;
  assign n6982 = n938 & n6896;
  assign n6983 = ~n926 & ~n6980;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = n6942 & ~n6984;
  assign n6986 = Ni38 & ~n6979;
  assign n6987 = n6897 & ~n6986;
  assign n6988 = n6948 & ~n6987;
  assign n6989 = ~n6985 & ~n6988;
  assign n6990 = ~n6981 & n6989;
  assign n6991 = n6978 & n6990;
  assign n6992 = n6886 & ~n6991;
  assign n6993 = ~Ni39 & n6905;
  assign n6994 = n6909 & ~n6993;
  assign n6995 = ~n6956 & ~n6994;
  assign n6996 = ~n899 & n6910;
  assign n6997 = ~n883 & n6912;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = ~n6995 & n6998;
  assign n7000 = ~n6992 & n6999;
  assign n7001 = n867 & ~n7000;
  assign n7002 = ~n6965 & ~n7001;
  assign n7003 = Pi21 & ~Pi20;
  assign n7004 = ~n6990 & n7003;
  assign n7005 = Pi21 & Pi20;
  assign n7006 = ~n6953 & n7005;
  assign n7007 = ~n7004 & ~n7006;
  assign n7008 = ~Pi22 & ~n7007;
  assign n7009 = ~n708 & n718;
  assign n7010 = n18 & n7009;
  assign n7011 = ~n864 & ~n7010;
  assign n7012 = ~Pi20 & n6978;
  assign n7013 = Pi20 & n6937;
  assign n7014 = ~Pi21 & ~n7013;
  assign n7015 = ~n7012 & n7014;
  assign n7016 = ~n7011 & ~n7015;
  assign n7017 = ~n7008 & n7016;
  assign n7018 = n7002 & n7017;
  assign n7019 = n869 & ~n7018;
  assign n7020 = ~n6890 & ~n6920;
  assign n7021 = n653 & n7020;
  assign n7022 = n6935 & ~n7021;
  assign n7023 = ~Pi21 & ~n7022;
  assign n7024 = Ni38 & ~n995;
  assign n7025 = n6897 & ~n7024;
  assign n7026 = Ni32 & ~n7025;
  assign n7027 = ~n995 & n6938;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = ~Pi22 & ~n7028;
  assign n7030 = ~n7011 & ~n7029;
  assign n7031 = ~n7023 & n7030;
  assign n7032 = n7022 & n7028;
  assign n7033 = n6886 & ~n7032;
  assign n7034 = ~n879 & n6912;
  assign n7035 = ~n1019 & n6910;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = ~n7033 & n7036;
  assign n7038 = n6909 & n7037;
  assign n7039 = n864 & ~n7038;
  assign n7040 = n7031 & ~n7039;
  assign n7041 = n730 & ~n7040;
  assign n7042 = n1610 & ~n7041;
  assign n7043 = ~Pi22 & n6902;
  assign n7044 = ~Pi21 & ~n6894;
  assign n7045 = ~n7011 & ~n7044;
  assign n7046 = ~n7043 & n7045;
  assign n7047 = Pi19 & ~n7046;
  assign n7048 = Pi17 & n7047;
  assign n7049 = n1672 & ~n7048;
  assign n7050 = ~n7042 & ~n7049;
  assign n7051 = ~n1010 & n6910;
  assign n7052 = ~n873 & ~n6943;
  assign n7053 = n927 & n928;
  assign n7054 = ~n939 & ~n7053;
  assign n7055 = n7052 & ~n7054;
  assign n7056 = Ni32 & ~n7055;
  assign n7057 = ~Ni37 & n6938;
  assign n7058 = ~n7053 & n7057;
  assign n7059 = ~n7056 & ~n7058;
  assign n7060 = n2029 & n3216;
  assign n7061 = ~n939 & ~n7060;
  assign n7062 = n6927 & ~n7061;
  assign n7063 = ~Ni32 & ~n7062;
  assign n7064 = n5092 & ~n7060;
  assign n7065 = ~n7063 & ~n7064;
  assign n7066 = n7059 & n7065;
  assign n7067 = n6886 & ~n7066;
  assign n7068 = ~n6907 & ~n6958;
  assign n7069 = ~n1006 & n6912;
  assign n7070 = n7068 & ~n7069;
  assign n7071 = ~n7067 & n7070;
  assign n7072 = ~n7051 & n7071;
  assign n7073 = n949 & ~n7072;
  assign n7074 = ~n1001 & n6910;
  assign n7075 = ~n873 & ~n6982;
  assign n7076 = ~n926 & ~n996;
  assign n7077 = n7075 & ~n7076;
  assign n7078 = Ni32 & ~n7077;
  assign n7079 = ~n996 & n7057;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = n2334 & n3216;
  assign n7082 = ~n926 & ~n7081;
  assign n7083 = n6967 & ~n7082;
  assign n7084 = ~Ni32 & ~n7083;
  assign n7085 = n5092 & ~n7081;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = n7080 & n7086;
  assign n7088 = n6886 & ~n7087;
  assign n7089 = ~n997 & n6912;
  assign n7090 = n6994 & ~n7089;
  assign n7091 = ~n7088 & n7090;
  assign n7092 = ~n7074 & n7091;
  assign n7093 = n867 & ~n7092;
  assign n7094 = ~n7073 & ~n7093;
  assign n7095 = Pi20 & n7065;
  assign n7096 = ~Pi20 & n7086;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~Pi21 & n7097;
  assign n7099 = n7003 & ~n7080;
  assign n7100 = n7005 & ~n7059;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = ~Pi22 & ~n7101;
  assign n7103 = ~n7011 & ~n7102;
  assign n7104 = ~n7098 & n7103;
  assign n7105 = n7094 & n7104;
  assign n7106 = n994 & ~n7105;
  assign n7107 = ~n7050 & ~n7106;
  assign n7108 = ~n7019 & n7107;
  assign n7109 = ~n6917 & n7108;
  assign n7110 = ~n1100 & n6910;
  assign n7111 = n878 & ~n973;
  assign n7112 = ~n939 & ~n7111;
  assign n7113 = n6927 & ~n7112;
  assign n7114 = n856 & ~n7113;
  assign n7115 = ~Ni32 & n908;
  assign n7116 = ~n973 & n6920;
  assign n7117 = ~n6890 & ~n7116;
  assign n7118 = n7115 & n7117;
  assign n7119 = ~n7114 & ~n7118;
  assign n7120 = n973 & n6887;
  assign n7121 = n6935 & ~n7120;
  assign n7122 = n7119 & n7121;
  assign n7123 = ~n973 & n995;
  assign n7124 = ~n873 & n7123;
  assign n7125 = n6938 & ~n7124;
  assign n7126 = ~n939 & ~n7124;
  assign n7127 = ~n6943 & ~n7126;
  assign n7128 = n6947 & ~n7127;
  assign n7129 = Ni38 & ~n7123;
  assign n7130 = n6897 & ~n7129;
  assign n7131 = Ni32 & n908;
  assign n7132 = ~n7130 & n7131;
  assign n7133 = ~n7128 & ~n7132;
  assign n7134 = ~n7125 & n7133;
  assign n7135 = n7122 & n7134;
  assign n7136 = n6886 & ~n7135;
  assign n7137 = ~Ni35 & n6909;
  assign n7138 = Ni35 & n7068;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = ~n1091 & n6912;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = ~n7136 & n7141;
  assign n7143 = ~n7110 & n7142;
  assign n7144 = n949 & ~n7143;
  assign n7145 = ~n956 & n6920;
  assign n7146 = ~n6890 & ~n7145;
  assign n7147 = n7115 & n7146;
  assign n7148 = n878 & ~n956;
  assign n7149 = ~n926 & ~n7148;
  assign n7150 = n6967 & ~n7149;
  assign n7151 = n856 & ~n7150;
  assign n7152 = ~n7147 & ~n7151;
  assign n7153 = n956 & n6887;
  assign n7154 = n6935 & ~n7153;
  assign n7155 = n7152 & n7154;
  assign n7156 = ~n956 & n995;
  assign n7157 = ~n873 & n7156;
  assign n7158 = n6938 & ~n7157;
  assign n7159 = ~n926 & ~n7157;
  assign n7160 = ~n6982 & ~n7159;
  assign n7161 = n6947 & ~n7160;
  assign n7162 = Ni38 & ~n7156;
  assign n7163 = n6897 & ~n7162;
  assign n7164 = n7131 & ~n7163;
  assign n7165 = ~n7161 & ~n7164;
  assign n7166 = ~n7158 & n7165;
  assign n7167 = n7155 & n7166;
  assign n7168 = n6886 & ~n7167;
  assign n7169 = ~n917 & n6910;
  assign n7170 = ~n905 & n6912;
  assign n7171 = ~n6994 & ~n7137;
  assign n7172 = ~n7170 & ~n7171;
  assign n7173 = ~n7169 & n7172;
  assign n7174 = ~n7168 & n7173;
  assign n7175 = n867 & ~n7174;
  assign n7176 = ~n7144 & ~n7175;
  assign n7177 = n7003 & ~n7166;
  assign n7178 = n7005 & ~n7134;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = ~Pi22 & ~n7179;
  assign n7181 = ~Pi20 & n7155;
  assign n7182 = Pi20 & n7122;
  assign n7183 = ~Pi21 & ~n7182;
  assign n7184 = ~n7181 & n7183;
  assign n7185 = ~n7011 & ~n7184;
  assign n7186 = ~n7180 & n7185;
  assign n7187 = n7176 & n7186;
  assign n7188 = n903 & ~n7187;
  assign n7189 = ~n959 & n6912;
  assign n7190 = ~n965 & n6938;
  assign n7191 = ~n926 & ~n965;
  assign n7192 = ~n6982 & ~n7191;
  assign n7193 = n6947 & ~n7192;
  assign n7194 = Ni38 & ~n958;
  assign n7195 = n6897 & ~n7194;
  assign n7196 = n7131 & ~n7195;
  assign n7197 = ~n7193 & ~n7196;
  assign n7198 = ~n7190 & n7197;
  assign n7199 = n877 & ~n957;
  assign n7200 = ~n892 & ~n7199;
  assign n7201 = ~n957 & n6891;
  assign n7202 = Ni37 & ~n7201;
  assign n7203 = ~n7200 & ~n7202;
  assign n7204 = ~n6966 & n7203;
  assign n7205 = n856 & ~n7204;
  assign n7206 = ~n6890 & ~n7201;
  assign n7207 = n7115 & n7206;
  assign n7208 = n957 & n6887;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = ~n6889 & n7209;
  assign n7211 = ~n7205 & n7210;
  assign n7212 = n7198 & n7211;
  assign n7213 = n6886 & ~n7212;
  assign n7214 = ~n969 & n6910;
  assign n7215 = ~n7171 & ~n7214;
  assign n7216 = ~n7213 & n7215;
  assign n7217 = ~n7189 & n7216;
  assign n7218 = n867 & ~n7217;
  assign n7219 = ~n988 & n6910;
  assign n7220 = ~n984 & n6938;
  assign n7221 = ~n939 & ~n984;
  assign n7222 = ~n6943 & ~n7221;
  assign n7223 = n6947 & ~n7222;
  assign n7224 = Ni38 & ~n975;
  assign n7225 = n6897 & ~n7224;
  assign n7226 = n7131 & ~n7225;
  assign n7227 = ~n7223 & ~n7226;
  assign n7228 = ~n7220 & n7227;
  assign n7229 = n877 & ~n974;
  assign n7230 = ~n980 & ~n7229;
  assign n7231 = ~n974 & n6891;
  assign n7232 = Ni37 & ~n7231;
  assign n7233 = ~n7230 & ~n7232;
  assign n7234 = ~n6926 & n7233;
  assign n7235 = n856 & ~n7234;
  assign n7236 = ~n6890 & ~n7231;
  assign n7237 = n7115 & n7236;
  assign n7238 = n974 & n6887;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = ~n6889 & n7239;
  assign n7241 = ~n7235 & n7240;
  assign n7242 = n7228 & n7241;
  assign n7243 = n6886 & ~n7242;
  assign n7244 = ~n976 & n6912;
  assign n7245 = ~n7139 & ~n7244;
  assign n7246 = ~n7243 & n7245;
  assign n7247 = ~n7219 & n7246;
  assign n7248 = n949 & ~n7247;
  assign n7249 = ~n7218 & ~n7248;
  assign n7250 = n7003 & ~n7198;
  assign n7251 = n7005 & ~n7228;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = ~Pi22 & ~n7252;
  assign n7254 = Pi20 & n7241;
  assign n7255 = ~Pi20 & n7211;
  assign n7256 = ~Pi21 & ~n7255;
  assign n7257 = ~n7254 & n7256;
  assign n7258 = ~n7011 & ~n7257;
  assign n7259 = ~n7253 & n7258;
  assign n7260 = n7249 & n7259;
  assign n7261 = n955 & ~n7260;
  assign n7262 = ~n7188 & ~n7261;
  assign n7263 = ~n1056 & n6912;
  assign n7264 = ~n1063 & n6938;
  assign n7265 = ~n939 & ~n1063;
  assign n7266 = ~n6943 & ~n7265;
  assign n7267 = n6942 & ~n7266;
  assign n7268 = Ni38 & ~n1055;
  assign n7269 = n6897 & ~n7268;
  assign n7270 = n6948 & ~n7269;
  assign n7271 = ~n7267 & ~n7270;
  assign n7272 = ~n7264 & n7271;
  assign n7273 = n877 & ~n1054;
  assign n7274 = ~n980 & ~n7273;
  assign n7275 = ~n1054 & n6891;
  assign n7276 = Ni37 & ~n7275;
  assign n7277 = ~n7274 & ~n7276;
  assign n7278 = ~n6926 & n7277;
  assign n7279 = n6924 & ~n7278;
  assign n7280 = ~n6890 & ~n7275;
  assign n7281 = n6919 & n7280;
  assign n7282 = ~Ni41 & n6933;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 = ~n6889 & n7283;
  assign n7285 = ~n7279 & n7284;
  assign n7286 = n7272 & n7285;
  assign n7287 = n6886 & ~n7286;
  assign n7288 = ~n1067 & n6910;
  assign n7289 = ~n6960 & ~n7288;
  assign n7290 = ~n7287 & n7289;
  assign n7291 = ~n7263 & n7290;
  assign n7292 = n949 & ~n7291;
  assign n7293 = ~n1045 & n6938;
  assign n7294 = ~n926 & ~n1045;
  assign n7295 = ~n6982 & ~n7294;
  assign n7296 = n6942 & ~n7295;
  assign n7297 = Ni38 & ~n1038;
  assign n7298 = n6897 & ~n7297;
  assign n7299 = n6948 & ~n7298;
  assign n7300 = ~n7296 & ~n7299;
  assign n7301 = ~n7293 & n7300;
  assign n7302 = n7003 & ~n7301;
  assign n7303 = n7005 & ~n7272;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = ~Pi22 & ~n7304;
  assign n7306 = ~n7011 & ~n7305;
  assign n7307 = n877 & ~n1037;
  assign n7308 = ~n892 & ~n7307;
  assign n7309 = ~n1037 & n6891;
  assign n7310 = Ni37 & ~n7309;
  assign n7311 = ~n7308 & ~n7310;
  assign n7312 = ~n6966 & n7311;
  assign n7313 = n6924 & ~n7312;
  assign n7314 = ~n6890 & ~n7309;
  assign n7315 = n6919 & n7314;
  assign n7316 = ~Ni41 & n6973;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = ~n6889 & n7317;
  assign n7319 = ~n7313 & n7318;
  assign n7320 = ~Pi20 & n7319;
  assign n7321 = Pi20 & n7285;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = ~Pi21 & n7322;
  assign n7324 = n7306 & ~n7323;
  assign n7325 = n7301 & n7319;
  assign n7326 = n6886 & ~n7325;
  assign n7327 = ~n1049 & n6910;
  assign n7328 = ~n1039 & n6912;
  assign n7329 = ~n7327 & ~n7328;
  assign n7330 = ~n7326 & n7329;
  assign n7331 = ~n6995 & n7330;
  assign n7332 = n867 & ~n7331;
  assign n7333 = n7324 & ~n7332;
  assign n7334 = ~n7292 & n7333;
  assign n7335 = n1035 & ~n7334;
  assign n7336 = ~n930 & n6912;
  assign n7337 = ~n926 & ~n929;
  assign n7338 = n7075 & ~n7337;
  assign n7339 = Ni32 & ~n7338;
  assign n7340 = ~n929 & n7057;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = n877 & ~n927;
  assign n7343 = ~n926 & ~n7342;
  assign n7344 = n6967 & ~n7343;
  assign n7345 = ~Ni32 & ~n7344;
  assign n7346 = n5092 & ~n7342;
  assign n7347 = ~n7345 & ~n7346;
  assign n7348 = n7341 & n7347;
  assign n7349 = n6886 & ~n7348;
  assign n7350 = ~n934 & n6910;
  assign n7351 = n6994 & ~n7350;
  assign n7352 = ~n7349 & n7351;
  assign n7353 = ~n7336 & n7352;
  assign n7354 = n867 & ~n7353;
  assign n7355 = ~n946 & n6910;
  assign n7356 = ~n941 & n7057;
  assign n7357 = ~n939 & ~n941;
  assign n7358 = n7052 & ~n7357;
  assign n7359 = Ni32 & ~n7358;
  assign n7360 = ~n7356 & ~n7359;
  assign n7361 = n877 & ~n940;
  assign n7362 = n5092 & ~n7361;
  assign n7363 = ~n939 & ~n7361;
  assign n7364 = n6927 & ~n7363;
  assign n7365 = ~Ni32 & ~n7364;
  assign n7366 = ~n7362 & ~n7365;
  assign n7367 = n7360 & n7366;
  assign n7368 = n6886 & ~n7367;
  assign n7369 = ~n942 & n6912;
  assign n7370 = n7068 & ~n7369;
  assign n7371 = ~n7368 & n7370;
  assign n7372 = ~n7355 & n7371;
  assign n7373 = n949 & ~n7372;
  assign n7374 = ~n7354 & ~n7373;
  assign n7375 = n7003 & ~n7341;
  assign n7376 = n7005 & ~n7360;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = ~Pi22 & ~n7377;
  assign n7379 = ~Pi20 & n7347;
  assign n7380 = Pi20 & n7366;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = ~Pi21 & n7381;
  assign n7383 = ~n7378 & ~n7382;
  assign n7384 = ~n7011 & n7383;
  assign n7385 = n7374 & n7384;
  assign n7386 = n924 & ~n7385;
  assign n7387 = ~n7335 & ~n7386;
  assign n7388 = n7262 & n7387;
  assign n7389 = n7109 & n7388;
  assign n7390 = ~n1121 & n6910;
  assign n7391 = ~n6938 & ~n6942;
  assign n7392 = ~n7163 & ~n7391;
  assign n7393 = ~n7161 & ~n7392;
  assign n7394 = ~Ni32 & ~n822;
  assign n7395 = n7146 & n7394;
  assign n7396 = ~n7151 & ~n7395;
  assign n7397 = n7393 & n7396;
  assign n7398 = n6886 & ~n7397;
  assign n7399 = ~n816 & n6993;
  assign n7400 = ~n6907 & ~n7399;
  assign n7401 = ~n6957 & ~n7400;
  assign n7402 = ~n7170 & ~n7401;
  assign n7403 = ~n7398 & n7402;
  assign n7404 = ~n7390 & n7403;
  assign n7405 = n867 & ~n7404;
  assign n7406 = n7003 & ~n7393;
  assign n7407 = ~n7130 & ~n7391;
  assign n7408 = ~n7128 & ~n7407;
  assign n7409 = n7005 & ~n7408;
  assign n7410 = ~n7406 & ~n7409;
  assign n7411 = ~Pi22 & ~n7410;
  assign n7412 = ~Pi20 & n7396;
  assign n7413 = n7117 & n7394;
  assign n7414 = ~n7114 & ~n7413;
  assign n7415 = Pi20 & n7414;
  assign n7416 = ~n7412 & ~n7415;
  assign n7417 = ~Pi21 & n7416;
  assign n7418 = ~n7011 & ~n7417;
  assign n7419 = ~n7411 & n7418;
  assign n7420 = n7408 & n7414;
  assign n7421 = n6886 & ~n7420;
  assign n7422 = ~n1141 & n6910;
  assign n7423 = Ni39 & ~n816;
  assign n7424 = n6905 & n7423;
  assign n7425 = ~n6907 & ~n7424;
  assign n7426 = ~n6957 & ~n7425;
  assign n7427 = ~n7140 & ~n7426;
  assign n7428 = ~n7422 & n7427;
  assign n7429 = ~n7421 & n7428;
  assign n7430 = n949 & ~n7429;
  assign n7431 = n7419 & ~n7430;
  assign n7432 = ~n7405 & n7431;
  assign n7433 = n903 & ~n7432;
  assign n7434 = n1110 & n6910;
  assign n7435 = n6896 & n6938;
  assign n7436 = Ni38 & n7079;
  assign n7437 = ~n7078 & ~n7436;
  assign n7438 = ~n7435 & n7437;
  assign n7439 = n5092 & n6925;
  assign n7440 = Ni38 & n7085;
  assign n7441 = ~n7084 & ~n7440;
  assign n7442 = ~n7439 & n7441;
  assign n7443 = n7438 & n7442;
  assign n7444 = n6886 & ~n7443;
  assign n7445 = ~n7089 & n7400;
  assign n7446 = ~n7444 & n7445;
  assign n7447 = ~n7434 & n7446;
  assign n7448 = n867 & ~n7447;
  assign n7449 = n7003 & ~n7438;
  assign n7450 = Ni38 & n7058;
  assign n7451 = ~n7056 & ~n7450;
  assign n7452 = ~n7435 & n7451;
  assign n7453 = n7005 & ~n7452;
  assign n7454 = ~n7449 & ~n7453;
  assign n7455 = ~Pi22 & ~n7454;
  assign n7456 = Ni38 & n7064;
  assign n7457 = ~n7063 & ~n7456;
  assign n7458 = ~n7439 & n7457;
  assign n7459 = Pi20 & n7458;
  assign n7460 = ~Pi20 & n7442;
  assign n7461 = ~Pi21 & ~n7460;
  assign n7462 = ~n7459 & n7461;
  assign n7463 = ~n7455 & ~n7462;
  assign n7464 = n7452 & n7458;
  assign n7465 = n6886 & ~n7464;
  assign n7466 = ~n1114 & n7051;
  assign n7467 = n7425 & ~n7466;
  assign n7468 = ~n7069 & n7467;
  assign n7469 = ~n7465 & n7468;
  assign n7470 = n949 & ~n7469;
  assign n7471 = n7463 & ~n7470;
  assign n7472 = ~n7011 & n7471;
  assign n7473 = ~n7448 & n7472;
  assign n7474 = n994 & ~n7473;
  assign n7475 = n1146 & n6910;
  assign n7476 = Ni38 & n7356;
  assign n7477 = ~n7359 & ~n7476;
  assign n7478 = ~n7435 & n7477;
  assign n7479 = Ni38 & n7362;
  assign n7480 = ~n7365 & ~n7479;
  assign n7481 = ~n7439 & n7480;
  assign n7482 = n7478 & n7481;
  assign n7483 = n6886 & ~n7482;
  assign n7484 = ~n7369 & n7425;
  assign n7485 = ~n7483 & n7484;
  assign n7486 = ~n7475 & n7485;
  assign n7487 = n949 & ~n7486;
  assign n7488 = Ni38 & n7340;
  assign n7489 = ~n7435 & ~n7488;
  assign n7490 = ~n7339 & n7489;
  assign n7491 = n7003 & ~n7490;
  assign n7492 = n7005 & ~n7478;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = ~Pi22 & ~n7493;
  assign n7495 = Ni38 & n7346;
  assign n7496 = ~n7439 & ~n7495;
  assign n7497 = ~n7345 & n7496;
  assign n7498 = ~Pi20 & n7497;
  assign n7499 = Pi20 & n7481;
  assign n7500 = ~Pi21 & ~n7499;
  assign n7501 = ~n7498 & n7500;
  assign n7502 = ~n7494 & ~n7501;
  assign n7503 = ~n1131 & n6910;
  assign n7504 = n7490 & n7497;
  assign n7505 = n6886 & ~n7504;
  assign n7506 = ~n7336 & n7400;
  assign n7507 = ~n7505 & n7506;
  assign n7508 = ~n7503 & n7507;
  assign n7509 = n867 & ~n7508;
  assign n7510 = ~n7011 & ~n7509;
  assign n7511 = n7502 & n7510;
  assign n7512 = ~n7487 & n7511;
  assign n7513 = n924 & ~n7512;
  assign n7514 = ~n6938 & ~n6947;
  assign n7515 = ~n7298 & ~n7514;
  assign n7516 = ~n7296 & ~n7515;
  assign n7517 = ~Ni32 & ~n908;
  assign n7518 = n7314 & n7517;
  assign n7519 = ~n7313 & ~n7518;
  assign n7520 = n7516 & n7519;
  assign n7521 = n6886 & ~n7520;
  assign n7522 = Ni35 & ~n6907;
  assign n7523 = ~n7400 & ~n7522;
  assign n7524 = ~n1164 & n6910;
  assign n7525 = ~n7328 & ~n7524;
  assign n7526 = ~n7523 & n7525;
  assign n7527 = ~n7521 & n7526;
  assign n7528 = n867 & ~n7527;
  assign n7529 = ~n7269 & ~n7514;
  assign n7530 = ~n7267 & ~n7529;
  assign n7531 = n7280 & n7517;
  assign n7532 = ~n7279 & ~n7531;
  assign n7533 = n7530 & n7532;
  assign n7534 = n6886 & ~n7533;
  assign n7535 = ~n7425 & ~n7522;
  assign n7536 = ~n1168 & n6910;
  assign n7537 = ~n7263 & ~n7536;
  assign n7538 = ~n7535 & n7537;
  assign n7539 = ~n7534 & n7538;
  assign n7540 = n949 & ~n7539;
  assign n7541 = ~n7528 & ~n7540;
  assign n7542 = Pi20 & n7532;
  assign n7543 = ~Pi20 & n7519;
  assign n7544 = ~Pi21 & ~n7543;
  assign n7545 = ~n7542 & n7544;
  assign n7546 = n7003 & ~n7516;
  assign n7547 = n7005 & ~n7530;
  assign n7548 = ~n7546 & ~n7547;
  assign n7549 = ~Pi22 & ~n7548;
  assign n7550 = ~n7011 & ~n7549;
  assign n7551 = ~n7545 & n7550;
  assign n7552 = n7541 & n7551;
  assign n7553 = n1035 & ~n7552;
  assign n7554 = ~Pi22 & ~n7025;
  assign n7555 = ~Pi21 & n7020;
  assign n7556 = ~n7011 & ~n7555;
  assign n7557 = ~n7554 & n7556;
  assign n7558 = ~n1017 & n6910;
  assign n7559 = ~n6907 & ~n7558;
  assign n7560 = n659 & n7026;
  assign n7561 = ~Ni32 & n6886;
  assign n7562 = n7020 & n7561;
  assign n7563 = ~n7034 & ~n7562;
  assign n7564 = ~n7560 & n7563;
  assign n7565 = n7559 & n7564;
  assign n7566 = n864 & ~n7565;
  assign n7567 = n7557 & ~n7566;
  assign n7568 = n730 & ~n7567;
  assign n7569 = n1178 & ~n7568;
  assign n7570 = ~n6907 & ~n6913;
  assign n7571 = ~n1025 & n6910;
  assign n7572 = n6892 & n7561;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = n707 & ~n6899;
  assign n7575 = n7573 & ~n7574;
  assign n7576 = n7570 & n7575;
  assign n7577 = n1030 & ~n7576;
  assign n7578 = ~Pi22 & ~n6899;
  assign n7579 = ~Pi21 & n6892;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n7011 & n7580;
  assign n7582 = Pi19 & ~n7581;
  assign n7583 = Pi17 & n7582;
  assign n7584 = ~n7577 & ~n7583;
  assign n7585 = n1769 & n7584;
  assign n7586 = ~n7569 & ~n7585;
  assign n7587 = ~n7553 & ~n7586;
  assign n7588 = ~n7513 & n7587;
  assign n7589 = ~n7474 & n7588;
  assign n7590 = ~n1137 & n6910;
  assign n7591 = ~n6950 & ~n7514;
  assign n7592 = ~n6946 & ~n7591;
  assign n7593 = n6922 & n7517;
  assign n7594 = ~n6931 & ~n7593;
  assign n7595 = n7592 & n7594;
  assign n7596 = n6886 & ~n7595;
  assign n7597 = ~n6918 & ~n7535;
  assign n7598 = ~n7596 & n7597;
  assign n7599 = ~n7590 & n7598;
  assign n7600 = n949 & ~n7599;
  assign n7601 = ~n6987 & ~n7514;
  assign n7602 = ~n6985 & ~n7601;
  assign n7603 = n6975 & n7517;
  assign n7604 = ~n6971 & ~n7603;
  assign n7605 = n7602 & n7604;
  assign n7606 = n6886 & ~n7605;
  assign n7607 = ~n1125 & n6910;
  assign n7608 = ~n6997 & ~n7523;
  assign n7609 = ~n7607 & n7608;
  assign n7610 = ~n7606 & n7609;
  assign n7611 = n867 & ~n7610;
  assign n7612 = ~n7600 & ~n7611;
  assign n7613 = n7003 & ~n7602;
  assign n7614 = n7005 & ~n7592;
  assign n7615 = ~n7613 & ~n7614;
  assign n7616 = ~Pi22 & ~n7615;
  assign n7617 = ~Pi20 & n7604;
  assign n7618 = Pi20 & n7594;
  assign n7619 = ~n7617 & ~n7618;
  assign n7620 = ~Pi21 & n7619;
  assign n7621 = ~n7011 & ~n7620;
  assign n7622 = ~n7616 & n7621;
  assign n7623 = n7612 & n7622;
  assign n7624 = n869 & ~n7623;
  assign n7625 = n7206 & n7394;
  assign n7626 = ~n7205 & ~n7625;
  assign n7627 = ~n7195 & ~n7391;
  assign n7628 = ~n7193 & ~n7627;
  assign n7629 = n7626 & n7628;
  assign n7630 = n6886 & ~n7629;
  assign n7631 = ~n1154 & n6910;
  assign n7632 = ~n7189 & ~n7401;
  assign n7633 = ~n7631 & n7632;
  assign n7634 = ~n7630 & n7633;
  assign n7635 = n867 & ~n7634;
  assign n7636 = n7236 & n7394;
  assign n7637 = ~n7235 & ~n7636;
  assign n7638 = ~n7225 & ~n7391;
  assign n7639 = ~n7223 & ~n7638;
  assign n7640 = n7637 & n7639;
  assign n7641 = n6886 & ~n7640;
  assign n7642 = ~n1158 & n6910;
  assign n7643 = ~n7244 & ~n7642;
  assign n7644 = ~n7641 & n7643;
  assign n7645 = ~n7426 & n7644;
  assign n7646 = n949 & ~n7645;
  assign n7647 = ~n7635 & ~n7646;
  assign n7648 = ~Pi20 & n7626;
  assign n7649 = Pi20 & n7637;
  assign n7650 = ~Pi21 & ~n7649;
  assign n7651 = ~n7648 & n7650;
  assign n7652 = n7003 & ~n7628;
  assign n7653 = n7005 & ~n7639;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~Pi22 & ~n7654;
  assign n7656 = ~n7011 & ~n7655;
  assign n7657 = ~n7651 & n7656;
  assign n7658 = n7647 & n7657;
  assign n7659 = n955 & ~n7658;
  assign n7660 = ~n7624 & ~n7659;
  assign n7661 = n7589 & n7660;
  assign n7662 = ~n7433 & n7661;
  assign n7663 = P__cmxcl_1 & ~n7662;
  assign n7664 = ~n7389 & n7663;
  assign n7665 = n18 & ~n7664;
  assign n7666 = n6885 & n7665;
  assign n7667 = ~n18 & ~n1068;
  assign n7668 = n7291 & ~n7667;
  assign n7669 = n1643 & ~n7668;
  assign n7670 = ~Pi19 & ~n7324;
  assign n7671 = ~n18 & ~n1050;
  assign n7672 = n7331 & ~n7671;
  assign n7673 = n1625 & ~n7672;
  assign n7674 = ~n18 & ~n1174;
  assign n7675 = ~n1346 & ~n7674;
  assign n7676 = n6916 & n7675;
  assign n7677 = n1814 & ~n7676;
  assign n7678 = ~n7047 & ~n7677;
  assign n7679 = ~n7673 & n7678;
  assign n7680 = ~n7670 & n7679;
  assign n7681 = ~n7669 & n7680;
  assign n7682 = n1672 & ~n7681;
  assign n7683 = Pi19 & ~n7557;
  assign n7684 = ~n18 & ~n1126;
  assign n7685 = n7610 & ~n7684;
  assign n7686 = n1625 & ~n7685;
  assign n7687 = ~Pi19 & ~n7622;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n18 & ~n1138;
  assign n7690 = n7599 & ~n7689;
  assign n7691 = n1643 & ~n7690;
  assign n7692 = ~n18 & ~n1179;
  assign n7693 = n7565 & ~n7692;
  assign n7694 = n1814 & ~n7693;
  assign n7695 = ~n7691 & ~n7694;
  assign n7696 = n7688 & n7695;
  assign n7697 = ~n7683 & n7696;
  assign n7698 = n1178 & ~n7697;
  assign n7699 = ~n18 & ~n1169;
  assign n7700 = n7539 & ~n7699;
  assign n7701 = n1643 & ~n7700;
  assign n7702 = n7576 & ~n7674;
  assign n7703 = n1814 & ~n7702;
  assign n7704 = ~n7582 & ~n7703;
  assign n7705 = ~Pi19 & ~n7551;
  assign n7706 = ~n18 & ~n1165;
  assign n7707 = n7527 & ~n7706;
  assign n7708 = n1625 & ~n7707;
  assign n7709 = ~n7705 & ~n7708;
  assign n7710 = n7704 & n7709;
  assign n7711 = ~n7701 & n7710;
  assign n7712 = n1769 & ~n7711;
  assign n7713 = ~n18 & ~n1087;
  assign n7714 = n6964 & ~n7713;
  assign n7715 = n1643 & ~n7714;
  assign n7716 = ~Pi19 & ~n7017;
  assign n7717 = ~n7715 & ~n7716;
  assign n7718 = ~n18 & ~n1020;
  assign n7719 = n7038 & ~n7718;
  assign n7720 = n1814 & ~n7719;
  assign n7721 = ~n18 & ~n900;
  assign n7722 = n7000 & ~n7721;
  assign n7723 = n1625 & ~n7722;
  assign n7724 = Pi19 & ~n7031;
  assign n7725 = ~n7723 & ~n7724;
  assign n7726 = ~n7720 & n7725;
  assign n7727 = n7717 & n7726;
  assign n7728 = n1610 & ~n7727;
  assign n7729 = ~n7712 & ~n7728;
  assign n7730 = ~n7698 & n7729;
  assign n7731 = ~n7682 & n7730;
  assign n7732 = Pi17 & n7731;
  assign n7733 = ~n18 & ~n1142;
  assign n7734 = n7429 & ~n7733;
  assign n7735 = n1611 & ~n7734;
  assign n7736 = ~n18 & ~n1116;
  assign n7737 = n7469 & ~n7736;
  assign n7738 = n1643 & ~n7737;
  assign n7739 = ~n7735 & ~n7738;
  assign n7740 = ~n18 & ~n1111;
  assign n7741 = n7447 & ~n7740;
  assign n7742 = n1625 & ~n7741;
  assign n7743 = n7419 & ~n7742;
  assign n7744 = ~n18 & ~n1122;
  assign n7745 = n7404 & ~n7744;
  assign n7746 = n1636 & ~n7745;
  assign n7747 = ~Pi19 & ~n7463;
  assign n7748 = ~n7746 & ~n7747;
  assign n7749 = n7743 & n7748;
  assign n7750 = n7739 & n7749;
  assign n7751 = n1178 & ~n7750;
  assign n7752 = ~n18 & ~n1011;
  assign n7753 = n7072 & ~n7752;
  assign n7754 = n1643 & ~n7753;
  assign n7755 = ~n18 & ~n1101;
  assign n7756 = n7143 & ~n7755;
  assign n7757 = n1611 & ~n7756;
  assign n7758 = n7186 & ~n7757;
  assign n7759 = ~n18 & ~n918;
  assign n7760 = n7174 & ~n7759;
  assign n7761 = n1636 & ~n7760;
  assign n7762 = ~Pi19 & ~n7104;
  assign n7763 = ~n18 & ~n1002_1;
  assign n7764 = n7092 & ~n7763;
  assign n7765 = n1625 & ~n7764;
  assign n7766 = ~n7762 & ~n7765;
  assign n7767 = ~n7761 & n7766;
  assign n7768 = n7758 & n7767;
  assign n7769 = ~n7754 & n7768;
  assign n7770 = n1610 & ~n7769;
  assign n7771 = ~n18 & ~n1159;
  assign n7772 = n7645 & ~n7771;
  assign n7773 = n1611 & ~n7772;
  assign n7774 = ~n18 & ~n1147;
  assign n7775 = n7486 & ~n7774;
  assign n7776 = n1643 & ~n7775;
  assign n7777 = ~n18 & ~n1155;
  assign n7778 = n7634 & ~n7777;
  assign n7779 = n1636 & ~n7778;
  assign n7780 = n7657 & ~n7779;
  assign n7781 = ~n7776 & n7780;
  assign n7782 = ~Pi19 & ~n7502;
  assign n7783 = ~n18 & ~n1132;
  assign n7784 = n7508 & ~n7783;
  assign n7785 = n1625 & ~n7784;
  assign n7786 = ~n7782 & ~n7785;
  assign n7787 = n7781 & n7786;
  assign n7788 = ~n7773 & n7787;
  assign n7789 = n1769 & ~n7788;
  assign n7790 = ~n18 & ~n970;
  assign n7791 = n7217 & ~n7790;
  assign n7792 = n1636 & ~n7791;
  assign n7793 = ~n18 & ~n989;
  assign n7794 = n7247 & ~n7793;
  assign n7795 = n1611 & ~n7794;
  assign n7796 = ~n18 & ~n935;
  assign n7797 = n7353 & ~n7796;
  assign n7798 = n1625 & ~n7797;
  assign n7799 = ~n7795 & ~n7798;
  assign n7800 = ~Pi19 & ~n7383;
  assign n7801 = ~n18 & ~n947;
  assign n7802 = n7372 & ~n7801;
  assign n7803 = n1643 & ~n7802;
  assign n7804 = ~n7800 & ~n7803;
  assign n7805 = n7259 & n7804;
  assign n7806 = n7799 & n7805;
  assign n7807 = ~n7792 & n7806;
  assign n7808 = n1672 & ~n7807;
  assign n7809 = ~n7789 & ~n7808;
  assign n7810 = ~n7770 & n7809;
  assign n7811 = ~n7751 & n7810;
  assign n7812 = ~Pi17 & n7811;
  assign n7813 = ~n863 & ~n7812;
  assign n7814 = ~n7732 & n7813;
  assign n7815 = ~Pi25 & ~n7647;
  assign n7816 = n950 & ~n7772;
  assign n7817 = n868 & ~n7778;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = n7657 & n7818;
  assign n7820 = ~n7815 & n7819;
  assign n7821 = n738 & ~n7820;
  assign n7822 = ~Pi25 & n1191;
  assign n7823 = n1031 & ~n7702;
  assign n7824 = ~n7822 & ~n7823;
  assign n7825 = n7584 & n7824;
  assign n7826 = ~Pi25 & ~n7541;
  assign n7827 = n868 & ~n7707;
  assign n7828 = n950 & ~n7700;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = n7551 & n7829;
  assign n7831 = ~n7826 & n7830;
  assign n7832 = n736 & ~n7831;
  assign n7833 = n950 & n7774;
  assign n7834 = n868 & n7783;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = n7512 & n7835;
  assign n7837 = n923 & ~n7836;
  assign n7838 = ~n7832 & ~n7837;
  assign n7839 = n7825 & n7838;
  assign n7840 = ~n7821 & n7839;
  assign n7841 = n1769 & ~n7840;
  assign n7842 = n950 & ~n7753;
  assign n7843 = ~Pi25 & ~n7094;
  assign n7844 = n868 & ~n7764;
  assign n7845 = n7104 & ~n7844;
  assign n7846 = ~n7843 & n7845;
  assign n7847 = ~n7842 & n7846;
  assign n7848 = n923 & ~n7847;
  assign n7849 = n868 & ~n7722;
  assign n7850 = ~Pi25 & ~n7002;
  assign n7851 = n950 & ~n7714;
  assign n7852 = n7017 & ~n7851;
  assign n7853 = ~n7850 & n7852;
  assign n7854 = ~n7849 & n7853;
  assign n7855 = n736 & ~n7854;
  assign n7856 = ~Pi25 & ~n7176;
  assign n7857 = n950 & ~n7756;
  assign n7858 = n868 & ~n7760;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = n7186 & n7859;
  assign n7861 = ~n7856 & n7860;
  assign n7862 = n738 & ~n7861;
  assign n7863 = n1031 & ~n7719;
  assign n7864 = ~n7041 & ~n7863;
  assign n7865 = ~n7822 & n7864;
  assign n7866 = ~n7862 & n7865;
  assign n7867 = ~n7855 & n7866;
  assign n7868 = ~n7848 & n7867;
  assign n7869 = n1610 & ~n7868;
  assign n7870 = n1031 & ~n7693;
  assign n7871 = n867 & n7744;
  assign n7872 = n949 & n7733;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = Pi25 & ~n7873;
  assign n7875 = n7432 & ~n7874;
  assign n7876 = n738 & ~n7875;
  assign n7877 = n868 & n7740;
  assign n7878 = n950 & n7736;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = n7473 & n7879;
  assign n7881 = n923 & ~n7880;
  assign n7882 = ~n7876 & ~n7881;
  assign n7883 = n950 & ~n7690;
  assign n7884 = ~Pi25 & ~n7612;
  assign n7885 = n868 & ~n7685;
  assign n7886 = n7622 & ~n7885;
  assign n7887 = ~n7884 & n7886;
  assign n7888 = ~n7883 & n7887;
  assign n7889 = n736 & ~n7888;
  assign n7890 = ~n7568 & ~n7822;
  assign n7891 = ~n7889 & n7890;
  assign n7892 = n7882 & n7891;
  assign n7893 = ~n7870 & n7892;
  assign n7894 = n1178 & ~n7893;
  assign n7895 = ~Pi25 & ~n7374;
  assign n7896 = n868 & ~n7797;
  assign n7897 = n950 & ~n7802;
  assign n7898 = ~n7896 & ~n7897;
  assign n7899 = n7384 & n7898;
  assign n7900 = ~n7895 & n7899;
  assign n7901 = n923 & ~n7900;
  assign n7902 = n949 & n7667;
  assign n7903 = n867 & n7671;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = Pi25 & ~n7904;
  assign n7906 = n7334 & ~n7905;
  assign n7907 = n736 & ~n7906;
  assign n7908 = ~n7901 & ~n7907;
  assign n7909 = n950 & ~n7794;
  assign n7910 = ~Pi25 & ~n7249;
  assign n7911 = n868 & ~n7791;
  assign n7912 = n7259 & ~n7911;
  assign n7913 = ~n7910 & n7912;
  assign n7914 = ~n7909 & n7913;
  assign n7915 = n738 & ~n7914;
  assign n7916 = Pi25 & ~n7675;
  assign n7917 = n6916 & ~n7916;
  assign n7918 = n1030 & ~n7917;
  assign n7919 = ~n7048 & ~n7918;
  assign n7920 = ~n7915 & n7919;
  assign n7921 = n7908 & n7920;
  assign n7922 = ~n7822 & n7921;
  assign n7923 = n1672 & ~n7922;
  assign n7924 = ~n7894 & ~n7923;
  assign n7925 = ~n7869 & n7924;
  assign n7926 = ~n7841 & n7925;
  assign n7927 = n863 & ~n7926;
  assign n7928 = ~n7814 & ~n7927;
  assign n7929 = ~n6885 & n7928;
  assign n1027 = n7666 | n7929;
  assign n7931 = ~P__cmxig_1 & n569;
  assign n7932 = P__cmxcl_1 & ~n7931;
  assign n7933 = Ni14 & ~n7932;
  assign n7934 = n568 & n604;
  assign n7935 = P__cmxcl_1 & ~n569;
  assign n7936 = ~n7934 & n7935;
  assign n7937 = ~Ni14 & n7936;
  assign n1032_1 = n7933 | n7937;
  assign n7939 = P__cmxcl_1 & n583;
  assign n7940 = Ni13 & ~n7939;
  assign n7941 = P__cmxig_1 & n571;
  assign n7942 = ~Pi27 & Ni12;
  assign n7943 = Ni11 & ~n677;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = P__cmxcl_1 & n678;
  assign n7946 = ~n7944 & n7945;
  assign n7947 = ~n7941 & ~n7946;
  assign n1037_1 = n7940 | ~n7947;
  assign n7949 = ~Ni12 & ~n7939;
  assign n7950 = Ni12 & n583;
  assign n7951 = P__cmxcl_1 & n7950;
  assign n7952 = ~n7949 & ~n7951;
  assign n1042 = ~n676 & n7952;
  assign n7954 = ~Ni11 & ~n7939;
  assign n7955 = n677 & n679;
  assign n7956 = Ni11 & n7950;
  assign n7957 = ~n582 & ~n7956;
  assign n7958 = ~n7955 & n7957;
  assign n7959 = P__cmxcl_1 & ~n7958;
  assign n1047_1 = ~n7954 & ~n7959;
  assign n7961 = ~Ni10 & ~P__cmxcl_1;
  assign n7962 = P__cmxcl_1 & n616;
  assign n7963 = ~Ni9 & ~n687;
  assign n7964 = Ni8 & ~n7963;
  assign n7965 = ~n577 & n578;
  assign n7966 = Ni10 & P__cmxcl_1;
  assign n7967 = ~Ni10 & ~Ni7;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = ~n7965 & ~n7968;
  assign n7970 = ~n7964 & n7969;
  assign n7971 = ~n7962 & ~n7970;
  assign n1052_1 = ~n7961 & n7971;
  assign n7973 = P__cmxig_0 & n578;
  assign n7974 = Ni7 & ~n691;
  assign n7975 = ~Pi24 & Ni8;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = ~n7973 & n7976;
  assign n7978 = n7966 & ~n7977;
  assign n7979 = ~Ni9 & ~n7978;
  assign n1057 = ~n7962 & ~n7979;
  assign n7981 = ~Ni8 & ~n7962;
  assign n7982 = Ni8 & P__cmxcl_1;
  assign n7983 = ~n616 & ~n689;
  assign n7984 = n7982 & ~n7983;
  assign n1062_1 = ~n7981 & ~n7984;
  assign n7986 = ~Ni7 & ~n7962;
  assign n7987 = n691 & n693;
  assign n7988 = Ni8 & Ni7;
  assign n7989 = n616 & n7988;
  assign n7990 = ~n578 & ~n7989;
  assign n7991 = ~n7987 & n7990;
  assign n7992 = P__cmxcl_1 & ~n7991;
  assign n1067_1 = ~n7986 & ~n7992;
  assign n7994 = n651 & n663;
  assign n7995 = Ni5 & ~Ni4;
  assign n7996 = Ni30 & n7995;
  assign n7997 = Ni31 & ~Ni2;
  assign n7998 = Ni3 & n7997;
  assign n7999 = ~n7996 & n7998;
  assign n8000 = n578 & ~n616;
  assign n8001 = ~n690 & ~n7987;
  assign n8002 = ~n8000 & n8001;
  assign n8003 = ~n855 & ~n8002;
  assign n8004 = ~Ni31 & n5370;
  assign n8005 = ~Pi26 & n3534;
  assign n8006 = ~n8004 & n8005;
  assign n8007 = Ni33 & ~n583;
  assign n8008 = ~Ni12 & n8007;
  assign n8009 = ~Ni31 & n3096;
  assign n8010 = ~n3122 & ~n8009;
  assign n8011 = n4046 & n8010;
  assign n8012 = ~n8008 & ~n8011;
  assign n8013 = ~n8006 & n8012;
  assign n8014 = ~Ni11 & ~n8013;
  assign n8015 = Ni30 & ~n652;
  assign n8016 = Ni33 & n681;
  assign n8017 = n8015 & ~n8016;
  assign n8018 = ~n8014 & n8017;
  assign n8019 = ~n8003 & n8018;
  assign n8020 = P__cmxcl_1 & n8019;
  assign n8021 = ~n7999 & ~n8020;
  assign n8022 = ~n7994 & n8021;
  assign n8023 = ~Ni6 & ~n8022;
  assign n8024 = Ni6 & ~n7997;
  assign n8025 = ~P__cmxcl_1 & ~n8024;
  assign n8026 = ~n8000 & n8015;
  assign n8027 = ~n8008 & n8026;
  assign n8028 = n582 & ~n583;
  assign n8029 = n855 & ~n8028;
  assign n8030 = Ni6 & ~n8029;
  assign n8031 = ~n8027 & n8030;
  assign n8032 = P__cmxcl_1 & ~n8031;
  assign n8033 = ~n8025 & ~n8032;
  assign n1072 = n8023 | n8033;
  assign n8035 = ~Ni14 & ~n855;
  assign n8036 = ~n672 & ~n8035;
  assign n8037 = n4427 & ~n8036;
  assign n8038 = ~n582 & ~n3087;
  assign n8039 = n677 & n855;
  assign n8040 = n680 & ~n8039;
  assign n8041 = n8038 & ~n8040;
  assign n8042 = ~n8037 & n8041;
  assign n8043 = Pi23 & ~n8042;
  assign n8044 = Pi26 & ~n8010;
  assign n8045 = n680 & ~n8044;
  assign n8046 = ~Pi26 & n8009;
  assign n8047 = n3534 & ~n8046;
  assign n8048 = ~n8045 & ~n8047;
  assign n8049 = ~n3122 & ~n8048;
  assign n8050 = ~n3122 & ~n8038;
  assign n8051 = Pi24 & ~n8042;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = ~n8049 & n8052;
  assign n8054 = ~n3141 & n4046;
  assign n8055 = n637 & n8004;
  assign n8056 = n8054 & ~n8055;
  assign n8057 = n8053 & ~n8056;
  assign n8058 = ~n8043 & n8057;
  assign n8059 = n4819 & ~n8058;
  assign n8060 = Ni14 & ~n3141;
  assign n8061 = Ni12 & n8060;
  assign n8062 = n8036 & n8038;
  assign n8063 = ~Ni12 & ~n8039;
  assign n8064 = n8062 & ~n8063;
  assign n8065 = ~n8061 & n8064;
  assign n8066 = ~Ni9 & ~n7988;
  assign n8067 = Ni10 & Ni7;
  assign n8068 = ~Ni8 & ~n8067;
  assign n8069 = n8066 & ~n8068;
  assign n8070 = ~n8065 & ~n8069;
  assign n8071 = n691 & n8004;
  assign n8072 = n8054 & ~n8071;
  assign n8073 = ~Pi23 & ~n8042;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = n8053 & n8074;
  assign n8076 = n694 & ~n8075;
  assign n8077 = ~n8070 & ~n8076;
  assign n8078 = n4046 & ~n8004;
  assign n8079 = Pi24 & ~n8050;
  assign n8080 = n8042 & ~n8054;
  assign n8081 = ~n8079 & ~n8080;
  assign n8082 = ~n8049 & ~n8081;
  assign n8083 = ~n8078 & n8082;
  assign n8084 = n4682 & ~n8083;
  assign n8085 = n8077 & ~n8084;
  assign n8086 = ~n8059 & n8085;
  assign n8087 = ~Ni6 & ~n8086;
  assign n8088 = ~n8031 & ~n8087;
  assign n8089 = Ni5 & ~n8088;
  assign n8090 = P__cmxcl_1 & n8089;
  assign n8091 = n650 & n652;
  assign n8092 = ~n8020 & ~n8091;
  assign n8093 = n660 & ~n8092;
  assign n8094 = Ni31 & Ni6;
  assign n8095 = n651 & ~n8094;
  assign n8096 = ~n656 & n8095;
  assign n8097 = Ni5 & n8094;
  assign n8098 = n664 & ~n8097;
  assign n8099 = ~Ni2 & ~n8098;
  assign n8100 = Ni5 & ~n8099;
  assign n8101 = ~n663 & n8098;
  assign n8102 = n8094 & n8101;
  assign n8103 = ~n8100 & ~n8102;
  assign n8104 = ~n8096 & n8103;
  assign n8105 = ~n8093 & n8104;
  assign n1077 = n8090 | ~n8105;
  assign n8107 = ~Ni5 & ~n8086;
  assign n8108 = ~n8089 & ~n8107;
  assign n8109 = Ni4 & ~n8108;
  assign n8110 = n7995 & n8019;
  assign n8111 = Ni6 & n8110;
  assign n8112 = ~n8109 & ~n8111;
  assign n8113 = P__cmxcl_1 & ~n8112;
  assign n8114 = n651 & n8094;
  assign n8115 = ~n660 & n8098;
  assign n8116 = Ni4 & Ni2;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = ~n8101 & n8117;
  assign n8119 = ~n8114 & n8118;
  assign n1082 = n8113 | ~n8119;
  assign P__cmx1ad_35 = 1'b0;
  assign P__cmx1ad_34 = 1'b0;
  assign P__cmx1ad_33 = 1'b0;
  assign P__cmx1ad_32 = 1'b0;
  assign P__cmx1ad_11 = 1'b0;
  assign P__cmx1ad_10 = 1'b0;
  assign P__cmx1ad_8 = 1'b0;
  assign P__cmx0ad_35 = 1'b0;
  assign P__cmx0ad_34 = 1'b0;
  assign P__cmx0ad_33 = 1'b0;
  assign P__cmx0ad_32 = 1'b0;
  assign P__cmx0ad_11 = 1'b0;
  assign P__cmx0ad_10 = 1'b0;
  assign P__cmx0ad_8 = 1'b0;
  assign P__cmxcl_0 = P__cmxcl_1;
  assign n1086 = P__cmxcl_1;
  always @ (posedge clock) begin
    Ni48 <= n932;
    Ni47 <= n937;
    Ni46 <= n942_1;
    Ni45 <= n947_1;
    Ni44 <= n952_1;
    Ni43 <= n957_1;
    Ni42 <= n962;
    Ni41 <= n967_1;
    Ni40 <= n972_1;
    Ni39 <= n977;
    Ni38 <= n982_1;
    Ni37 <= n987_1;
    Ni36 <= n992;
    Ni35 <= n997_1;
    Ni34 <= n1002;
    Ni33 <= n1007_1;
    Ni32 <= n1012;
    Ni31 <= n1017_1;
    Ni30 <= n1022_1;
    n18 <= n1027;
    Ni14 <= n1032_1;
    Ni13 <= n1037_1;
    Ni12 <= n1042;
    Ni11 <= n1047_1;
    Ni10 <= n1052_1;
    Ni9 <= n1057;
    Ni8 <= n1062_1;
    Ni7 <= n1067_1;
    Ni6 <= n1072;
    Ni5 <= n1077;
    Ni4 <= n1082;
    Ni3 <= n1086;
    Ni2 <= n1091_1;
  end
endmodule


