// Benchmark "ksa_128" written by ABC on Sat Apr 23 20:18:09 2016

module ksa_128 ( 
    a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7, a8, b8,
    a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15, b15,
    a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22, b22,
    a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29, b29,
    a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36, b36,
    a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43, b43,
    a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50, b50,
    a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57, b57,
    a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64, b64,
    a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71, b71,
    a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78, b78,
    a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85, b85,
    a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92, b92,
    a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99, b99,
    a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105, b105,
    a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111, b111,
    a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117, b117,
    a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123, b123,
    a124, b124, a125, b125, a126, b126, a127, b127,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128  );
  input  a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7,
    a8, b8, a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15,
    b15, a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22,
    b22, a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29,
    b29, a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36,
    b36, a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43,
    b43, a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50,
    b50, a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57,
    b57, a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64,
    b64, a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71,
    b71, a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78,
    b78, a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85,
    b85, a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92,
    b92, a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99,
    b99, a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105,
    b105, a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111,
    b111, a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117,
    b117, a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123,
    b123, a124, b124, a125, b125, a126, b126, a127, b127;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128;
  wire n386, n387, n389, n390, n391, n392, n393, n395, n396, n397, n398,
    n399, n400, n402, n403, n404, n405, n406, n407, n408, n409, n410, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424, n425,
    n426, n427, n428, n429, n431, n432, n433, n434, n435, n436, n437, n438,
    n439, n441, n442, n443, n444, n445, n446, n447, n448, n450, n451, n452,
    n453, n454, n455, n456, n457, n459, n460, n461, n462, n463, n464, n465,
    n466, n468, n469, n470, n471, n472, n473, n474, n475, n477, n478, n479,
    n480, n481, n482, n483, n484, n486, n487, n488, n489, n490, n491, n492,
    n493, n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506,
    n507, n508, n509, n510, n511, n513, n514, n515, n516, n517, n518, n519,
    n520, n522, n523, n524, n525, n526, n527, n528, n529, n531, n532, n533,
    n534, n535, n536, n537, n538, n540, n541, n542, n543, n544, n545, n546,
    n547, n549, n550, n551, n552, n553, n554, n555, n556, n558, n559, n560,
    n561, n562, n563, n564, n565, n567, n568, n569, n570, n571, n572, n573,
    n574, n576, n577, n578, n579, n580, n581, n582, n583, n585, n586, n587,
    n588, n589, n590, n591, n592, n594, n595, n596, n597, n598, n599, n600,
    n601, n603, n604, n605, n606, n607, n608, n609, n610, n612, n613, n614,
    n615, n616, n617, n618, n619, n621, n622, n623, n624, n625, n626, n627,
    n628, n630, n631, n632, n633, n634, n635, n636, n637, n639, n640, n641,
    n642, n643, n644, n645, n646, n648, n649, n650, n651, n652, n653, n654,
    n655, n657, n658, n659, n660, n661, n662, n663, n664, n666, n667, n668,
    n669, n670, n671, n672, n673, n675, n676, n677, n678, n679, n680, n681,
    n682, n684, n685, n686, n687, n688, n689, n690, n691, n693, n694, n695,
    n696, n697, n698, n699, n700, n702, n703, n704, n705, n706, n707, n708,
    n709, n711, n712, n713, n714, n715, n716, n717, n718, n720, n721, n722,
    n723, n724, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735,
    n736, n738, n739, n740, n741, n742, n743, n744, n745, n747, n748, n749,
    n750, n751, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762,
    n763, n765, n766, n767, n768, n769, n770, n771, n772, n774, n775, n776,
    n777, n778, n779, n780, n781, n783, n784, n785, n786, n787, n788, n789,
    n790, n792, n793, n794, n795, n796, n797, n798, n799, n801, n802, n803,
    n804, n805, n806, n807, n808, n810, n811, n812, n813, n814, n815, n816,
    n817, n819, n820, n821, n822, n823, n824, n825, n826, n828, n829, n830,
    n831, n832, n833, n834, n835, n837, n838, n839, n840, n841, n842, n843,
    n844, n846, n847, n848, n849, n850, n851, n852, n853, n855, n856, n857,
    n858, n859, n860, n861, n862, n864, n865, n866, n867, n868, n869, n870,
    n871, n873, n874, n875, n876, n877, n878, n879, n880, n882, n883, n884,
    n885, n886, n887, n888, n889, n891, n892, n893, n894, n895, n896, n897,
    n898, n900, n901, n902, n903, n904, n905, n906, n907, n909, n910, n911,
    n912, n913, n914, n915, n916, n918, n919, n920, n921, n922, n923, n924,
    n925, n927, n928, n929, n930, n931, n932, n933, n934, n936, n937, n938,
    n939, n940, n941, n942, n943, n945, n946, n947, n948, n949, n950, n951,
    n952, n954, n955, n956, n957, n958, n959, n960, n961, n963, n964, n965,
    n966, n967, n968, n969, n970, n972, n973, n974, n975, n976, n977, n978,
    n979, n981, n982, n983, n984, n985, n986, n987, n988, n990, n991, n992,
    n993, n994, n995, n996, n997, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1531, n1532, n1533,
    n1534;
  assign n386 = a0 & b0;
  assign n387 = ~a0 & ~b0;
  assign s0 = ~n386 & ~n387;
  assign n389 = a1 & b1;
  assign n390 = ~a1 & ~b1;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & n391;
  assign n393 = ~n386 & ~n391;
  assign s1 = ~n392 & ~n393;
  assign n395 = ~n389 & ~n392;
  assign n396 = a2 & b2;
  assign n397 = ~a2 & ~b2;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n395 & n398;
  assign n400 = n395 & ~n398;
  assign s2 = ~n399 & ~n400;
  assign n402 = n392 & n398;
  assign n403 = ~n389 & ~n396;
  assign n404 = ~n397 & ~n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = a3 & b3;
  assign n407 = ~a3 & ~b3;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n405 & n408;
  assign n410 = n405 & ~n408;
  assign s3 = ~n409 & ~n410;
  assign n412 = n399 & n408;
  assign n413 = ~n396 & ~n406;
  assign n414 = ~n407 & ~n413;
  assign n415 = ~n412 & ~n414;
  assign n416 = a4 & b4;
  assign n417 = ~a4 & ~b4;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n415 & n418;
  assign n420 = n415 & ~n418;
  assign s4 = ~n419 & ~n420;
  assign n422 = a5 & b5;
  assign n423 = ~a5 & ~b5;
  assign n424 = ~n422 & ~n423;
  assign n425 = ~n406 & ~n416;
  assign n426 = ~n409 & n425;
  assign n427 = ~n417 & ~n426;
  assign n428 = ~n424 & ~n427;
  assign n429 = n424 & n427;
  assign s5 = ~n428 & ~n429;
  assign n431 = n419 & n424;
  assign n432 = ~n416 & ~n422;
  assign n433 = ~n423 & ~n432;
  assign n434 = ~n431 & ~n433;
  assign n435 = a6 & b6;
  assign n436 = ~a6 & ~b6;
  assign n437 = ~n435 & ~n436;
  assign n438 = n434 & ~n437;
  assign n439 = ~n434 & n437;
  assign s6 = ~n438 & ~n439;
  assign n441 = a7 & b7;
  assign n442 = ~a7 & ~b7;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~n422 & ~n435;
  assign n445 = ~n429 & n444;
  assign n446 = ~n436 & ~n445;
  assign n447 = n443 & n446;
  assign n448 = ~n443 & ~n446;
  assign s7 = ~n447 & ~n448;
  assign n450 = a8 & b8;
  assign n451 = ~a8 & ~b8;
  assign n452 = ~n450 & ~n451;
  assign n453 = ~n435 & ~n441;
  assign n454 = ~n439 & n453;
  assign n455 = ~n442 & ~n454;
  assign n456 = ~n452 & ~n455;
  assign n457 = n452 & n455;
  assign s8 = ~n456 & ~n457;
  assign n459 = a9 & b9;
  assign n460 = ~a9 & ~b9;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n441 & ~n450;
  assign n463 = ~n447 & n462;
  assign n464 = ~n451 & ~n463;
  assign n465 = n461 & n464;
  assign n466 = ~n461 & ~n464;
  assign s9 = ~n465 & ~n466;
  assign n468 = a10 & b10;
  assign n469 = ~a10 & ~b10;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~n450 & ~n459;
  assign n472 = ~n457 & n471;
  assign n473 = ~n460 & ~n472;
  assign n474 = ~n470 & ~n473;
  assign n475 = n470 & n473;
  assign s10 = ~n474 & ~n475;
  assign n477 = a11 & b11;
  assign n478 = ~a11 & ~b11;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n459 & ~n468;
  assign n481 = ~n465 & n480;
  assign n482 = ~n469 & ~n481;
  assign n483 = ~n479 & ~n482;
  assign n484 = n479 & n482;
  assign s11 = ~n483 & ~n484;
  assign n486 = a12 & b12;
  assign n487 = ~a12 & ~b12;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n468 & ~n477;
  assign n490 = ~n475 & n489;
  assign n491 = ~n478 & ~n490;
  assign n492 = ~n488 & ~n491;
  assign n493 = n488 & n491;
  assign s12 = ~n492 & ~n493;
  assign n495 = a13 & b13;
  assign n496 = ~a13 & ~b13;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n477 & ~n486;
  assign n499 = ~n484 & n498;
  assign n500 = ~n487 & ~n499;
  assign n501 = ~n497 & ~n500;
  assign n502 = n497 & n500;
  assign s13 = ~n501 & ~n502;
  assign n504 = a14 & b14;
  assign n505 = ~a14 & ~b14;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~n486 & ~n495;
  assign n508 = ~n493 & n507;
  assign n509 = ~n496 & ~n508;
  assign n510 = ~n506 & ~n509;
  assign n511 = n506 & n509;
  assign s14 = ~n510 & ~n511;
  assign n513 = a15 & b15;
  assign n514 = ~a15 & ~b15;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n495 & ~n504;
  assign n517 = ~n502 & n516;
  assign n518 = ~n505 & ~n517;
  assign n519 = ~n515 & ~n518;
  assign n520 = n515 & n518;
  assign s15 = ~n519 & ~n520;
  assign n522 = a16 & b16;
  assign n523 = ~a16 & ~b16;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n504 & ~n513;
  assign n526 = ~n511 & n525;
  assign n527 = ~n514 & ~n526;
  assign n528 = ~n524 & ~n527;
  assign n529 = n524 & n527;
  assign s16 = ~n528 & ~n529;
  assign n531 = a17 & b17;
  assign n532 = ~a17 & ~b17;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n513 & ~n522;
  assign n535 = ~n520 & n534;
  assign n536 = ~n523 & ~n535;
  assign n537 = ~n533 & ~n536;
  assign n538 = n533 & n536;
  assign s17 = ~n537 & ~n538;
  assign n540 = a18 & b18;
  assign n541 = ~a18 & ~b18;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~n522 & ~n531;
  assign n544 = ~n529 & n543;
  assign n545 = ~n532 & ~n544;
  assign n546 = ~n542 & ~n545;
  assign n547 = n542 & n545;
  assign s18 = ~n546 & ~n547;
  assign n549 = a19 & b19;
  assign n550 = ~a19 & ~b19;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n531 & ~n540;
  assign n553 = ~n538 & n552;
  assign n554 = ~n541 & ~n553;
  assign n555 = ~n551 & ~n554;
  assign n556 = n551 & n554;
  assign s19 = ~n555 & ~n556;
  assign n558 = a20 & b20;
  assign n559 = ~a20 & ~b20;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n540 & ~n549;
  assign n562 = ~n547 & n561;
  assign n563 = ~n550 & ~n562;
  assign n564 = ~n560 & ~n563;
  assign n565 = n560 & n563;
  assign s20 = ~n564 & ~n565;
  assign n567 = a21 & b21;
  assign n568 = ~a21 & ~b21;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n549 & ~n558;
  assign n571 = ~n556 & n570;
  assign n572 = ~n559 & ~n571;
  assign n573 = ~n569 & ~n572;
  assign n574 = n569 & n572;
  assign s21 = ~n573 & ~n574;
  assign n576 = a22 & b22;
  assign n577 = ~a22 & ~b22;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~n558 & ~n567;
  assign n580 = ~n565 & n579;
  assign n581 = ~n568 & ~n580;
  assign n582 = ~n578 & ~n581;
  assign n583 = n578 & n581;
  assign s22 = ~n582 & ~n583;
  assign n585 = a23 & b23;
  assign n586 = ~a23 & ~b23;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n567 & ~n576;
  assign n589 = ~n574 & n588;
  assign n590 = ~n577 & ~n589;
  assign n591 = ~n587 & ~n590;
  assign n592 = n587 & n590;
  assign s23 = ~n591 & ~n592;
  assign n594 = a24 & b24;
  assign n595 = ~a24 & ~b24;
  assign n596 = ~n594 & ~n595;
  assign n597 = ~n576 & ~n585;
  assign n598 = ~n583 & n597;
  assign n599 = ~n586 & ~n598;
  assign n600 = ~n596 & ~n599;
  assign n601 = n596 & n599;
  assign s24 = ~n600 & ~n601;
  assign n603 = a25 & b25;
  assign n604 = ~a25 & ~b25;
  assign n605 = ~n603 & ~n604;
  assign n606 = ~n585 & ~n594;
  assign n607 = ~n592 & n606;
  assign n608 = ~n595 & ~n607;
  assign n609 = ~n605 & ~n608;
  assign n610 = n605 & n608;
  assign s25 = ~n609 & ~n610;
  assign n612 = a26 & b26;
  assign n613 = ~a26 & ~b26;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n594 & ~n603;
  assign n616 = ~n601 & n615;
  assign n617 = ~n604 & ~n616;
  assign n618 = ~n614 & ~n617;
  assign n619 = n614 & n617;
  assign s26 = ~n618 & ~n619;
  assign n621 = a27 & b27;
  assign n622 = ~a27 & ~b27;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n603 & ~n612;
  assign n625 = ~n610 & n624;
  assign n626 = ~n613 & ~n625;
  assign n627 = ~n623 & ~n626;
  assign n628 = n623 & n626;
  assign s27 = ~n627 & ~n628;
  assign n630 = a28 & b28;
  assign n631 = ~a28 & ~b28;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n612 & ~n621;
  assign n634 = ~n619 & n633;
  assign n635 = ~n622 & ~n634;
  assign n636 = ~n632 & ~n635;
  assign n637 = n632 & n635;
  assign s28 = ~n636 & ~n637;
  assign n639 = a29 & b29;
  assign n640 = ~a29 & ~b29;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n621 & ~n630;
  assign n643 = ~n628 & n642;
  assign n644 = ~n631 & ~n643;
  assign n645 = ~n641 & ~n644;
  assign n646 = n641 & n644;
  assign s29 = ~n645 & ~n646;
  assign n648 = a30 & b30;
  assign n649 = ~a30 & ~b30;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n630 & ~n639;
  assign n652 = ~n637 & n651;
  assign n653 = ~n640 & ~n652;
  assign n654 = ~n650 & ~n653;
  assign n655 = n650 & n653;
  assign s30 = ~n654 & ~n655;
  assign n657 = a31 & b31;
  assign n658 = ~a31 & ~b31;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n639 & ~n648;
  assign n661 = ~n646 & n660;
  assign n662 = ~n649 & ~n661;
  assign n663 = ~n659 & ~n662;
  assign n664 = n659 & n662;
  assign s31 = ~n663 & ~n664;
  assign n666 = a32 & b32;
  assign n667 = ~a32 & ~b32;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n648 & ~n657;
  assign n670 = ~n655 & n669;
  assign n671 = ~n658 & ~n670;
  assign n672 = ~n668 & ~n671;
  assign n673 = n668 & n671;
  assign s32 = ~n672 & ~n673;
  assign n675 = a33 & b33;
  assign n676 = ~a33 & ~b33;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n657 & ~n666;
  assign n679 = ~n664 & n678;
  assign n680 = ~n667 & ~n679;
  assign n681 = ~n677 & ~n680;
  assign n682 = n677 & n680;
  assign s33 = ~n681 & ~n682;
  assign n684 = a34 & b34;
  assign n685 = ~a34 & ~b34;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n666 & ~n675;
  assign n688 = ~n673 & n687;
  assign n689 = ~n676 & ~n688;
  assign n690 = ~n686 & ~n689;
  assign n691 = n686 & n689;
  assign s34 = ~n690 & ~n691;
  assign n693 = a35 & b35;
  assign n694 = ~a35 & ~b35;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~n675 & ~n684;
  assign n697 = ~n682 & n696;
  assign n698 = ~n685 & ~n697;
  assign n699 = ~n695 & ~n698;
  assign n700 = n695 & n698;
  assign s35 = ~n699 & ~n700;
  assign n702 = a36 & b36;
  assign n703 = ~a36 & ~b36;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~n684 & ~n693;
  assign n706 = ~n691 & n705;
  assign n707 = ~n694 & ~n706;
  assign n708 = ~n704 & ~n707;
  assign n709 = n704 & n707;
  assign s36 = ~n708 & ~n709;
  assign n711 = a37 & b37;
  assign n712 = ~a37 & ~b37;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n693 & ~n702;
  assign n715 = ~n700 & n714;
  assign n716 = ~n703 & ~n715;
  assign n717 = ~n713 & ~n716;
  assign n718 = n713 & n716;
  assign s37 = ~n717 & ~n718;
  assign n720 = a38 & b38;
  assign n721 = ~a38 & ~b38;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~n702 & ~n711;
  assign n724 = ~n709 & n723;
  assign n725 = ~n712 & ~n724;
  assign n726 = ~n722 & ~n725;
  assign n727 = n722 & n725;
  assign s38 = ~n726 & ~n727;
  assign n729 = a39 & b39;
  assign n730 = ~a39 & ~b39;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n711 & ~n720;
  assign n733 = ~n718 & n732;
  assign n734 = ~n721 & ~n733;
  assign n735 = ~n731 & ~n734;
  assign n736 = n731 & n734;
  assign s39 = ~n735 & ~n736;
  assign n738 = a40 & b40;
  assign n739 = ~a40 & ~b40;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n720 & ~n729;
  assign n742 = ~n727 & n741;
  assign n743 = ~n730 & ~n742;
  assign n744 = ~n740 & ~n743;
  assign n745 = n740 & n743;
  assign s40 = ~n744 & ~n745;
  assign n747 = a41 & b41;
  assign n748 = ~a41 & ~b41;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~n729 & ~n738;
  assign n751 = ~n736 & n750;
  assign n752 = ~n739 & ~n751;
  assign n753 = ~n749 & ~n752;
  assign n754 = n749 & n752;
  assign s41 = ~n753 & ~n754;
  assign n756 = a42 & b42;
  assign n757 = ~a42 & ~b42;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n738 & ~n747;
  assign n760 = ~n745 & n759;
  assign n761 = ~n748 & ~n760;
  assign n762 = ~n758 & ~n761;
  assign n763 = n758 & n761;
  assign s42 = ~n762 & ~n763;
  assign n765 = a43 & b43;
  assign n766 = ~a43 & ~b43;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n747 & ~n756;
  assign n769 = ~n754 & n768;
  assign n770 = ~n757 & ~n769;
  assign n771 = ~n767 & ~n770;
  assign n772 = n767 & n770;
  assign s43 = ~n771 & ~n772;
  assign n774 = a44 & b44;
  assign n775 = ~a44 & ~b44;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n756 & ~n765;
  assign n778 = ~n763 & n777;
  assign n779 = ~n766 & ~n778;
  assign n780 = ~n776 & ~n779;
  assign n781 = n776 & n779;
  assign s44 = ~n780 & ~n781;
  assign n783 = a45 & b45;
  assign n784 = ~a45 & ~b45;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n765 & ~n774;
  assign n787 = ~n772 & n786;
  assign n788 = ~n775 & ~n787;
  assign n789 = ~n785 & ~n788;
  assign n790 = n785 & n788;
  assign s45 = ~n789 & ~n790;
  assign n792 = a46 & b46;
  assign n793 = ~a46 & ~b46;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n774 & ~n783;
  assign n796 = ~n781 & n795;
  assign n797 = ~n784 & ~n796;
  assign n798 = ~n794 & ~n797;
  assign n799 = n794 & n797;
  assign s46 = ~n798 & ~n799;
  assign n801 = a47 & b47;
  assign n802 = ~a47 & ~b47;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n783 & ~n792;
  assign n805 = ~n790 & n804;
  assign n806 = ~n793 & ~n805;
  assign n807 = ~n803 & ~n806;
  assign n808 = n803 & n806;
  assign s47 = ~n807 & ~n808;
  assign n810 = a48 & b48;
  assign n811 = ~a48 & ~b48;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n792 & ~n801;
  assign n814 = ~n799 & n813;
  assign n815 = ~n802 & ~n814;
  assign n816 = ~n812 & ~n815;
  assign n817 = n812 & n815;
  assign s48 = ~n816 & ~n817;
  assign n819 = a49 & b49;
  assign n820 = ~a49 & ~b49;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n801 & ~n810;
  assign n823 = ~n808 & n822;
  assign n824 = ~n811 & ~n823;
  assign n825 = ~n821 & ~n824;
  assign n826 = n821 & n824;
  assign s49 = ~n825 & ~n826;
  assign n828 = a50 & b50;
  assign n829 = ~a50 & ~b50;
  assign n830 = ~n828 & ~n829;
  assign n831 = ~n810 & ~n819;
  assign n832 = ~n817 & n831;
  assign n833 = ~n820 & ~n832;
  assign n834 = ~n830 & ~n833;
  assign n835 = n830 & n833;
  assign s50 = ~n834 & ~n835;
  assign n837 = a51 & b51;
  assign n838 = ~a51 & ~b51;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n819 & ~n828;
  assign n841 = ~n826 & n840;
  assign n842 = ~n829 & ~n841;
  assign n843 = ~n839 & ~n842;
  assign n844 = n839 & n842;
  assign s51 = ~n843 & ~n844;
  assign n846 = a52 & b52;
  assign n847 = ~a52 & ~b52;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n828 & ~n837;
  assign n850 = ~n835 & n849;
  assign n851 = ~n838 & ~n850;
  assign n852 = ~n848 & ~n851;
  assign n853 = n848 & n851;
  assign s52 = ~n852 & ~n853;
  assign n855 = a53 & b53;
  assign n856 = ~a53 & ~b53;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n837 & ~n846;
  assign n859 = ~n844 & n858;
  assign n860 = ~n847 & ~n859;
  assign n861 = ~n857 & ~n860;
  assign n862 = n857 & n860;
  assign s53 = ~n861 & ~n862;
  assign n864 = a54 & b54;
  assign n865 = ~a54 & ~b54;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n846 & ~n855;
  assign n868 = ~n853 & n867;
  assign n869 = ~n856 & ~n868;
  assign n870 = ~n866 & ~n869;
  assign n871 = n866 & n869;
  assign s54 = ~n870 & ~n871;
  assign n873 = a55 & b55;
  assign n874 = ~a55 & ~b55;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~n855 & ~n864;
  assign n877 = ~n862 & n876;
  assign n878 = ~n865 & ~n877;
  assign n879 = ~n875 & ~n878;
  assign n880 = n875 & n878;
  assign s55 = ~n879 & ~n880;
  assign n882 = a56 & b56;
  assign n883 = ~a56 & ~b56;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n864 & ~n873;
  assign n886 = ~n871 & n885;
  assign n887 = ~n874 & ~n886;
  assign n888 = ~n884 & ~n887;
  assign n889 = n884 & n887;
  assign s56 = ~n888 & ~n889;
  assign n891 = a57 & b57;
  assign n892 = ~a57 & ~b57;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n873 & ~n882;
  assign n895 = ~n880 & n894;
  assign n896 = ~n883 & ~n895;
  assign n897 = ~n893 & ~n896;
  assign n898 = n893 & n896;
  assign s57 = ~n897 & ~n898;
  assign n900 = a58 & b58;
  assign n901 = ~a58 & ~b58;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n882 & ~n891;
  assign n904 = ~n889 & n903;
  assign n905 = ~n892 & ~n904;
  assign n906 = ~n902 & ~n905;
  assign n907 = n902 & n905;
  assign s58 = ~n906 & ~n907;
  assign n909 = a59 & b59;
  assign n910 = ~a59 & ~b59;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n891 & ~n900;
  assign n913 = ~n898 & n912;
  assign n914 = ~n901 & ~n913;
  assign n915 = ~n911 & ~n914;
  assign n916 = n911 & n914;
  assign s59 = ~n915 & ~n916;
  assign n918 = a60 & b60;
  assign n919 = ~a60 & ~b60;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n900 & ~n909;
  assign n922 = ~n907 & n921;
  assign n923 = ~n910 & ~n922;
  assign n924 = ~n920 & ~n923;
  assign n925 = n920 & n923;
  assign s60 = ~n924 & ~n925;
  assign n927 = a61 & b61;
  assign n928 = ~a61 & ~b61;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n909 & ~n918;
  assign n931 = ~n916 & n930;
  assign n932 = ~n919 & ~n931;
  assign n933 = ~n929 & ~n932;
  assign n934 = n929 & n932;
  assign s61 = ~n933 & ~n934;
  assign n936 = a62 & b62;
  assign n937 = ~a62 & ~b62;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n918 & ~n927;
  assign n940 = ~n925 & n939;
  assign n941 = ~n928 & ~n940;
  assign n942 = ~n938 & ~n941;
  assign n943 = n938 & n941;
  assign s62 = ~n942 & ~n943;
  assign n945 = a63 & b63;
  assign n946 = ~a63 & ~b63;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~n927 & ~n936;
  assign n949 = ~n934 & n948;
  assign n950 = ~n937 & ~n949;
  assign n951 = ~n947 & ~n950;
  assign n952 = n947 & n950;
  assign s63 = ~n951 & ~n952;
  assign n954 = a64 & b64;
  assign n955 = ~a64 & ~b64;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n936 & ~n945;
  assign n958 = ~n943 & n957;
  assign n959 = ~n946 & ~n958;
  assign n960 = ~n956 & ~n959;
  assign n961 = n956 & n959;
  assign s64 = ~n960 & ~n961;
  assign n963 = a65 & b65;
  assign n964 = ~a65 & ~b65;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n945 & ~n954;
  assign n967 = ~n952 & n966;
  assign n968 = ~n955 & ~n967;
  assign n969 = ~n965 & ~n968;
  assign n970 = n965 & n968;
  assign s65 = ~n969 & ~n970;
  assign n972 = a66 & b66;
  assign n973 = ~a66 & ~b66;
  assign n974 = ~n972 & ~n973;
  assign n975 = ~n954 & ~n963;
  assign n976 = ~n961 & n975;
  assign n977 = ~n964 & ~n976;
  assign n978 = ~n974 & ~n977;
  assign n979 = n974 & n977;
  assign s66 = ~n978 & ~n979;
  assign n981 = a67 & b67;
  assign n982 = ~a67 & ~b67;
  assign n983 = ~n981 & ~n982;
  assign n984 = ~n963 & ~n972;
  assign n985 = ~n970 & n984;
  assign n986 = ~n973 & ~n985;
  assign n987 = ~n983 & ~n986;
  assign n988 = n983 & n986;
  assign s67 = ~n987 & ~n988;
  assign n990 = a68 & b68;
  assign n991 = ~a68 & ~b68;
  assign n992 = ~n990 & ~n991;
  assign n993 = ~n972 & ~n981;
  assign n994 = ~n979 & n993;
  assign n995 = ~n982 & ~n994;
  assign n996 = n992 & n995;
  assign n997 = ~n992 & ~n995;
  assign s68 = ~n996 & ~n997;
  assign n999 = a69 & b69;
  assign n1000 = ~a69 & ~b69;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~n981 & ~n990;
  assign n1003 = ~n988 & n1002;
  assign n1004 = ~n991 & ~n1003;
  assign n1005 = n1001 & n1004;
  assign n1006 = ~n1001 & ~n1004;
  assign s69 = ~n1005 & ~n1006;
  assign n1008 = a70 & b70;
  assign n1009 = ~a70 & ~b70;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = ~n990 & ~n999;
  assign n1012 = ~n996 & n1011;
  assign n1013 = ~n1000 & ~n1012;
  assign n1014 = n1010 & n1013;
  assign n1015 = ~n1010 & ~n1013;
  assign s70 = ~n1014 & ~n1015;
  assign n1017 = a71 & b71;
  assign n1018 = ~a71 & ~b71;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = ~n999 & ~n1008;
  assign n1021 = ~n1005 & n1020;
  assign n1022 = ~n1009 & ~n1021;
  assign n1023 = ~n1019 & ~n1022;
  assign n1024 = n1019 & n1022;
  assign s71 = ~n1023 & ~n1024;
  assign n1026 = a72 & b72;
  assign n1027 = ~a72 & ~b72;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1008 & ~n1017;
  assign n1030 = ~n1014 & n1029;
  assign n1031 = ~n1018 & ~n1030;
  assign n1032 = n1028 & n1031;
  assign n1033 = ~n1028 & ~n1031;
  assign s72 = ~n1032 & ~n1033;
  assign n1035 = a73 & b73;
  assign n1036 = ~a73 & ~b73;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = ~n1017 & ~n1026;
  assign n1039 = ~n1024 & n1038;
  assign n1040 = ~n1027 & ~n1039;
  assign n1041 = n1037 & n1040;
  assign n1042 = ~n1037 & ~n1040;
  assign s73 = ~n1041 & ~n1042;
  assign n1044 = a74 & b74;
  assign n1045 = ~a74 & ~b74;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = ~n1026 & ~n1035;
  assign n1048 = ~n1032 & n1047;
  assign n1049 = ~n1036 & ~n1048;
  assign n1050 = n1046 & n1049;
  assign n1051 = ~n1046 & ~n1049;
  assign s74 = ~n1050 & ~n1051;
  assign n1053 = a75 & b75;
  assign n1054 = ~a75 & ~b75;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1035 & ~n1044;
  assign n1057 = ~n1041 & n1056;
  assign n1058 = ~n1045 & ~n1057;
  assign n1059 = n1055 & n1058;
  assign n1060 = ~n1055 & ~n1058;
  assign s75 = ~n1059 & ~n1060;
  assign n1062 = a76 & b76;
  assign n1063 = ~a76 & ~b76;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n1044 & ~n1053;
  assign n1066 = ~n1050 & n1065;
  assign n1067 = ~n1054 & ~n1066;
  assign n1068 = ~n1064 & ~n1067;
  assign n1069 = n1064 & n1067;
  assign s76 = ~n1068 & ~n1069;
  assign n1071 = a77 & b77;
  assign n1072 = ~a77 & ~b77;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = ~n1053 & ~n1062;
  assign n1075 = ~n1059 & n1074;
  assign n1076 = ~n1063 & ~n1075;
  assign n1077 = ~n1073 & ~n1076;
  assign n1078 = n1073 & n1076;
  assign s77 = ~n1077 & ~n1078;
  assign n1080 = a78 & b78;
  assign n1081 = ~a78 & ~b78;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = ~n1062 & ~n1071;
  assign n1084 = ~n1069 & n1083;
  assign n1085 = ~n1072 & ~n1084;
  assign n1086 = ~n1082 & ~n1085;
  assign n1087 = n1082 & n1085;
  assign s78 = ~n1086 & ~n1087;
  assign n1089 = a79 & b79;
  assign n1090 = ~a79 & ~b79;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n1071 & ~n1080;
  assign n1093 = ~n1078 & n1092;
  assign n1094 = ~n1081 & ~n1093;
  assign n1095 = ~n1091 & ~n1094;
  assign n1096 = n1091 & n1094;
  assign s79 = ~n1095 & ~n1096;
  assign n1098 = a80 & b80;
  assign n1099 = ~a80 & ~b80;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n1080 & ~n1089;
  assign n1102 = ~n1087 & n1101;
  assign n1103 = ~n1090 & ~n1102;
  assign n1104 = n1100 & n1103;
  assign n1105 = ~n1100 & ~n1103;
  assign s80 = ~n1104 & ~n1105;
  assign n1107 = a81 & b81;
  assign n1108 = ~a81 & ~b81;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~n1089 & ~n1098;
  assign n1111 = ~n1096 & n1110;
  assign n1112 = ~n1099 & ~n1111;
  assign n1113 = n1109 & n1112;
  assign n1114 = ~n1109 & ~n1112;
  assign s81 = ~n1113 & ~n1114;
  assign n1116 = a82 & b82;
  assign n1117 = ~a82 & ~b82;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1098 & ~n1107;
  assign n1120 = ~n1104 & n1119;
  assign n1121 = ~n1108 & ~n1120;
  assign n1122 = n1118 & n1121;
  assign n1123 = ~n1118 & ~n1121;
  assign s82 = ~n1122 & ~n1123;
  assign n1125 = a83 & b83;
  assign n1126 = ~a83 & ~b83;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1107 & ~n1116;
  assign n1129 = ~n1113 & n1128;
  assign n1130 = ~n1117 & ~n1129;
  assign n1131 = n1127 & n1130;
  assign n1132 = ~n1127 & ~n1130;
  assign s83 = ~n1131 & ~n1132;
  assign n1134 = a84 & b84;
  assign n1135 = ~a84 & ~b84;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = ~n1116 & ~n1125;
  assign n1138 = ~n1122 & n1137;
  assign n1139 = ~n1126 & ~n1138;
  assign n1140 = n1136 & n1139;
  assign n1141 = ~n1136 & ~n1139;
  assign s84 = ~n1140 & ~n1141;
  assign n1143 = a85 & b85;
  assign n1144 = ~a85 & ~b85;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = ~n1125 & ~n1134;
  assign n1147 = ~n1131 & n1146;
  assign n1148 = ~n1135 & ~n1147;
  assign n1149 = n1145 & n1148;
  assign n1150 = ~n1145 & ~n1148;
  assign s85 = ~n1149 & ~n1150;
  assign n1152 = a86 & b86;
  assign n1153 = ~a86 & ~b86;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = ~n1134 & ~n1143;
  assign n1156 = ~n1140 & n1155;
  assign n1157 = ~n1144 & ~n1156;
  assign n1158 = n1154 & n1157;
  assign n1159 = ~n1154 & ~n1157;
  assign s86 = ~n1158 & ~n1159;
  assign n1161 = a87 & b87;
  assign n1162 = ~a87 & ~b87;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1143 & ~n1152;
  assign n1165 = ~n1149 & n1164;
  assign n1166 = ~n1153 & ~n1165;
  assign n1167 = n1163 & n1166;
  assign n1168 = ~n1163 & ~n1166;
  assign s87 = ~n1167 & ~n1168;
  assign n1170 = a88 & b88;
  assign n1171 = ~a88 & ~b88;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1152 & ~n1161;
  assign n1174 = ~n1158 & n1173;
  assign n1175 = ~n1162 & ~n1174;
  assign n1176 = n1172 & n1175;
  assign n1177 = ~n1172 & ~n1175;
  assign s88 = ~n1176 & ~n1177;
  assign n1179 = a89 & b89;
  assign n1180 = ~a89 & ~b89;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1161 & ~n1170;
  assign n1183 = ~n1167 & n1182;
  assign n1184 = ~n1171 & ~n1183;
  assign n1185 = n1181 & n1184;
  assign n1186 = ~n1181 & ~n1184;
  assign s89 = ~n1185 & ~n1186;
  assign n1188 = a90 & b90;
  assign n1189 = ~a90 & ~b90;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = ~n1170 & ~n1179;
  assign n1192 = ~n1176 & n1191;
  assign n1193 = ~n1180 & ~n1192;
  assign n1194 = n1190 & n1193;
  assign n1195 = ~n1190 & ~n1193;
  assign s90 = ~n1194 & ~n1195;
  assign n1197 = a91 & b91;
  assign n1198 = ~a91 & ~b91;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~n1179 & ~n1188;
  assign n1201 = ~n1185 & n1200;
  assign n1202 = ~n1189 & ~n1201;
  assign n1203 = n1199 & n1202;
  assign n1204 = ~n1199 & ~n1202;
  assign s91 = ~n1203 & ~n1204;
  assign n1206 = a92 & b92;
  assign n1207 = ~a92 & ~b92;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = ~n1188 & ~n1197;
  assign n1210 = ~n1194 & n1209;
  assign n1211 = ~n1198 & ~n1210;
  assign n1212 = n1208 & n1211;
  assign n1213 = ~n1208 & ~n1211;
  assign s92 = ~n1212 & ~n1213;
  assign n1215 = a93 & b93;
  assign n1216 = ~a93 & ~b93;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~n1197 & ~n1206;
  assign n1219 = ~n1203 & n1218;
  assign n1220 = ~n1207 & ~n1219;
  assign n1221 = n1217 & n1220;
  assign n1222 = ~n1217 & ~n1220;
  assign s93 = ~n1221 & ~n1222;
  assign n1224 = a94 & b94;
  assign n1225 = ~a94 & ~b94;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~n1206 & ~n1215;
  assign n1228 = ~n1212 & n1227;
  assign n1229 = ~n1216 & ~n1228;
  assign n1230 = n1226 & n1229;
  assign n1231 = ~n1226 & ~n1229;
  assign s94 = ~n1230 & ~n1231;
  assign n1233 = a95 & b95;
  assign n1234 = ~a95 & ~b95;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1215 & ~n1224;
  assign n1237 = ~n1221 & n1236;
  assign n1238 = ~n1225 & ~n1237;
  assign n1239 = n1235 & n1238;
  assign n1240 = ~n1235 & ~n1238;
  assign s95 = ~n1239 & ~n1240;
  assign n1242 = a96 & b96;
  assign n1243 = ~a96 & ~b96;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1224 & ~n1233;
  assign n1246 = ~n1230 & n1245;
  assign n1247 = ~n1234 & ~n1246;
  assign n1248 = n1244 & n1247;
  assign n1249 = ~n1244 & ~n1247;
  assign s96 = ~n1248 & ~n1249;
  assign n1251 = a97 & b97;
  assign n1252 = ~a97 & ~b97;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1233 & ~n1242;
  assign n1255 = ~n1239 & n1254;
  assign n1256 = ~n1243 & ~n1255;
  assign n1257 = n1253 & n1256;
  assign n1258 = ~n1253 & ~n1256;
  assign s97 = ~n1257 & ~n1258;
  assign n1260 = a98 & b98;
  assign n1261 = ~a98 & ~b98;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~n1242 & ~n1251;
  assign n1264 = ~n1248 & n1263;
  assign n1265 = ~n1252 & ~n1264;
  assign n1266 = n1262 & n1265;
  assign n1267 = ~n1262 & ~n1265;
  assign s98 = ~n1266 & ~n1267;
  assign n1269 = a99 & b99;
  assign n1270 = ~a99 & ~b99;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~n1251 & ~n1260;
  assign n1273 = ~n1257 & n1272;
  assign n1274 = ~n1261 & ~n1273;
  assign n1275 = n1271 & n1274;
  assign n1276 = ~n1271 & ~n1274;
  assign s99 = ~n1275 & ~n1276;
  assign n1278 = a100 & b100;
  assign n1279 = ~a100 & ~b100;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~n1260 & ~n1269;
  assign n1282 = ~n1266 & n1281;
  assign n1283 = ~n1270 & ~n1282;
  assign n1284 = n1280 & n1283;
  assign n1285 = ~n1280 & ~n1283;
  assign s100 = ~n1284 & ~n1285;
  assign n1287 = a101 & b101;
  assign n1288 = ~a101 & ~b101;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~n1269 & ~n1278;
  assign n1291 = ~n1275 & n1290;
  assign n1292 = ~n1279 & ~n1291;
  assign n1293 = n1289 & n1292;
  assign n1294 = ~n1289 & ~n1292;
  assign s101 = ~n1293 & ~n1294;
  assign n1296 = a102 & b102;
  assign n1297 = ~a102 & ~b102;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1278 & ~n1287;
  assign n1300 = ~n1284 & n1299;
  assign n1301 = ~n1288 & ~n1300;
  assign n1302 = n1298 & n1301;
  assign n1303 = ~n1298 & ~n1301;
  assign s102 = ~n1302 & ~n1303;
  assign n1305 = a103 & b103;
  assign n1306 = ~a103 & ~b103;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1287 & ~n1296;
  assign n1309 = ~n1293 & n1308;
  assign n1310 = ~n1297 & ~n1309;
  assign n1311 = n1307 & n1310;
  assign n1312 = ~n1307 & ~n1310;
  assign s103 = ~n1311 & ~n1312;
  assign n1314 = a104 & b104;
  assign n1315 = ~a104 & ~b104;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = ~n1296 & ~n1305;
  assign n1318 = ~n1302 & n1317;
  assign n1319 = ~n1306 & ~n1318;
  assign n1320 = n1316 & n1319;
  assign n1321 = ~n1316 & ~n1319;
  assign s104 = ~n1320 & ~n1321;
  assign n1323 = a105 & b105;
  assign n1324 = ~a105 & ~b105;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = ~n1305 & ~n1314;
  assign n1327 = ~n1311 & n1326;
  assign n1328 = ~n1315 & ~n1327;
  assign n1329 = n1325 & n1328;
  assign n1330 = ~n1325 & ~n1328;
  assign s105 = ~n1329 & ~n1330;
  assign n1332 = a106 & b106;
  assign n1333 = ~a106 & ~b106;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1314 & ~n1323;
  assign n1336 = ~n1320 & n1335;
  assign n1337 = ~n1324 & ~n1336;
  assign n1338 = n1334 & n1337;
  assign n1339 = ~n1334 & ~n1337;
  assign s106 = ~n1338 & ~n1339;
  assign n1341 = a107 & b107;
  assign n1342 = ~a107 & ~b107;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1323 & ~n1332;
  assign n1345 = ~n1329 & n1344;
  assign n1346 = ~n1333 & ~n1345;
  assign n1347 = ~n1343 & ~n1346;
  assign n1348 = n1343 & n1346;
  assign s107 = ~n1347 & ~n1348;
  assign n1350 = a108 & b108;
  assign n1351 = ~a108 & ~b108;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~n1332 & ~n1341;
  assign n1354 = ~n1338 & n1353;
  assign n1355 = ~n1342 & ~n1354;
  assign n1356 = n1352 & n1355;
  assign n1357 = ~n1352 & ~n1355;
  assign s108 = ~n1356 & ~n1357;
  assign n1359 = a109 & b109;
  assign n1360 = ~a109 & ~b109;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = ~n1341 & ~n1350;
  assign n1363 = ~n1348 & n1362;
  assign n1364 = ~n1351 & ~n1363;
  assign n1365 = n1361 & n1364;
  assign n1366 = ~n1361 & ~n1364;
  assign s109 = ~n1365 & ~n1366;
  assign n1368 = a110 & b110;
  assign n1369 = ~a110 & ~b110;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1350 & ~n1359;
  assign n1372 = ~n1356 & n1371;
  assign n1373 = ~n1360 & ~n1372;
  assign n1374 = n1370 & n1373;
  assign n1375 = ~n1370 & ~n1373;
  assign s110 = ~n1374 & ~n1375;
  assign n1377 = a111 & b111;
  assign n1378 = ~a111 & ~b111;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = ~n1359 & ~n1368;
  assign n1381 = ~n1365 & n1380;
  assign n1382 = ~n1369 & ~n1381;
  assign n1383 = ~n1379 & ~n1382;
  assign n1384 = n1379 & n1382;
  assign s111 = ~n1383 & ~n1384;
  assign n1386 = a112 & b112;
  assign n1387 = ~a112 & ~b112;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~n1368 & ~n1377;
  assign n1390 = ~n1374 & n1389;
  assign n1391 = ~n1378 & ~n1390;
  assign n1392 = n1388 & n1391;
  assign n1393 = ~n1388 & ~n1391;
  assign s112 = ~n1392 & ~n1393;
  assign n1395 = a113 & b113;
  assign n1396 = ~a113 & ~b113;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1377 & ~n1386;
  assign n1399 = ~n1384 & n1398;
  assign n1400 = ~n1387 & ~n1399;
  assign n1401 = ~n1397 & ~n1400;
  assign n1402 = n1397 & n1400;
  assign s113 = ~n1401 & ~n1402;
  assign n1404 = a114 & b114;
  assign n1405 = ~a114 & ~b114;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1386 & ~n1395;
  assign n1408 = ~n1392 & n1407;
  assign n1409 = ~n1396 & ~n1408;
  assign n1410 = ~n1406 & ~n1409;
  assign n1411 = n1406 & n1409;
  assign s114 = ~n1410 & ~n1411;
  assign n1413 = a115 & b115;
  assign n1414 = ~a115 & ~b115;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~n1395 & ~n1404;
  assign n1417 = ~n1402 & n1416;
  assign n1418 = ~n1405 & ~n1417;
  assign n1419 = ~n1415 & ~n1418;
  assign n1420 = n1415 & n1418;
  assign s115 = ~n1419 & ~n1420;
  assign n1422 = a116 & b116;
  assign n1423 = ~a116 & ~b116;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1404 & ~n1413;
  assign n1426 = ~n1411 & n1425;
  assign n1427 = ~n1414 & ~n1426;
  assign n1428 = ~n1424 & ~n1427;
  assign n1429 = n1424 & n1427;
  assign s116 = ~n1428 & ~n1429;
  assign n1431 = a117 & b117;
  assign n1432 = ~a117 & ~b117;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1413 & ~n1422;
  assign n1435 = ~n1420 & n1434;
  assign n1436 = ~n1423 & ~n1435;
  assign n1437 = n1433 & n1436;
  assign n1438 = ~n1433 & ~n1436;
  assign s117 = ~n1437 & ~n1438;
  assign n1440 = a118 & b118;
  assign n1441 = ~a118 & ~b118;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = ~n1422 & ~n1431;
  assign n1444 = ~n1429 & n1443;
  assign n1445 = ~n1432 & ~n1444;
  assign n1446 = ~n1442 & ~n1445;
  assign n1447 = n1442 & n1445;
  assign s118 = ~n1446 & ~n1447;
  assign n1449 = a119 & b119;
  assign n1450 = ~a119 & ~b119;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = ~n1431 & ~n1440;
  assign n1453 = ~n1437 & n1452;
  assign n1454 = ~n1441 & ~n1453;
  assign n1455 = ~n1451 & ~n1454;
  assign n1456 = n1451 & n1454;
  assign s119 = ~n1455 & ~n1456;
  assign n1458 = a120 & b120;
  assign n1459 = ~a120 & ~b120;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = ~n1440 & ~n1449;
  assign n1462 = ~n1447 & n1461;
  assign n1463 = ~n1450 & ~n1462;
  assign n1464 = ~n1460 & ~n1463;
  assign n1465 = n1460 & n1463;
  assign s120 = ~n1464 & ~n1465;
  assign n1467 = a121 & b121;
  assign n1468 = ~a121 & ~b121;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n1449 & ~n1458;
  assign n1471 = ~n1456 & n1470;
  assign n1472 = ~n1459 & ~n1471;
  assign n1473 = ~n1469 & ~n1472;
  assign n1474 = n1469 & n1472;
  assign s121 = ~n1473 & ~n1474;
  assign n1476 = a122 & b122;
  assign n1477 = ~a122 & ~b122;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = ~n1458 & ~n1467;
  assign n1480 = ~n1465 & n1479;
  assign n1481 = ~n1468 & ~n1480;
  assign n1482 = n1478 & n1481;
  assign n1483 = ~n1478 & ~n1481;
  assign s122 = ~n1482 & ~n1483;
  assign n1485 = a123 & b123;
  assign n1486 = ~a123 & ~b123;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~n1467 & ~n1476;
  assign n1489 = ~n1474 & n1488;
  assign n1490 = ~n1477 & ~n1489;
  assign n1491 = n1487 & n1490;
  assign n1492 = ~n1487 & ~n1490;
  assign s123 = ~n1491 & ~n1492;
  assign n1494 = a124 & b124;
  assign n1495 = ~a124 & ~b124;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1476 & ~n1485;
  assign n1498 = ~n1482 & n1497;
  assign n1499 = ~n1486 & ~n1498;
  assign n1500 = n1496 & n1499;
  assign n1501 = ~n1496 & ~n1499;
  assign s124 = ~n1500 & ~n1501;
  assign n1503 = a125 & b125;
  assign n1504 = ~a125 & ~b125;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1485 & ~n1494;
  assign n1507 = ~n1491 & n1506;
  assign n1508 = ~n1495 & ~n1507;
  assign n1509 = n1505 & n1508;
  assign n1510 = ~n1505 & ~n1508;
  assign s125 = ~n1509 & ~n1510;
  assign n1512 = n1494 & ~n1504;
  assign n1513 = n1500 & n1505;
  assign n1514 = ~n1503 & ~n1513;
  assign n1515 = ~n1512 & n1514;
  assign n1516 = a126 & b126;
  assign n1517 = ~a126 & ~b126;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1515 & ~n1518;
  assign n1520 = n1515 & n1518;
  assign s126 = n1519 | n1520;
  assign n1522 = a127 & b127;
  assign n1523 = ~a127 & ~b127;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1503 & ~n1516;
  assign n1526 = ~n1509 & n1525;
  assign n1527 = ~n1517 & ~n1526;
  assign n1528 = ~n1524 & n1527;
  assign n1529 = n1524 & ~n1527;
  assign s127 = n1528 | n1529;
  assign n1531 = ~n1512 & n1525;
  assign n1532 = ~n1513 & n1531;
  assign n1533 = ~n1523 & ~n1532;
  assign n1534 = ~n1517 & n1533;
  assign s128 = n1522 | n1534;
endmodule


