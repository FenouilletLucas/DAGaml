// Benchmark "pair" written by ABC on Tue May 16 16:07:51 2017

module pair ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, c0, c1, c2, c3, c4,
    c5, d0, d1, d2, d3, d4, d5, e0, e1, e2, e3, e4, e5, f0, f1, f2, f3, f4,
    f5, g0, g1, g2, g3, g4, g5, h0, h1, h2, h3, h4, h5, i0, i1, i2, i3, i4,
    i5, j0, j1, j2, j3, j4, j5, k0, k1, k2, k3, k4, k5, l0, l1, l2, l3, l4,
    l5, m0, m1, m2, m3, m4, m5, n0, n1, n2, n3, n4, n5, o0, o1, o2, o3, o4,
    o5, p0, p1, p2, p3, p4, p5, q0, q1, q2, q3, q4, q5, r0, r1, r2, r3, r4,
    r5, s0, s1, s2, s3, s4, t0, t1, t2, t3, t4, u0, u1, u2, u3, u4, v0, v1,
    v2, v3, v4, w0, w1, w2, w3, w4, x0, x1, x2, x3, x4, y0, y1, y2, y3, y4,
    z0, z1, z2, z3, z4,
    y10, a6, a7, a8, a9, b6, b7, b8, b9, c6, c7, c8, c9, d6, d7, d8, d9,
    e6, e7, e8, e9, f6, f7, f8, f9, g6, g7, g8, g9, h6, h7, h8, h9, i6, i7,
    i8, i9, j6, j7, j8, j9, k6, k7, k8, k9, l6, l7, l8, l9, m6, m7, m8, m9,
    n6, n7, n8, n9, o6, o7, o8, o9, p6, p7, p8, p9, q6, q7, q8, q9, a10,
    r6, r7, r8, r9, s5, s6, s7, s8, s9, t5, t6, t7, t8, t9, u5, u6, u7, u8,
    u9, v5, v6, v7, v8, v9, w5, w6, w7, w8, w9, x5, x6, x7, x8, x9, y5, y6,
    y7, y8, y9, z5, z6, z7, z8, z9, b10, c10, d10, e10, f10, g10, h10, i10,
    j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10,
    x10  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, c0, c1, c2,
    c3, c4, c5, d0, d1, d2, d3, d4, d5, e0, e1, e2, e3, e4, e5, f0, f1, f2,
    f3, f4, f5, g0, g1, g2, g3, g4, g5, h0, h1, h2, h3, h4, h5, i0, i1, i2,
    i3, i4, i5, j0, j1, j2, j3, j4, j5, k0, k1, k2, k3, k4, k5, l0, l1, l2,
    l3, l4, l5, m0, m1, m2, m3, m4, m5, n0, n1, n2, n3, n4, n5, o0, o1, o2,
    o3, o4, o5, p0, p1, p2, p3, p4, p5, q0, q1, q2, q3, q4, q5, r0, r1, r2,
    r3, r4, r5, s0, s1, s2, s3, s4, t0, t1, t2, t3, t4, u0, u1, u2, u3, u4,
    v0, v1, v2, v3, v4, w0, w1, w2, w3, w4, x0, x1, x2, x3, x4, y0, y1, y2,
    y3, y4, z0, z1, z2, z3, z4;
  output y10, a6, a7, a8, a9, b6, b7, b8, b9, c6, c7, c8, c9, d6, d7, d8, d9,
    e6, e7, e8, e9, f6, f7, f8, f9, g6, g7, g8, g9, h6, h7, h8, h9, i6, i7,
    i8, i9, j6, j7, j8, j9, k6, k7, k8, k9, l6, l7, l8, l9, m6, m7, m8, m9,
    n6, n7, n8, n9, o6, o7, o8, o9, p6, p7, p8, p9, q6, q7, q8, q9, a10,
    r6, r7, r8, r9, s5, s6, s7, s8, s9, t5, t6, t7, t8, t9, u5, u6, u7, u8,
    u9, v5, v6, v7, v8, v9, w5, w6, w7, w8, w9, x5, x6, x7, x8, x9, y5, y6,
    y7, y8, y9, z5, z6, z7, z8, z9, b10, c10, d10, e10, f10, g10, h10, i10,
    j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10,
    x10;
  wire n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n501, n502, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n634, n635, n636, n637, n638, n639, n640, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n718, n719, n720,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n736, n737, n738, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n788, n789, n790, n791, n792, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n845, n846, n847, n848, n849, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n903, n904, n905, n906, n907, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n959, n960, n961, n962, n963, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1019, n1020, n1021, n1022, n1023, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1066, n1067, n1068, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101, n1102, n1103,
    n1104, n1106, n1107, n1108, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1157, n1158, n1159,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1170, n1171,
    n1172, n1174, n1175, n1176, n1178, n1179, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1204, n1205, n1206,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1237, n1238, n1239, n1240,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1262, n1263,
    n1265, n1266, n1267, n1268, n1269, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1675, n1676, n1677, n1678, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1737, n1738,
    n1739, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1817, n1818, n1819, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1873, n1874, n1875, n1877, n1878, n1879, n1880, n1881,
    n1883, n1884, n1885, n1886, n1887, n1889, n1890, n1891, n1892, n1893,
    n1895, n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1909, n1910, n1911, n1912, n1913, n1915, n1916, n1917,
    n1918, n1919, n1921, n1922, n1923, n1924, n1926, n1927, n1928, n1929,
    n1930, n1931, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1950, n1951, n1952,
    n1953, n1955, n1956, n1957, n1959, n1960, n1961, n1962, n1963, n1964,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042;
  assign n311 = ~l5 & ~m5;
  assign n312 = n5 & n311;
  assign n313 = ~z & n312;
  assign n314 = ~b0 & ~n313;
  assign n315 = l5 & m5;
  assign n316 = n5 & n315;
  assign n317 = ~z & n316;
  assign n318 = ~c0 & ~n317;
  assign n319 = ~p5 & n318;
  assign n320 = ~n314 & n319;
  assign n321 = ~p5 & ~q5;
  assign n322 = ~n314 & n321;
  assign n323 = ~q5 & ~n318;
  assign n324 = n314 & n323;
  assign n325 = ~r5 & n318;
  assign n326 = n314 & n325;
  assign n327 = ~q5 & ~r5;
  assign n328 = n314 & n327;
  assign n329 = ~n318 & n321;
  assign n330 = ~p5 & ~r5;
  assign n331 = n318 & n330;
  assign n332 = ~r5 & n321;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n329 & n333;
  assign n335 = ~n328 & n334;
  assign n336 = ~n326 & n335;
  assign n337 = ~n324 & n336;
  assign n338 = ~n322 & n337;
  assign n339 = ~n320 & n338;
  assign n340 = ~n321 & ~n330;
  assign n341 = ~n327 & n340;
  assign n342 = q5 & ~n341;
  assign n343 = ~z & n342;
  assign n344 = r5 & ~n341;
  assign n345 = ~z & n344;
  assign n346 = p5 & ~n341;
  assign n347 = ~z & n346;
  assign n348 = ~n345 & ~n347;
  assign n349 = ~n343 & n348;
  assign y10 = n339 & ~n349;
  assign n351 = k0 & q3;
  assign n352 = l0 & m3;
  assign n353 = f3 & m0;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n351 & n354;
  assign n356 = n0 & p5;
  assign n357 = o0 & r5;
  assign n358 = m5 & p0;
  assign n359 = m4 & q0;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~n356 & n361;
  assign n363 = h4 & r0;
  assign n364 = d4 & s0;
  assign n365 = t0 & w4;
  assign n366 = r4 & u0;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~n364 & n367;
  assign n369 = ~n363 & n368;
  assign n370 = n362 & n369;
  assign a6 = ~n355 | ~n370;
  assign n372 = ~x0 & ~y0;
  assign n373 = ~z0 & n372;
  assign n374 = ~a1 & n373;
  assign n375 = ~b1 & n374;
  assign n376 = ~c1 & n375;
  assign n377 = ~v0 & w0;
  assign n378 = ~p1 & ~n376;
  assign n379 = ~q1 & n378;
  assign n380 = ~p1 & ~r1;
  assign n381 = ~q1 & n380;
  assign n382 = ~n372 & ~n376;
  assign n383 = ~q1 & n382;
  assign n384 = ~r1 & ~n372;
  assign n385 = ~q1 & n384;
  assign n386 = ~n373 & ~n376;
  assign n387 = ~p1 & n386;
  assign n388 = ~r1 & ~n373;
  assign n389 = ~p1 & n388;
  assign n390 = ~n373 & n382;
  assign n391 = ~n373 & n384;
  assign n392 = n377 & ~n391;
  assign n393 = ~n390 & n392;
  assign n394 = ~n389 & n393;
  assign n395 = ~n387 & n394;
  assign n396 = ~n385 & n395;
  assign n397 = ~n383 & n396;
  assign n398 = ~n381 & n397;
  assign n399 = ~n379 & n398;
  assign n400 = ~l1 & ~m1;
  assign n401 = ~n1 & n400;
  assign v6 = b | n401;
  assign n403 = n399 & v6;
  assign n404 = ~h & ~n403;
  assign n405 = ~h1 & ~i1;
  assign n406 = ~j1 & ~o1;
  assign n407 = ~k1 & o1;
  assign n408 = ~n406 & ~n407;
  assign n409 = j1 & ~n408;
  assign n410 = e1 & ~f1;
  assign n411 = n409 & ~n410;
  assign n412 = ~n409 & n410;
  assign n413 = ~n411 & ~n412;
  assign n414 = n410 & ~n413;
  assign n415 = n405 & n414;
  assign n6 = i1 | n415;
  assign n417 = ~g1 & ~n6;
  assign n418 = ~i & n417;
  assign n419 = ~s1 & ~n418;
  assign n420 = s1 & n418;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n404 & n421;
  assign n423 = ~t1 & n422;
  assign n424 = t1 & ~n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = l1 & ~m1;
  assign n427 = ~n1 & n426;
  assign n428 = ~b & n427;
  assign n429 = ~w0 & n376;
  assign n430 = ~d1 & n429;
  assign n431 = v0 & n430;
  assign n432 = ~v6 & ~n428;
  assign n433 = ~n428 & ~n431;
  assign n434 = ~n432 & ~n433;
  assign n435 = n425 & ~n434;
  assign n436 = ~x2 & n425;
  assign n437 = ~x2 & n434;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n435 & n438;
  assign a7 = ~b & n439;
  assign n441 = v6 & ~n417;
  assign n442 = ~g & ~n441;
  assign n443 = ~l1 & m1;
  assign n444 = ~n1 & n443;
  assign n445 = ~b & n444;
  assign n446 = ~b & ~n445;
  assign n447 = ~n442 & ~n446;
  assign n448 = n405 & ~n413;
  assign n449 = n409 & n448;
  assign n450 = ~h1 & ~n449;
  assign n451 = ~v0 & n430;
  assign n452 = n417 & n450;
  assign n453 = n451 & ~n452;
  assign n454 = ~b & ~n1;
  assign n455 = l1 & m1;
  assign n456 = n454 & n455;
  assign n457 = r1 & ~v0;
  assign n458 = ~v6 & n457;
  assign n459 = ~n453 & n457;
  assign n460 = ~v6 & ~n456;
  assign n461 = ~n453 & ~n456;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~n459 & n462;
  assign n464 = ~n458 & n463;
  assign n465 = ~f & ~n464;
  assign n466 = p1 & n456;
  assign n467 = ~j & n466;
  assign n468 = q1 & n456;
  assign n469 = ~j & n468;
  assign n470 = q2 & r2;
  assign n471 = ~n469 & ~n470;
  assign n472 = ~s2 & ~n467;
  assign n473 = ~n467 & n471;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~q2 & ~r2;
  assign n476 = ~n469 & ~n475;
  assign n477 = ~n467 & n476;
  assign n478 = s2 & ~n467;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n442 & n474;
  assign n481 = n442 & n479;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n465 & ~n482;
  assign n484 = ~t2 & n483;
  assign n485 = t2 & ~n483;
  assign n486 = ~n484 & ~n485;
  assign n487 = n446 & ~n486;
  assign a8 = n447 | n487;
  assign n489 = ~d5 & ~e5;
  assign n490 = ~g5 & ~o5;
  assign n491 = ~i5 & o5;
  assign n492 = ~n490 & ~n491;
  assign n493 = g5 & ~n492;
  assign n494 = a5 & ~b5;
  assign n495 = n493 & ~n494;
  assign n496 = ~n493 & n494;
  assign n497 = ~n495 & ~n496;
  assign n498 = n494 & ~n497;
  assign n499 = n489 & n498;
  assign j10 = e5 | n499;
  assign n501 = ~c5 & ~j10;
  assign n502 = ~n5 & n311;
  assign v10 = z | n502;
  assign n504 = ~n501 & v10;
  assign n505 = ~e0 & ~n504;
  assign n506 = ~l5 & m5;
  assign n507 = ~n5 & n506;
  assign n508 = ~z & n507;
  assign n509 = ~z & ~n508;
  assign n510 = ~n505 & ~n509;
  assign n511 = n489 & ~n497;
  assign n512 = n493 & n511;
  assign n513 = ~d5 & ~n512;
  assign n514 = ~t4 & ~u4;
  assign n515 = ~v4 & n514;
  assign n516 = ~w4 & n515;
  assign n517 = ~x4 & n516;
  assign n518 = ~y4 & n517;
  assign n519 = ~s4 & n518;
  assign n520 = ~z4 & n519;
  assign n521 = ~r4 & n520;
  assign n522 = n501 & n513;
  assign n523 = n521 & ~n522;
  assign n524 = ~j5 & k5;
  assign n525 = ~r4 & r5;
  assign n526 = ~v10 & n525;
  assign n527 = ~n523 & n525;
  assign n528 = ~v10 & ~n524;
  assign n529 = ~n523 & ~n524;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n527 & n530;
  assign n532 = ~n526 & n531;
  assign n533 = ~d0 & ~n532;
  assign n534 = ~z & ~n5;
  assign n535 = n315 & n534;
  assign n536 = p5 & n535;
  assign n537 = ~h0 & n536;
  assign n538 = q5 & n535;
  assign n539 = ~h0 & n538;
  assign n540 = f3 & g3;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~h3 & ~n537;
  assign n543 = ~n537 & n541;
  assign n544 = ~n542 & ~n543;
  assign n545 = i3 & n544;
  assign n546 = ~h0 & ~n545;
  assign n547 = k3 & ~n546;
  assign n548 = p3 & n547;
  assign n549 = ~h0 & ~n548;
  assign n550 = q3 & ~n549;
  assign n551 = r3 & s3;
  assign n552 = n550 & n551;
  assign n553 = ~f3 & ~g3;
  assign n554 = ~n539 & ~n553;
  assign n555 = ~n537 & n554;
  assign n556 = h3 & ~n537;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~i3 & n557;
  assign n559 = ~h0 & ~n558;
  assign n560 = j3 & ~n559;
  assign n561 = ~p3 & n560;
  assign n562 = ~h0 & ~n561;
  assign n563 = ~q3 & ~n562;
  assign n564 = ~r3 & n563;
  assign n565 = ~s3 & n564;
  assign n566 = ~n505 & ~n552;
  assign n567 = ~n552 & ~n565;
  assign n568 = n505 & ~n565;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n566 & n569;
  assign n571 = ~n533 & n570;
  assign n572 = ~t3 & n571;
  assign n573 = t3 & ~n571;
  assign n574 = ~n572 & ~n573;
  assign n575 = n509 & ~n574;
  assign a9 = n510 | n575;
  assign n577 = ~q3 & ~r3;
  assign n578 = ~s3 & n577;
  assign n579 = ~t3 & n578;
  assign n580 = n3 & ~o3;
  assign n581 = ~p3 & n580;
  assign n582 = n579 & n581;
  assign n583 = k0 & n582;
  assign n584 = l0 & l3;
  assign n585 = p3 & q3;
  assign n586 = s3 & t3;
  assign n587 = r3 & n586;
  assign n588 = n585 & n587;
  assign n589 = m0 & n588;
  assign n590 = ~n584 & ~n589;
  assign n591 = ~n583 & n590;
  assign n592 = n0 & q5;
  assign n593 = o0 & ~n509;
  assign n594 = n5 & p0;
  assign n595 = ~j0 & ~p5;
  assign n596 = ~j0 & q5;
  assign n597 = e4 & f4;
  assign n598 = d4 & n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = i4 & ~n599;
  assign n601 = n595 & ~n600;
  assign n602 = g4 & ~n601;
  assign n603 = p4 & n602;
  assign n604 = q0 & n603;
  assign n605 = ~n594 & ~n604;
  assign n606 = ~n593 & n605;
  assign n607 = ~n592 & n606;
  assign n608 = g4 & r0;
  assign n609 = s0 & n533;
  assign n610 = t0 & v4;
  assign n611 = l5 & u0;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n609 & n612;
  assign n614 = ~n608 & n613;
  assign n615 = n607 & n614;
  assign b6 = ~n591 | ~n615;
  assign n617 = s1 & t1;
  assign n618 = ~s1 & ~t1;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n418 & ~n617;
  assign n621 = n418 & ~n618;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n619 & n622;
  assign n624 = ~n404 & n623;
  assign n625 = ~u1 & n624;
  assign n626 = u1 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n434 & n627;
  assign n629 = ~y2 & n627;
  assign n630 = ~y2 & n434;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n628 & n631;
  assign b7 = ~b & n632;
  assign n634 = ~w2 & ~x2;
  assign n635 = ~y2 & n634;
  assign n636 = ~z2 & n635;
  assign n637 = n446 & n636;
  assign n638 = n442 & ~n446;
  assign n639 = n442 & n636;
  assign n640 = ~n638 & ~n639;
  assign b8 = n637 | ~n640;
  assign n642 = l5 & ~m5;
  assign n643 = ~n5 & n642;
  assign n644 = ~z & n643;
  assign n645 = r4 & n520;
  assign n646 = ~v10 & ~n644;
  assign n647 = ~n644 & ~n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~r4 & s4;
  assign n650 = ~n514 & ~n518;
  assign n651 = ~n515 & n650;
  assign n652 = ~r5 & ~n514;
  assign n653 = ~n515 & n652;
  assign n654 = ~p5 & ~n518;
  assign n655 = ~n515 & n654;
  assign n656 = n330 & ~n515;
  assign n657 = ~q5 & ~n518;
  assign n658 = ~n514 & n657;
  assign n659 = n327 & ~n514;
  assign n660 = n321 & ~n518;
  assign n661 = ~n332 & n649;
  assign n662 = ~n660 & n661;
  assign n663 = ~n659 & n662;
  assign n664 = ~n658 & n663;
  assign n665 = ~n656 & n664;
  assign n666 = ~n655 & n665;
  assign n667 = ~n653 & n666;
  assign n668 = ~n651 & n667;
  assign n669 = v10 & n668;
  assign n670 = ~f0 & ~n669;
  assign n671 = ~u3 & ~n670;
  assign n672 = u3 & n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~l3 & n648;
  assign n675 = ~l3 & n673;
  assign n676 = ~n648 & n673;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n674 & n677;
  assign b9 = ~z & n678;
  assign n680 = ~m1 & n1;
  assign n681 = l1 & n680;
  assign n682 = ~b & n681;
  assign n683 = r1 & n456;
  assign n684 = v0 & n683;
  assign n685 = v6 & n452;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~b & n686;
  assign n688 = ~n682 & n687;
  assign n689 = ~r1 & n417;
  assign n690 = n417 & ~n456;
  assign n691 = ~n689 & ~n690;
  assign n692 = n450 & ~n691;
  assign n693 = ~v0 & n692;
  assign n694 = v0 & ~n692;
  assign n695 = ~n693 & ~n694;
  assign c6 = n688 & n695;
  assign n697 = t1 & u1;
  assign n698 = s1 & n697;
  assign n699 = ~k & ~n698;
  assign n700 = ~t1 & ~u1;
  assign n701 = ~s1 & n700;
  assign n702 = ~k & ~n701;
  assign n703 = n699 & n702;
  assign n704 = ~n418 & n699;
  assign n705 = n418 & n702;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n703 & n706;
  assign n708 = ~n404 & n707;
  assign n709 = ~v1 & n708;
  assign n710 = v1 & ~n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n434 & n711;
  assign n713 = ~z2 & n711;
  assign n714 = ~z2 & n434;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~n712 & n715;
  assign c7 = b | n716;
  assign n718 = w2 & x2;
  assign n719 = y2 & n718;
  assign n720 = z2 & n719;
  assign c8 = n446 & n720;
  assign n722 = ~g0 & n501;
  assign n723 = ~u3 & ~n722;
  assign n724 = u3 & n722;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n670 & n725;
  assign n727 = ~v3 & n726;
  assign n728 = v3 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~m3 & n648;
  assign n731 = ~m3 & n729;
  assign n732 = ~n648 & n729;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n730 & n733;
  assign c9 = ~z & n734;
  assign n736 = ~w0 & ~n694;
  assign n737 = w0 & n694;
  assign n738 = ~n736 & ~n737;
  assign d6 = n688 & n738;
  assign n740 = v1 & ~n699;
  assign n741 = ~v1 & ~n702;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n418 & ~n740;
  assign n744 = n418 & ~n741;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n742 & n745;
  assign n747 = ~n404 & n746;
  assign n748 = ~w1 & n747;
  assign n749 = w1 & ~n747;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~n434 & n750;
  assign n752 = ~a3 & n750;
  assign n753 = ~a3 & n434;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n751 & n754;
  assign d7 = b | n755;
  assign n757 = t2 & n474;
  assign n758 = ~j & ~n757;
  assign n759 = ~t2 & n479;
  assign n760 = ~j & ~n759;
  assign n761 = n758 & n760;
  assign n762 = ~n442 & n758;
  assign n763 = n442 & n760;
  assign n764 = ~n762 & ~n763;
  assign n765 = ~n761 & n764;
  assign n766 = ~n465 & n765;
  assign n767 = ~w2 & ~n766;
  assign n768 = w2 & n766;
  assign n769 = ~n767 & ~n768;
  assign d8 = n446 & n769;
  assign n771 = u3 & v3;
  assign n772 = ~u3 & ~v3;
  assign n773 = ~n722 & ~n771;
  assign n774 = ~n771 & ~n772;
  assign n775 = n722 & ~n772;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n773 & n776;
  assign n778 = ~n670 & n777;
  assign n779 = ~w3 & n778;
  assign n780 = w3 & ~n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~n3 & n648;
  assign n783 = ~n3 & n781;
  assign n784 = ~n648 & n781;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n782 & n785;
  assign d9 = ~z & n786;
  assign n788 = v0 & w0;
  assign n789 = ~n692 & n788;
  assign n790 = ~x0 & ~n789;
  assign n791 = x0 & n789;
  assign n792 = ~n790 & ~n791;
  assign e6 = n688 & n792;
  assign n794 = v1 & w1;
  assign n795 = ~n699 & n794;
  assign n796 = ~w1 & n741;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n418 & ~n795;
  assign n799 = n418 & ~n796;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~n797 & n800;
  assign n802 = ~n404 & n801;
  assign n803 = ~x1 & n802;
  assign n804 = x1 & ~n802;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n434 & n805;
  assign n807 = ~b3 & n805;
  assign n808 = ~b3 & n434;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n806 & n809;
  assign e7 = b | n810;
  assign n812 = w2 & ~n758;
  assign n813 = ~w2 & ~n760;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n442 & ~n812;
  assign n816 = n442 & ~n813;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~n814 & n817;
  assign n819 = ~n465 & n818;
  assign n820 = ~x2 & ~n819;
  assign n821 = x2 & n819;
  assign n822 = ~n820 & ~n821;
  assign e8 = n446 & n822;
  assign n824 = v3 & w3;
  assign n825 = u3 & n824;
  assign n826 = ~i0 & ~n825;
  assign n827 = ~v3 & ~w3;
  assign n828 = ~u3 & n827;
  assign n829 = ~i0 & ~n828;
  assign n830 = ~n722 & n826;
  assign n831 = n826 & n829;
  assign n832 = n722 & n829;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n830 & n833;
  assign n835 = ~n670 & n834;
  assign n836 = ~x3 & n835;
  assign n837 = x3 & ~n835;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~o3 & n648;
  assign n840 = ~o3 & n838;
  assign n841 = ~n648 & n838;
  assign n842 = ~n840 & ~n841;
  assign n843 = ~n839 & n842;
  assign e9 = z | n843;
  assign n845 = x0 & n788;
  assign n846 = ~n692 & n845;
  assign n847 = ~y0 & ~n846;
  assign n848 = y0 & n846;
  assign n849 = ~n847 & ~n848;
  assign f6 = n688 & n849;
  assign n851 = w1 & x1;
  assign n852 = v1 & n851;
  assign n853 = ~n699 & n852;
  assign n854 = ~k & ~n853;
  assign n855 = ~w1 & ~x1;
  assign n856 = ~v1 & n855;
  assign n857 = ~n702 & n856;
  assign n858 = ~k & ~n857;
  assign n859 = n854 & n858;
  assign n860 = ~n418 & n854;
  assign n861 = n418 & n858;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n859 & n862;
  assign n864 = ~n404 & n863;
  assign n865 = ~y1 & n864;
  assign n866 = y1 & ~n864;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n434 & n867;
  assign n869 = ~c3 & n867;
  assign n870 = ~c3 & n434;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n868 & n871;
  assign f7 = ~b & n872;
  assign n874 = n718 & ~n758;
  assign n875 = ~x2 & n813;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n442 & ~n874;
  assign n878 = n442 & ~n875;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~n876 & n879;
  assign n881 = ~n465 & n880;
  assign n882 = ~y2 & ~n881;
  assign n883 = y2 & n881;
  assign n884 = ~n882 & ~n883;
  assign f8 = n446 & n884;
  assign n886 = x3 & ~n826;
  assign n887 = ~x3 & ~n829;
  assign n888 = ~n722 & ~n886;
  assign n889 = ~n886 & ~n887;
  assign n890 = n722 & ~n887;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n888 & n891;
  assign n893 = ~n670 & n892;
  assign n894 = ~y3 & n893;
  assign n895 = y3 & ~n893;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~p3 & n648;
  assign n898 = ~p3 & n896;
  assign n899 = ~n648 & n896;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n897 & n900;
  assign f9 = z | n901;
  assign n903 = y0 & n845;
  assign n904 = ~n692 & n903;
  assign n905 = ~z0 & ~n904;
  assign n906 = z0 & n904;
  assign n907 = ~n905 & ~n906;
  assign g6 = n688 & n907;
  assign n909 = y1 & ~n854;
  assign n910 = ~y1 & ~n858;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n418 & ~n909;
  assign n913 = n418 & ~n910;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~n911 & n914;
  assign n916 = ~n404 & n915;
  assign n917 = ~z1 & n916;
  assign n918 = z1 & ~n916;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n434 & n919;
  assign n921 = ~d3 & n919;
  assign n922 = ~d3 & n434;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n920 & n923;
  assign g7 = b | n924;
  assign n926 = x2 & y2;
  assign n927 = w2 & n926;
  assign n928 = ~n758 & n927;
  assign n929 = ~y2 & n875;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n442 & ~n928;
  assign n932 = n442 & ~n929;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n930 & n933;
  assign n935 = ~n465 & n934;
  assign n936 = ~z2 & n935;
  assign n937 = z2 & ~n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = n446 & ~n938;
  assign g8 = n447 | n939;
  assign n941 = x3 & y3;
  assign n942 = ~n826 & n941;
  assign n943 = ~y3 & n887;
  assign n944 = ~n722 & ~n942;
  assign n945 = ~n942 & ~n943;
  assign n946 = n722 & ~n943;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~n944 & n947;
  assign n949 = ~n670 & n948;
  assign n950 = ~z3 & n949;
  assign n951 = z3 & ~n949;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~q3 & n648;
  assign n954 = ~q3 & n952;
  assign n955 = ~n648 & n952;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n953 & n956;
  assign g9 = z | n957;
  assign n959 = z0 & n903;
  assign n960 = ~n692 & n959;
  assign n961 = ~a1 & ~n960;
  assign n962 = a1 & n960;
  assign n963 = ~n961 & ~n962;
  assign h6 = n688 & n963;
  assign n965 = y1 & z1;
  assign n966 = ~n854 & n965;
  assign n967 = ~z1 & n910;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~n418 & ~n966;
  assign n970 = n418 & ~n967;
  assign n971 = ~n969 & ~n970;
  assign n972 = ~n968 & n971;
  assign n973 = ~n404 & n972;
  assign n974 = ~a2 & n973;
  assign n975 = a2 & ~n973;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n434 & n976;
  assign n978 = ~e3 & n976;
  assign n979 = ~e3 & n434;
  assign n980 = ~n978 & ~n979;
  assign n981 = ~n977 & n980;
  assign h7 = b | n981;
  assign n983 = v2 & ~n758;
  assign n984 = u2 & ~n760;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n442 & ~n983;
  assign n987 = n442 & ~n984;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n985 & n988;
  assign n990 = ~n465 & n989;
  assign n991 = ~a3 & n990;
  assign n992 = a3 & ~n990;
  assign n993 = ~n991 & ~n992;
  assign n994 = n446 & ~n993;
  assign h8 = n447 | n994;
  assign n996 = y3 & z3;
  assign n997 = x3 & n996;
  assign n998 = ~n826 & n997;
  assign n999 = ~i0 & ~n998;
  assign n1000 = ~y3 & ~z3;
  assign n1001 = ~x3 & n1000;
  assign n1002 = ~n829 & n1001;
  assign n1003 = ~i0 & ~n1002;
  assign n1004 = ~n722 & n999;
  assign n1005 = n999 & n1003;
  assign n1006 = n722 & n1003;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1004 & n1007;
  assign n1009 = ~n670 & n1008;
  assign n1010 = ~a4 & n1009;
  assign n1011 = a4 & ~n1009;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~r3 & n648;
  assign n1014 = ~r3 & n1012;
  assign n1015 = ~n648 & n1012;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n1013 & n1016;
  assign h9 = ~z & n1017;
  assign n1019 = a1 & n959;
  assign n1020 = ~n692 & n1019;
  assign n1021 = ~b1 & ~n1020;
  assign n1022 = b1 & n1020;
  assign n1023 = ~n1021 & ~n1022;
  assign i6 = n688 & n1023;
  assign i7 = b | ~b2;
  assign n1026 = a3 & n983;
  assign n1027 = ~j & ~n1026;
  assign n1028 = ~a3 & n984;
  assign n1029 = ~j & ~n1028;
  assign n1030 = n1027 & n1029;
  assign n1031 = ~n442 & n1027;
  assign n1032 = n442 & n1029;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = ~n1030 & n1033;
  assign n1035 = ~n465 & n1034;
  assign n1036 = ~b3 & n1035;
  assign n1037 = b3 & ~n1035;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = n446 & ~n1038;
  assign i8 = n447 | n1039;
  assign n1041 = a4 & ~n999;
  assign n1042 = ~a4 & ~n1003;
  assign n1043 = ~n722 & ~n1041;
  assign n1044 = ~n1041 & ~n1042;
  assign n1045 = n722 & ~n1042;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = ~n1043 & n1046;
  assign n1048 = ~n670 & n1047;
  assign n1049 = ~b4 & n1048;
  assign n1050 = b4 & ~n1048;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = ~s3 & n648;
  assign n1053 = ~s3 & n1051;
  assign n1054 = ~n648 & n1051;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1052 & n1055;
  assign i9 = z | n1056;
  assign n1058 = a1 & z0;
  assign n1059 = b1 & n1058;
  assign n1060 = n903 & n1059;
  assign n1061 = ~n692 & n1060;
  assign n1062 = ~c1 & ~n1061;
  assign n1063 = c1 & n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign j6 = n688 & n1064;
  assign n1066 = ~b2 & ~c2;
  assign n1067 = b2 & c2;
  assign n1068 = ~n1066 & ~n1067;
  assign j7 = b | n1068;
  assign n1070 = b3 & ~n1027;
  assign n1071 = ~b3 & ~n1029;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = n442 & ~n1071;
  assign n1074 = ~n442 & ~n1070;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = ~n1072 & n1075;
  assign n1077 = ~n465 & n1076;
  assign n1078 = ~c3 & ~n1077;
  assign n1079 = c3 & n1077;
  assign n1080 = ~n1078 & ~n1079;
  assign j8 = n446 & n1080;
  assign n1082 = a4 & b4;
  assign n1083 = ~n999 & n1082;
  assign n1084 = ~b4 & n1042;
  assign n1085 = ~n722 & ~n1083;
  assign n1086 = ~n1083 & ~n1084;
  assign n1087 = n722 & ~n1084;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n1085 & n1088;
  assign n1090 = ~n670 & n1089;
  assign n1091 = ~c4 & n1090;
  assign n1092 = c4 & ~n1090;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = ~t3 & n648;
  assign n1095 = ~t3 & n1093;
  assign n1096 = ~n648 & n1093;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n1094 & n1097;
  assign j9 = z | n1098;
  assign n1100 = c1 & ~n692;
  assign n1101 = n1060 & n1100;
  assign n1102 = d1 & n1101;
  assign n1103 = ~d1 & ~n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign k6 = n688 & n1104;
  assign n1106 = ~d2 & ~n1067;
  assign n1107 = d2 & n1067;
  assign n1108 = ~n1106 & ~n1107;
  assign k7 = b | n1108;
  assign n1110 = c3 & n1070;
  assign n1111 = ~c3 & n1071;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n442 & ~n1110;
  assign n1114 = n442 & ~n1111;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~n1112 & n1115;
  assign n1117 = ~n465 & n1116;
  assign n1118 = ~d3 & n1117;
  assign n1119 = d3 & ~n1117;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = n446 & ~n1120;
  assign k8 = n447 | n1121;
  assign k9 = z | ~d4;
  assign n1124 = ~l & ~p1;
  assign n1125 = ~l & q1;
  assign n1126 = c2 & d2;
  assign n1127 = b2 & n1126;
  assign n1128 = ~n1125 & ~n1127;
  assign n1129 = g2 & ~n1128;
  assign n1130 = n1124 & ~n1129;
  assign n1131 = ~e2 & ~n1130;
  assign n1132 = e2 & n1130;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = e2 & ~n1130;
  assign n1135 = n2 & n1134;
  assign n1136 = ~n682 & ~n1135;
  assign n1137 = n1133 & n1136;
  assign n1138 = ~s1 & n1133;
  assign n1139 = ~s1 & ~n1136;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1137 & n1140;
  assign l7 = b | n1141;
  assign n1143 = c3 & d3;
  assign n1144 = n1070 & n1143;
  assign n1145 = ~d3 & n1111;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n442 & ~n1144;
  assign n1148 = n442 & ~n1145;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = ~n1146 & n1149;
  assign n1151 = ~n465 & n1150;
  assign n1152 = ~e3 & n1151;
  assign n1153 = e3 & ~n1151;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = n446 & ~n1154;
  assign l8 = n447 | n1155;
  assign n1157 = ~d4 & ~e4;
  assign n1158 = d4 & e4;
  assign n1159 = ~n1157 & ~n1158;
  assign l9 = z | n1159;
  assign n1161 = ~f2 & n1134;
  assign n1162 = f2 & ~n1134;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = n1136 & n1163;
  assign n1165 = ~t1 & n1163;
  assign n1166 = ~t1 & ~n1136;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1164 & n1167;
  assign m7 = b | n1168;
  assign n1170 = ~f3 & n533;
  assign n1171 = f3 & ~n533;
  assign n1172 = ~n1170 & ~n1171;
  assign m8 = n509 & n1172;
  assign n1174 = ~f4 & ~n1158;
  assign n1175 = f4 & n1158;
  assign n1176 = ~n1174 & ~n1175;
  assign m9 = z | n1176;
  assign n1178 = ~g2 & n1128;
  assign n1179 = ~n1129 & ~n1178;
  assign n7 = b | n1179;
  assign n1181 = ~f3 & ~n505;
  assign n1182 = f3 & n505;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n533 & n1183;
  assign n1185 = ~g3 & ~n1184;
  assign n1186 = g3 & n1184;
  assign n1187 = ~n1185 & ~n1186;
  assign n8 = n509 & n1187;
  assign n1189 = ~m5 & n5;
  assign n1190 = l5 & n1189;
  assign n1191 = ~z & n1190;
  assign n1192 = ~n603 & ~n1191;
  assign n1193 = ~g4 & ~n601;
  assign n1194 = g4 & n601;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1192 & n1195;
  assign n1197 = ~u3 & n1195;
  assign n1198 = ~u3 & ~n1192;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~n1196 & n1199;
  assign n9 = z | n1200;
  assign n1202 = ~b & ~n682;
  assign n1203 = ~n410 & n1202;
  assign n1204 = ~h1 & n1202;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = h1 & ~n1205;
  assign o6 = n449 | n1206;
  assign n1208 = f2 & n1134;
  assign n1209 = ~h2 & n1208;
  assign n1210 = h2 & ~n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = n1136 & n1211;
  assign n1213 = ~u1 & n1211;
  assign n1214 = ~u1 & ~n1136;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = ~n1212 & n1215;
  assign o7 = b | n1216;
  assign n1218 = ~n505 & n541;
  assign n1219 = n541 & n554;
  assign n1220 = n505 & n554;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n1218 & n1221;
  assign n1223 = ~n533 & n1222;
  assign n1224 = ~h3 & ~n1223;
  assign n1225 = h3 & n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign o8 = n509 & n1226;
  assign n1228 = ~h4 & n602;
  assign n1229 = h4 & ~n602;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = n1192 & n1230;
  assign n1232 = ~v3 & n1230;
  assign n1233 = ~v3 & ~n1192;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~n1231 & n1234;
  assign o9 = z | n1235;
  assign n1237 = ~i1 & n1202;
  assign n1238 = ~n409 & n1202;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = i1 & ~n1239;
  assign p6 = n415 | n1240;
  assign n1242 = f2 & h2;
  assign n1243 = n1134 & n1242;
  assign n1244 = ~i2 & n1243;
  assign n1245 = i2 & ~n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = n1136 & n1246;
  assign n1248 = ~v1 & n1246;
  assign n1249 = ~v1 & ~n1136;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n1247 & n1250;
  assign p7 = b | n1251;
  assign n1253 = ~n505 & n544;
  assign n1254 = n505 & n557;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n533 & ~n1255;
  assign n1257 = ~i3 & n1256;
  assign n1258 = i3 & ~n1256;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = n509 & ~n1259;
  assign p8 = n510 | n1260;
  assign n1262 = ~i4 & n599;
  assign n1263 = ~n600 & ~n1262;
  assign p9 = z | n1263;
  assign n1265 = ~n428 & ~n682;
  assign n1266 = j1 & n1135;
  assign n1267 = ~j1 & ~n1135;
  assign n1268 = ~b & ~n1267;
  assign n1269 = ~n1266 & n1268;
  assign q6 = ~n1265 | n1269;
  assign n1271 = i2 & n1243;
  assign n1272 = ~j2 & n1271;
  assign n1273 = j2 & ~n1271;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = n1136 & n1274;
  assign n1276 = ~w1 & n1274;
  assign n1277 = ~w1 & ~n1136;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~n1275 & n1278;
  assign q7 = b | n1279;
  assign n1281 = ~l3 & ~m3;
  assign n1282 = ~n3 & n1281;
  assign n1283 = ~o3 & n1282;
  assign n1284 = n505 & ~n509;
  assign n1285 = n505 & n1283;
  assign n1286 = n509 & n1283;
  assign n1287 = ~n1285 & ~n1286;
  assign q8 = n1284 | ~n1287;
  assign n1289 = h4 & n602;
  assign n1290 = ~j4 & n1289;
  assign n1291 = j4 & ~n1289;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = n1192 & n1292;
  assign n1294 = ~w3 & n1292;
  assign n1295 = ~w3 & ~n1192;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1293 & n1296;
  assign q9 = z | n1297;
  assign n1299 = r5 & n535;
  assign n1300 = r4 & n1299;
  assign n1301 = v10 & n522;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~z & n1302;
  assign n1304 = ~n1191 & n1303;
  assign n1305 = ~r5 & n501;
  assign n1306 = n501 & ~n535;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = n513 & ~n1307;
  assign n1309 = r4 & s4;
  assign n1310 = ~n1308 & n1309;
  assign n1311 = ~t4 & ~n1310;
  assign n1312 = t4 & n1310;
  assign n1313 = ~n1311 & ~n1312;
  assign a10 = n1304 & n1313;
  assign n1315 = i2 & j2;
  assign n1316 = n1243 & n1315;
  assign n1317 = ~l & ~n1316;
  assign n1318 = ~k2 & ~n1317;
  assign n1319 = k2 & n1317;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = n1136 & n1320;
  assign n1322 = ~x1 & n1320;
  assign n1323 = ~x1 & ~n1136;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1321 & n1324;
  assign r7 = b | n1325;
  assign n1327 = l3 & m3;
  assign n1328 = n3 & n1327;
  assign n1329 = o3 & n1328;
  assign r8 = n509 & n1329;
  assign n1331 = h4 & j4;
  assign n1332 = n602 & n1331;
  assign n1333 = ~k4 & n1332;
  assign n1334 = k4 & ~n1332;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = n1192 & n1335;
  assign n1337 = ~x3 & n1335;
  assign n1338 = ~x3 & ~n1192;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n1336 & n1339;
  assign r9 = z | n1340;
  assign n1342 = m & e3;
  assign n1343 = n & a3;
  assign n1344 = o & t2;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1342 & n1345;
  assign n1347 = p & a2;
  assign n1348 = q & x1;
  assign n1349 = r & u1;
  assign n1350 = s & o2;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1348 & n1351;
  assign n1353 = ~n1347 & n1352;
  assign n1354 = t & j2;
  assign n1355 = u & g2;
  assign n1356 = v & d1;
  assign n1357 = w & y0;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~n1355 & n1358;
  assign n1360 = ~n1354 & n1359;
  assign n1361 = n1353 & n1360;
  assign s5 = ~n1346 | ~n1361;
  assign n1363 = n410 & n445;
  assign n1364 = d3 & e3;
  assign n1365 = c3 & n1364;
  assign n1366 = ~b3 & ~c3;
  assign n1367 = ~d3 & n1366;
  assign n1368 = ~e3 & n1367;
  assign n1369 = y2 & ~z2;
  assign n1370 = ~a3 & n1369;
  assign n1371 = n1368 & n1370;
  assign n1372 = n410 & ~n1371;
  assign n1373 = n1365 & n1372;
  assign n1374 = n456 & ~n1373;
  assign n1375 = ~n428 & ~n1374;
  assign n1376 = ~n1363 & n1375;
  assign s6 = ~b & ~n1376;
  assign n1378 = k2 & ~n1317;
  assign n1379 = ~l2 & n1378;
  assign n1380 = l2 & ~n1378;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = n1136 & n1381;
  assign n1383 = ~y1 & n1381;
  assign n1384 = ~y1 & ~n1136;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n1382 & n1385;
  assign s7 = b | n1386;
  assign n1388 = ~n505 & n546;
  assign n1389 = n546 & n559;
  assign n1390 = n505 & n559;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1388 & n1391;
  assign n1393 = ~n533 & n1392;
  assign n1394 = ~l3 & ~n1393;
  assign n1395 = l3 & n1393;
  assign n1396 = ~n1394 & ~n1395;
  assign s8 = n509 & n1396;
  assign n1398 = k4 & n1332;
  assign n1399 = ~l4 & n1398;
  assign n1400 = l4 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = n1192 & n1401;
  assign n1403 = ~y3 & n1401;
  assign n1404 = ~y3 & ~n1192;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1402 & n1405;
  assign s9 = z | n1406;
  assign n1408 = m & d3;
  assign n1409 = n & z2;
  assign n1410 = o & s2;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~n1408 & n1411;
  assign n1413 = p & z1;
  assign n1414 = q & w1;
  assign n1415 = r & t1;
  assign n1416 = s & m2;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = ~n1414 & n1417;
  assign n1419 = ~n1413 & n1418;
  assign n1420 = t & i2;
  assign n1421 = u & d2;
  assign n1422 = v & c1;
  assign n1423 = w & x0;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1421 & n1424;
  assign n1426 = ~n1420 & n1425;
  assign n1427 = n1419 & n1426;
  assign t5 = ~n1412 | ~n1427;
  assign n1429 = n1 & n455;
  assign n1430 = ~b & n1429;
  assign n1431 = ~m1 & n1371;
  assign n1432 = ~n1430 & n1431;
  assign n1433 = ~m1 & n410;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = ~m1 & ~n456;
  assign n1436 = ~n1430 & n1435;
  assign n1437 = ~n1 & n1371;
  assign n1438 = ~n1430 & n1437;
  assign n1439 = ~n1 & n410;
  assign n1440 = ~n1430 & n1439;
  assign n1441 = ~n1 & ~n456;
  assign n1442 = ~n1430 & n1441;
  assign n1443 = ~n1440 & ~n1442;
  assign n1444 = ~n1438 & n1443;
  assign n1445 = ~n1436 & n1444;
  assign n1446 = ~n1434 & n1445;
  assign n1447 = ~n1432 & n1446;
  assign n1448 = n1 & n400;
  assign n1449 = ~b & n1448;
  assign n1450 = n456 & n1371;
  assign n1451 = ~c & r1;
  assign n1452 = ~n1102 & n1451;
  assign n1453 = ~c & ~d1;
  assign n1454 = ~r1 & n1453;
  assign n1455 = ~n1102 & n1453;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1452 & n1456;
  assign n1458 = v6 & n1457;
  assign n1459 = ~n1450 & ~n1458;
  assign n1460 = ~n445 & n1459;
  assign n1461 = ~n1449 & n1460;
  assign n1462 = ~n1447 & n1461;
  assign t6 = ~b & ~n1462;
  assign n1464 = k2 & l2;
  assign n1465 = ~n1317 & n1464;
  assign n1466 = ~m2 & n1465;
  assign n1467 = m2 & ~n1465;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = n1136 & n1468;
  assign n1470 = ~z1 & n1468;
  assign n1471 = ~z1 & ~n1136;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n1469 & n1472;
  assign t7 = b | n1473;
  assign n1475 = l3 & ~n546;
  assign n1476 = ~l3 & ~n559;
  assign n1477 = ~n505 & ~n1475;
  assign n1478 = ~n1475 & ~n1476;
  assign n1479 = n505 & ~n1476;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = ~n1477 & n1480;
  assign n1482 = ~n533 & n1481;
  assign n1483 = ~m3 & ~n1482;
  assign n1484 = m3 & n1482;
  assign n1485 = ~n1483 & ~n1484;
  assign t8 = n509 & n1485;
  assign n1487 = k4 & l4;
  assign n1488 = n1332 & n1487;
  assign n1489 = ~j0 & ~n1488;
  assign n1490 = ~m4 & ~n1489;
  assign n1491 = m4 & n1489;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n1192 & n1492;
  assign n1494 = ~z3 & n1492;
  assign n1495 = ~z3 & ~n1192;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1493 & n1496;
  assign t9 = z | n1497;
  assign n1499 = m & c3;
  assign n1500 = n & y2;
  assign n1501 = o & r2;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1499 & n1502;
  assign n1504 = p & y1;
  assign n1505 = q & v1;
  assign n1506 = r & s1;
  assign n1507 = s & l2;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1505 & n1508;
  assign n1510 = ~n1504 & n1509;
  assign n1511 = t & h2;
  assign n1512 = u & c2;
  assign n1513 = v & b1;
  assign n1514 = w & w0;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1512 & n1515;
  assign n1517 = ~n1511 & n1516;
  assign n1518 = n1510 & n1517;
  assign u5 = ~n1503 | ~n1518;
  assign n1520 = ~n1365 & ~n1430;
  assign n1521 = n1371 & ~n1430;
  assign n1522 = ~n410 & ~n1430;
  assign n1523 = ~n456 & ~n1430;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1521 & n1524;
  assign n1526 = ~n1520 & n1525;
  assign n1527 = ~n428 & ~n1371;
  assign n1528 = ~n1449 & n1527;
  assign n1529 = ~n428 & ~n456;
  assign n1530 = ~n1449 & n1529;
  assign n1531 = ~n1528 & ~n1530;
  assign n1532 = ~n1526 & ~n1531;
  assign u6 = ~b & ~n1532;
  assign n1534 = ~b & ~n1136;
  assign n1535 = j2 & k2;
  assign n1536 = i2 & n1535;
  assign n1537 = m2 & o2;
  assign n1538 = l2 & n1537;
  assign n1539 = n1536 & n1538;
  assign n1540 = n1242 & n1539;
  assign u7 = ~n1534 & n1540;
  assign n1542 = ~n546 & n1327;
  assign n1543 = ~m3 & n1476;
  assign n1544 = ~n505 & ~n1542;
  assign n1545 = ~n1542 & ~n1543;
  assign n1546 = n505 & ~n1543;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1544 & n1547;
  assign n1549 = ~n533 & n1548;
  assign n1550 = ~n3 & ~n1549;
  assign n1551 = n3 & n1549;
  assign n1552 = ~n1550 & ~n1551;
  assign u8 = n509 & n1552;
  assign n1554 = m4 & ~n1489;
  assign n1555 = ~n4 & n1554;
  assign n1556 = n4 & ~n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = n1192 & n1557;
  assign n1559 = ~a4 & n1557;
  assign n1560 = ~a4 & ~n1192;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1558 & n1561;
  assign u9 = z | n1562;
  assign n1564 = m & b3;
  assign n1565 = n & x2;
  assign n1566 = o & q2;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1564 & n1567;
  assign n1569 = p & p1;
  assign n1570 = q & r1;
  assign n1571 = r & m1;
  assign n1572 = s & k2;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1570 & n1573;
  assign n1575 = ~n1569 & n1574;
  assign n1576 = t & f2;
  assign n1577 = u & b2;
  assign n1578 = v & a1;
  assign n1579 = w & v0;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1577 & n1580;
  assign n1582 = ~n1576 & n1581;
  assign n1583 = n1575 & n1582;
  assign v5 = ~n1568 | ~n1583;
  assign n1585 = m2 & n1465;
  assign n1586 = ~o2 & n1585;
  assign n1587 = o2 & ~n1585;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = n1136 & n1588;
  assign n1590 = ~a2 & n1588;
  assign n1591 = ~a2 & ~n1136;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n1589 & n1592;
  assign v7 = b | n1593;
  assign n1595 = m3 & n3;
  assign n1596 = l3 & n1595;
  assign n1597 = ~n546 & n1596;
  assign n1598 = ~n3 & n1543;
  assign n1599 = ~n505 & ~n1597;
  assign n1600 = ~n1597 & ~n1598;
  assign n1601 = n505 & ~n1598;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1599 & n1602;
  assign n1604 = ~n533 & n1603;
  assign n1605 = ~o3 & n1604;
  assign n1606 = o3 & ~n1604;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n509 & ~n1607;
  assign v8 = n510 | n1608;
  assign n1610 = m4 & n4;
  assign n1611 = ~n1489 & n1610;
  assign n1612 = ~o4 & n1611;
  assign n1613 = o4 & ~n1611;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = n1192 & n1614;
  assign n1616 = ~b4 & n1614;
  assign n1617 = ~b4 & ~n1192;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = ~n1615 & n1618;
  assign v9 = z | n1619;
  assign n1621 = m & n1371;
  assign n1622 = n & w2;
  assign n1623 = o & n1365;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n1621 & n1624;
  assign n1626 = p & q1;
  assign n1627 = q & ~n446;
  assign n1628 = r & n1;
  assign n1629 = s & n1135;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = ~n1627 & n1630;
  assign n1632 = ~n1626 & n1631;
  assign n1633 = t & e2;
  assign n1634 = u & n465;
  assign n1635 = v & z0;
  assign n1636 = w & l1;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = ~n1634 & n1637;
  assign n1639 = ~n1633 & n1638;
  assign n1640 = n1632 & n1639;
  assign w5 = ~n1625 | ~n1640;
  assign n1642 = ~d & ~n1449;
  assign n1643 = ~e & ~n1430;
  assign n1644 = ~q1 & n1643;
  assign n1645 = ~n1642 & n1644;
  assign n1646 = ~q1 & ~r1;
  assign n1647 = ~n1642 & n1646;
  assign n1648 = ~r1 & ~n1643;
  assign n1649 = n1642 & n1648;
  assign n1650 = ~p1 & n1643;
  assign n1651 = n1642 & n1650;
  assign n1652 = n380 & n1642;
  assign n1653 = ~n1643 & n1646;
  assign n1654 = ~p1 & ~q1;
  assign n1655 = n1643 & n1654;
  assign n1656 = ~r1 & n1654;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = ~n1653 & n1657;
  assign n1659 = ~n1652 & n1658;
  assign n1660 = ~n1651 & n1659;
  assign n1661 = ~n1649 & n1660;
  assign n1662 = ~n1647 & n1661;
  assign n1663 = ~n1645 & n1662;
  assign n1664 = ~n380 & ~n1654;
  assign n1665 = ~n1646 & n1664;
  assign n1666 = q1 & ~n1665;
  assign n1667 = ~b & n1666;
  assign n1668 = r1 & ~n1665;
  assign n1669 = ~b & n1668;
  assign n1670 = p1 & ~n1665;
  assign n1671 = ~b & n1670;
  assign n1672 = ~n1669 & ~n1671;
  assign n1673 = ~n1667 & n1672;
  assign w6 = n1663 | n1673;
  assign n1675 = ~a & n1266;
  assign n1676 = ~a & p2;
  assign n1677 = p2 & ~n1266;
  assign n1678 = ~n1676 & ~n1677;
  assign w7 = n1675 | ~n1678;
  assign n1680 = ~n505 & ~n547;
  assign n1681 = ~n547 & ~n560;
  assign n1682 = n505 & ~n560;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1680 & n1683;
  assign n1685 = ~n533 & n1684;
  assign n1686 = ~p3 & n1685;
  assign n1687 = p3 & ~n1685;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = n509 & ~n1688;
  assign w8 = n510 | n1689;
  assign n1691 = ~z & ~n1192;
  assign n1692 = l4 & m4;
  assign n1693 = k4 & n1692;
  assign n1694 = o4 & q4;
  assign n1695 = n4 & n1694;
  assign n1696 = n1693 & n1695;
  assign n1697 = n1331 & n1696;
  assign w9 = ~n1691 & n1697;
  assign n1699 = k0 & t3;
  assign n1700 = l0 & p3;
  assign n1701 = i3 & m0;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1699 & n1702;
  assign n1704 = c4 & n0;
  assign n1705 = o0 & z3;
  assign n1706 = p0 & w3;
  assign n1707 = q0 & q4;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n1705 & n1708;
  assign n1710 = ~n1704 & n1709;
  assign n1711 = l4 & r0;
  assign n1712 = i4 & s0;
  assign n1713 = t0 & z4;
  assign n1714 = u0 & u4;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1712 & n1715;
  assign n1717 = ~n1711 & n1716;
  assign n1718 = n1710 & n1717;
  assign x5 = ~n1703 | ~n1718;
  assign n1720 = ~r1 & n1643;
  assign n1721 = ~n1642 & n1720;
  assign n1722 = n380 & ~n1642;
  assign n1723 = ~p1 & ~n1643;
  assign n1724 = n1642 & n1723;
  assign n1725 = n1642 & n1644;
  assign n1726 = n1642 & n1654;
  assign n1727 = n380 & ~n1643;
  assign n1728 = n1643 & n1646;
  assign n1729 = ~n1656 & ~n1728;
  assign n1730 = ~n1727 & n1729;
  assign n1731 = ~n1726 & n1730;
  assign n1732 = ~n1725 & n1731;
  assign n1733 = ~n1724 & n1732;
  assign n1734 = ~n1722 & n1733;
  assign n1735 = ~n1721 & n1734;
  assign x6 = ~n1673 & n1735;
  assign n1737 = ~q2 & n465;
  assign n1738 = q2 & ~n465;
  assign n1739 = ~n1737 & ~n1738;
  assign x7 = n446 & n1739;
  assign n1741 = ~n505 & n549;
  assign n1742 = n549 & n562;
  assign n1743 = n505 & n562;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = ~n1741 & n1744;
  assign n1746 = ~n533 & n1745;
  assign n1747 = ~q3 & n1746;
  assign n1748 = q3 & ~n1746;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n509 & ~n1749;
  assign x8 = n510 | n1750;
  assign n1752 = o4 & n1611;
  assign n1753 = ~q4 & n1752;
  assign n1754 = q4 & ~n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = n1192 & n1755;
  assign n1757 = ~c4 & n1755;
  assign n1758 = ~c4 & ~n1192;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1756 & n1759;
  assign x9 = z | n1760;
  assign n1762 = k0 & s3;
  assign n1763 = l0 & o3;
  assign n1764 = h3 & m0;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n1762 & n1765;
  assign n1767 = b4 & n0;
  assign n1768 = o0 & y3;
  assign n1769 = p0 & v3;
  assign n1770 = o4 & q0;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = ~n1768 & n1771;
  assign n1773 = ~n1767 & n1772;
  assign n1774 = k4 & r0;
  assign n1775 = f4 & s0;
  assign n1776 = t0 & y4;
  assign n1777 = t4 & u0;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1775 & n1778;
  assign n1780 = ~n1774 & n1779;
  assign n1781 = n1773 & n1780;
  assign y5 = ~n1766 | ~n1781;
  assign n1783 = ~n1642 & n1650;
  assign n1784 = ~n1642 & n1654;
  assign n1785 = ~q1 & ~n1643;
  assign n1786 = n1642 & n1785;
  assign n1787 = n1642 & n1720;
  assign n1788 = n1642 & n1646;
  assign n1789 = ~n1643 & n1654;
  assign n1790 = n380 & n1643;
  assign n1791 = ~n1656 & ~n1790;
  assign n1792 = ~n1789 & n1791;
  assign n1793 = ~n1788 & n1792;
  assign n1794 = ~n1787 & n1793;
  assign n1795 = ~n1786 & n1794;
  assign n1796 = ~n1784 & n1795;
  assign n1797 = ~n1783 & n1796;
  assign y6 = ~n1673 & n1797;
  assign n1799 = ~q2 & ~n442;
  assign n1800 = q2 & n442;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = ~n465 & n1801;
  assign n1803 = ~r2 & ~n1802;
  assign n1804 = r2 & n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign y7 = n446 & n1805;
  assign n1807 = ~n505 & ~n550;
  assign n1808 = ~n550 & ~n563;
  assign n1809 = n505 & ~n563;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1807 & n1810;
  assign n1812 = ~n533 & n1811;
  assign n1813 = ~r3 & ~n1812;
  assign n1814 = r3 & n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign y8 = n509 & n1815;
  assign n1817 = ~r4 & n1308;
  assign n1818 = r4 & ~n1308;
  assign n1819 = ~n1817 & ~n1818;
  assign y9 = n1304 & n1819;
  assign n1821 = k0 & r3;
  assign n1822 = l0 & n3;
  assign n1823 = g3 & m0;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~n1821 & n1824;
  assign n1826 = a4 & n0;
  assign n1827 = o0 & x3;
  assign n1828 = p0 & u3;
  assign n1829 = n4 & q0;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~n1827 & n1830;
  assign n1832 = ~n1826 & n1831;
  assign n1833 = j4 & r0;
  assign n1834 = e4 & s0;
  assign n1835 = t0 & x4;
  assign n1836 = s4 & u0;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1834 & n1837;
  assign n1839 = ~n1833 & n1838;
  assign n1840 = n1832 & n1839;
  assign z5 = ~n1825 | ~n1840;
  assign n1842 = ~s1 & ~n404;
  assign n1843 = s1 & n404;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n434 & n1844;
  assign n1846 = ~w2 & n1844;
  assign n1847 = ~w2 & n434;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1845 & n1848;
  assign z6 = ~b & n1849;
  assign n1851 = n471 & n476;
  assign n1852 = ~n442 & n471;
  assign n1853 = n442 & n476;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1851 & n1854;
  assign n1856 = ~n465 & n1855;
  assign n1857 = ~s2 & ~n1856;
  assign n1858 = s2 & n1856;
  assign n1859 = ~n1857 & ~n1858;
  assign z7 = n446 & n1859;
  assign n1861 = r3 & n550;
  assign n1862 = ~n505 & ~n1861;
  assign n1863 = ~n564 & ~n1861;
  assign n1864 = n505 & ~n564;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1862 & n1865;
  assign n1867 = ~n533 & n1866;
  assign n1868 = ~s3 & n1867;
  assign n1869 = s3 & ~n1867;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = n509 & ~n1870;
  assign z8 = n510 | n1871;
  assign n1873 = ~s4 & ~n1818;
  assign n1874 = s4 & n1818;
  assign n1875 = ~n1873 & ~n1874;
  assign z9 = n1304 & n1875;
  assign n1877 = t4 & n1309;
  assign n1878 = ~n1308 & n1877;
  assign n1879 = ~u4 & ~n1878;
  assign n1880 = u4 & n1878;
  assign n1881 = ~n1879 & ~n1880;
  assign b10 = n1304 & n1881;
  assign n1883 = u4 & n1877;
  assign n1884 = ~n1308 & n1883;
  assign n1885 = ~v4 & ~n1884;
  assign n1886 = v4 & n1884;
  assign n1887 = ~n1885 & ~n1886;
  assign c10 = n1304 & n1887;
  assign n1889 = v4 & n1883;
  assign n1890 = ~n1308 & n1889;
  assign n1891 = ~w4 & ~n1890;
  assign n1892 = w4 & n1890;
  assign n1893 = ~n1891 & ~n1892;
  assign d10 = n1304 & n1893;
  assign n1895 = w4 & n1889;
  assign n1896 = ~n1308 & n1895;
  assign n1897 = ~x4 & ~n1896;
  assign n1898 = x4 & n1896;
  assign n1899 = ~n1897 & ~n1898;
  assign e10 = n1304 & n1899;
  assign n1901 = v4 & w4;
  assign n1902 = x4 & n1901;
  assign n1903 = n1883 & n1902;
  assign n1904 = ~n1308 & n1903;
  assign n1905 = ~y4 & ~n1904;
  assign n1906 = y4 & n1904;
  assign n1907 = ~n1905 & ~n1906;
  assign f10 = n1304 & n1907;
  assign n1909 = y4 & ~n1308;
  assign n1910 = n1903 & n1909;
  assign n1911 = z4 & n1910;
  assign n1912 = ~z4 & ~n1910;
  assign n1913 = ~n1911 & ~n1912;
  assign g10 = n1304 & n1913;
  assign n1915 = ~z & ~n1191;
  assign n1916 = ~n494 & n1915;
  assign n1917 = ~d5 & n1915;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = d5 & ~n1918;
  assign k10 = n512 | n1919;
  assign n1921 = ~e5 & n1915;
  assign n1922 = ~n493 & n1915;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = e5 & ~n1923;
  assign l10 = n499 | n1924;
  assign n1926 = ~n644 & ~n1191;
  assign n1927 = ~f5 & ~g5;
  assign n1928 = h5 & n603;
  assign n1929 = ~h5 & ~n603;
  assign n1930 = ~z & ~n1929;
  assign n1931 = ~n1928 & n1930;
  assign o10 = ~n1926 | n1931;
  assign n1933 = ~h5 & o10;
  assign n1934 = ~z & n1933;
  assign n1935 = ~n1927 & n1934;
  assign n1936 = ~z & ~f5;
  assign n1937 = ~n1927 & n1936;
  assign n1938 = ~n1933 & n1936;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~n1935 & n1939;
  assign m10 = n1926 & n1940;
  assign n1942 = ~f5 & n1933;
  assign n1943 = n1926 & n1942;
  assign n1944 = ~g5 & ~n1933;
  assign n1945 = n1926 & n1944;
  assign n1946 = n1926 & n1927;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1943 & n1947;
  assign n10 = ~z & n1948;
  assign n1950 = ~z & ~n524;
  assign n1951 = j5 & n535;
  assign n1952 = ~j5 & ~n535;
  assign n1953 = ~n1951 & ~n1952;
  assign q10 = n1950 & n1953;
  assign n1955 = ~k5 & ~n1951;
  assign n1956 = k5 & n1951;
  assign n1957 = ~n1955 & ~n1956;
  assign r10 = n1950 & n1957;
  assign n1959 = n494 & n508;
  assign n1960 = n494 & ~n582;
  assign n1961 = n588 & n1960;
  assign n1962 = n535 & ~n1961;
  assign n1963 = ~n644 & ~n1962;
  assign n1964 = ~n1959 & n1963;
  assign s10 = ~z & ~n1964;
  assign n1966 = ~m5 & n582;
  assign n1967 = ~n317 & n1966;
  assign n1968 = ~m5 & n494;
  assign n1969 = ~n317 & n1968;
  assign n1970 = ~m5 & ~n535;
  assign n1971 = ~n317 & n1970;
  assign n1972 = ~n5 & n582;
  assign n1973 = ~n317 & n1972;
  assign n1974 = ~n5 & n494;
  assign n1975 = ~n317 & n1974;
  assign n1976 = ~n5 & ~n535;
  assign n1977 = ~n317 & n1976;
  assign n1978 = ~n1975 & ~n1977;
  assign n1979 = ~n1973 & n1978;
  assign n1980 = ~n1971 & n1979;
  assign n1981 = ~n1969 & n1980;
  assign n1982 = ~n1967 & n1981;
  assign n1983 = n535 & n582;
  assign n1984 = ~a0 & r5;
  assign n1985 = ~n1911 & n1984;
  assign n1986 = ~a0 & ~z4;
  assign n1987 = ~r5 & n1986;
  assign n1988 = ~n1911 & n1986;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1985 & n1989;
  assign n1991 = v10 & n1990;
  assign n1992 = ~n1983 & ~n1991;
  assign n1993 = ~n508 & n1992;
  assign n1994 = ~n313 & n1993;
  assign n1995 = ~n1982 & n1994;
  assign t10 = ~z & ~n1995;
  assign n1997 = ~n317 & ~n588;
  assign n1998 = ~n317 & n582;
  assign n1999 = ~n317 & ~n494;
  assign n2000 = ~n317 & ~n535;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = ~n1998 & n2001;
  assign n2003 = ~n1997 & n2002;
  assign n2004 = ~n582 & ~n644;
  assign n2005 = ~n313 & n2004;
  assign n2006 = ~n535 & ~n644;
  assign n2007 = ~n313 & n2006;
  assign n2008 = ~n2005 & ~n2007;
  assign n2009 = ~n2003 & ~n2008;
  assign u10 = ~z & ~n2009;
  assign n2011 = ~q5 & n318;
  assign n2012 = ~n314 & n2011;
  assign n2013 = ~n314 & n327;
  assign n2014 = ~r5 & ~n318;
  assign n2015 = n314 & n2014;
  assign n2016 = n314 & n319;
  assign n2017 = n314 & n330;
  assign n2018 = ~n318 & n327;
  assign n2019 = n318 & n321;
  assign n2020 = ~n332 & ~n2019;
  assign n2021 = ~n2018 & n2020;
  assign n2022 = ~n2017 & n2021;
  assign n2023 = ~n2016 & n2022;
  assign n2024 = ~n2015 & n2023;
  assign n2025 = ~n2013 & n2024;
  assign n2026 = ~n2012 & n2025;
  assign w10 = n349 | n2026;
  assign n2028 = ~n314 & n325;
  assign n2029 = ~n314 & n330;
  assign n2030 = ~p5 & ~n318;
  assign n2031 = n314 & n2030;
  assign n2032 = n314 & n2011;
  assign n2033 = n314 & n321;
  assign n2034 = ~n318 & n330;
  assign n2035 = n318 & n327;
  assign n2036 = ~n332 & ~n2035;
  assign n2037 = ~n2034 & n2036;
  assign n2038 = ~n2033 & n2037;
  assign n2039 = ~n2032 & n2038;
  assign n2040 = ~n2031 & n2039;
  assign n2041 = ~n2029 & n2040;
  assign n2042 = ~n2028 & n2041;
  assign x10 = ~n349 & n2042;
  assign l6 = a;
  assign m6 = e1;
  assign r6 = j1;
  assign h10 = y;
  assign i10 = a5;
  assign p10 = g5;
endmodule


