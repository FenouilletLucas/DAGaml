// Benchmark "apex6" written by ABC on Tue May 16 16:07:44 2017

module apex6 ( 
    A, B, C, STW_N, QPR0, QPR1, QPR2, QPR3, QPR4, ENWIN, INZZZE, XZFR0,
    XZFR1, VZZZE, RXZ0, RXZ1, INFIN, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, XZ161, XZ162, XZ163, I2ZZZ0, I2ZZZ1,
    I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, XZ160_N, I2ZZZ7, TXMESS_N,
    PZZZE, RYZ, AXZ0, AXZ1, COMPPAR, MMERR, V1ZZZ0, PSRW, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3,
    I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, RPTEN, XZ320, XZ321, XZ322, XZ323,
    XZ324, CBT0, CBT1, CBT2, ESRSUM, SLAD0, SLAD1, SLAD2, SLAD3, XZFS,
    RPTWIN, PFIN, PSYNC, OFS1, OFS2, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3,
    P2ZZZ4, TXWRD0, P2ZZZ5, TXWRD1, P2ZZZ6, TXWRD2, P2ZZZ7, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, INYBB0, INYBB1, INYBB2, INYBB3,
    INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, VYBB0, VYBB1, TXWRD10, TXWRD11,
    TXWRD12, TXWRD13, TXWRD14, TXWRD15, PYBB0, PYBB1, PYBB2, PYBB3, PYBB4,
    PYBB5, PYBB6, PYBB7, PYBB8, ICLR, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3,
    P1ZZZ4, P1ZZZ5, P1ZZZ6, P1ZZZ7, VFIN,
    V2ZZZ2_P, QPR3_P, XZ323_P, P1ZZZ4_P, I1ZZZ3_P, TXWRD5_P, STW_F,
    TXWRD13_P, V1ZZZ4_P, P2ZZZ1_P, I2ZZZ2_P, TXWRD0_P, A_P, V2ZZZ1_P,
    TXWRD8_P, QPR4_P, XZ324_P, P1ZZZ3_P, I1ZZZ4_P, V1ZZZ3_P, COMPPAR_P,
    XZFS_P, P2ZZZ4_P, I2ZZZ3_P, XZ160_F, B_P, TXMESS_F, TXWRD7_P, P1ZZZ6_P,
    V2ZZZ4_P, I1ZZZ5_P, TXWRD15_P, V1ZZZ6_P, XZ161_P, RPTWIN_P, P2ZZZ3_P,
    AXZ0_P, I2ZZZ4_P, TXWRD2_P, C_P, P1ZZZ5_P, V2ZZZ3_P, I1ZZZ6_P, FSESR_P,
    V1ZZZ5_P, XZ162_P, TXWRD10_P, P1ZZZ0_P, OFS1_P, P2ZZZ6_P, AXZ1_P,
    I2ZZZ5_P, TXWRD1_P, I1ZZZ7_P, TXWRD9_P, ENWIN_P, V1ZZZ0_P, V2ZZZ6_P,
    XZ163_P, OFS2_P, P2ZZZ5_P, I1ZZZ0_P, I2ZZZ6_P, QPR0_P, XZ320_P,
    P1ZZZ7_P, TXWRD4_P, RXZ0_P, V2ZZZ5_P, SBUFF, V1ZZZ7_P, P2ZZZ0_P,
    TXWRD12_P, I2ZZZ7_P, P1ZZZ2_P, V2ZZZ0_P, I1ZZZ1_P, QPR1_P, XZ321_P,
    TXWRD3_P, RXZ1_P, V1ZZZ2_P, XZFR0_P, TD_P, I2ZZZ0_P, P2ZZZ7_P,
    TXWRD11_P, P1ZZZ1_P, I1ZZZ2_P, RYZ_P, QPR2_P, XZ322_P, V2ZZZ7_P,
    TXWRD6_P, V1ZZZ1_P, XZFR1_P, TXWRD14_P, P2ZZZ2_P, I2ZZZ1_P  );
  input  A, B, C, STW_N, QPR0, QPR1, QPR2, QPR3, QPR4, ENWIN, INZZZE,
    XZFR0, XZFR1, VZZZE, RXZ0, RXZ1, INFIN, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, XZ161, XZ162, XZ163, I2ZZZ0, I2ZZZ1,
    I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, XZ160_N, I2ZZZ7, TXMESS_N,
    PZZZE, RYZ, AXZ0, AXZ1, COMPPAR, MMERR, V1ZZZ0, PSRW, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3,
    I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, RPTEN, XZ320, XZ321, XZ322, XZ323,
    XZ324, CBT0, CBT1, CBT2, ESRSUM, SLAD0, SLAD1, SLAD2, SLAD3, XZFS,
    RPTWIN, PFIN, PSYNC, OFS1, OFS2, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3,
    P2ZZZ4, TXWRD0, P2ZZZ5, TXWRD1, P2ZZZ6, TXWRD2, P2ZZZ7, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, INYBB0, INYBB1, INYBB2, INYBB3,
    INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, VYBB0, VYBB1, TXWRD10, TXWRD11,
    TXWRD12, TXWRD13, TXWRD14, TXWRD15, PYBB0, PYBB1, PYBB2, PYBB3, PYBB4,
    PYBB5, PYBB6, PYBB7, PYBB8, ICLR, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3,
    P1ZZZ4, P1ZZZ5, P1ZZZ6, P1ZZZ7, VFIN;
  output V2ZZZ2_P, QPR3_P, XZ323_P, P1ZZZ4_P, I1ZZZ3_P, TXWRD5_P, STW_F,
    TXWRD13_P, V1ZZZ4_P, P2ZZZ1_P, I2ZZZ2_P, TXWRD0_P, A_P, V2ZZZ1_P,
    TXWRD8_P, QPR4_P, XZ324_P, P1ZZZ3_P, I1ZZZ4_P, V1ZZZ3_P, COMPPAR_P,
    XZFS_P, P2ZZZ4_P, I2ZZZ3_P, XZ160_F, B_P, TXMESS_F, TXWRD7_P, P1ZZZ6_P,
    V2ZZZ4_P, I1ZZZ5_P, TXWRD15_P, V1ZZZ6_P, XZ161_P, RPTWIN_P, P2ZZZ3_P,
    AXZ0_P, I2ZZZ4_P, TXWRD2_P, C_P, P1ZZZ5_P, V2ZZZ3_P, I1ZZZ6_P, FSESR_P,
    V1ZZZ5_P, XZ162_P, TXWRD10_P, P1ZZZ0_P, OFS1_P, P2ZZZ6_P, AXZ1_P,
    I2ZZZ5_P, TXWRD1_P, I1ZZZ7_P, TXWRD9_P, ENWIN_P, V1ZZZ0_P, V2ZZZ6_P,
    XZ163_P, OFS2_P, P2ZZZ5_P, I1ZZZ0_P, I2ZZZ6_P, QPR0_P, XZ320_P,
    P1ZZZ7_P, TXWRD4_P, RXZ0_P, V2ZZZ5_P, SBUFF, V1ZZZ7_P, P2ZZZ0_P,
    TXWRD12_P, I2ZZZ7_P, P1ZZZ2_P, V2ZZZ0_P, I1ZZZ1_P, QPR1_P, XZ321_P,
    TXWRD3_P, RXZ1_P, V1ZZZ2_P, XZFR0_P, TD_P, I2ZZZ0_P, P2ZZZ7_P,
    TXWRD11_P, P1ZZZ1_P, I1ZZZ2_P, RYZ_P, QPR2_P, XZ322_P, V2ZZZ7_P,
    TXWRD6_P, V1ZZZ1_P, XZFR1_P, TXWRD14_P, P2ZZZ2_P, I2ZZZ1_P;
  wire n235, n236, n237, n238, n239, n241, n242, n243, n244, n245, n246,
    n248, n249, n250, n251, n252, n253, n255, n256, n257, n259, n260, n261,
    n262, n263, n264, n265, n267, n268, n269, n270, n271, n273, n274, n275,
    n276, n277, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n297, n298, n299, n300, n301,
    n302, n304, n305, n306, n307, n308, n309, n310, n311, n312, n314, n315,
    n316, n317, n318, n320, n321, n322, n323, n324, n326, n327, n328, n329,
    n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n355, n356,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n368, n369, n370,
    n371, n372, n373, n375, n376, n377, n378, n379, n380, n381, n382, n384,
    n385, n387, n388, n390, n391, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n432, n434, n435, n436, n438,
    n439, n441, n442, n444, n445, n446, n447, n448, n449, n450, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n477, n478, n480,
    n481, n483, n484, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n496, n497, n499, n500, n501, n502, n503, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n533, n534,
    n536, n537, n538, n539, n540, n542, n543, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561, n562,
    n563, n565, n566, n568, n569, n571, n572, n575, n576, n578, n579, n581,
    n582, n583, n584, n585, n586, n587, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n600, n601, n603, n604, n606, n607, n608, n609,
    n611, n612, n614, n615, n616, n617, n618, n619, n620, n621, n622, n624,
    n625, n627, n628, n629, n630, n631, n632, n633, n634, n635, n637, n638,
    n639, n640, n642, n643, n645, n646, n648, n649, n650, n651, n652, n653,
    n654, n656, n657, n659, n660, n662, n663, n665, n666, n667, n669, n670,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n726, n727, n730, n731, n733, n734, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n747, n748, n750, n751,
    n753, n754, n756, n757, n759, n760, n761, n763, n764, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n776, n777, n778, n779, n780, n781,
    n783, n784, n786, n787, n788, n789, n790, n791, n792, n793, n794, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n823, n824, n826, n827, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n840, n841, n843, n844, n847, n848, n849, n851, n852,
    n853, n855, n856, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n868, n869, n871, n872, n873, n874, n875, n876, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n888, n889, n891, n892;
  assign n235 = VZZZE & VYBB0;
  assign n236 = ~RYZ & n235;
  assign n237 = ~RYZ & ~n235;
  assign n238 = V2ZZZ3 & n236;
  assign n239 = V2ZZZ2 & n237;
  assign V2ZZZ2_P = n238 | n239;
  assign n241 = ~INFIN & ~PFIN;
  assign n242 = TXMESS_N & ~VFIN;
  assign n243 = n241 & n242;
  assign n244 = QPR0 & ~n243;
  assign n245 = QPR1 & n244;
  assign n246 = QPR2 & n245;
  assign TXMESS_F = RYZ | n243;
  assign n248 = QPR0 & QPR1;
  assign n249 = ~TXMESS_F & n248;
  assign n250 = QPR3 & ~n246;
  assign n251 = ~RYZ & n250;
  assign n252 = QPR2 & ~QPR3;
  assign n253 = n249 & n252;
  assign QPR3_P = n251 | n253;
  assign n255 = XZ321 & XZ322;
  assign n256 = ~PSYNC & ~ICLR;
  assign n257 = XZ320 & n256;
  assign XZ320_P = ~XZ320 & n256;
  assign n259 = ~XZ321 & n256;
  assign n260 = ~XZ320_P & ~n259;
  assign n261 = ~XZ322 & n256;
  assign n262 = n260 & ~n261;
  assign n263 = XZ323 & ~n262;
  assign n264 = ~XZ323 & n257;
  assign n265 = n255 & n264;
  assign XZ323_P = n263 | n265;
  assign n267 = ~PZZZE & PYBB0;
  assign n268 = ~RYZ & n267;
  assign n269 = ~RYZ & ~n267;
  assign n270 = PYBB5 & n268;
  assign n271 = P1ZZZ4 & n269;
  assign P1ZZZ4_P = n270 | n271;
  assign n273 = ~INZZZE & INYBB0;
  assign n274 = ~RYZ & n273;
  assign n275 = ~RYZ & ~n273;
  assign n276 = INYBB4 & n274;
  assign n277 = I1ZZZ3 & n275;
  assign I1ZZZ3_P = n276 | n277;
  assign n279 = ~INFIN & ~RYZ;
  assign n280 = ~PFIN & n279;
  assign n281 = ~B & ~C;
  assign n282 = ~TXMESS_N & ~n281;
  assign n283 = ~VFIN & n282;
  assign n284 = ~VFIN & ~n282;
  assign n285 = TXWRD6 & n283;
  assign n286 = TXWRD5 & n284;
  assign n287 = V1ZZZ5 & VFIN;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~n285 & n288;
  assign n290 = PFIN & n279;
  assign n291 = INFIN & ~RYZ;
  assign n292 = n280 & ~n289;
  assign n293 = P1ZZZ5 & n290;
  assign n294 = I1ZZZ5 & n291;
  assign n295 = ~n293 & ~n294;
  assign TXWRD5_P = n292 | ~n295;
  assign n297 = ~TXMESS_N & AXZ0;
  assign n298 = AXZ1 & n297;
  assign n299 = A & n298;
  assign n300 = ~STW_N & ~n299;
  assign n301 = ~VFIN & n241;
  assign n302 = ~n300 & n301;
  assign STW_F = RYZ | n302;
  assign n304 = TXWRD14 & n283;
  assign n305 = TXWRD13 & n284;
  assign n306 = V2ZZZ5 & VFIN;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~n304 & n307;
  assign n309 = n280 & ~n308;
  assign n310 = I2ZZZ5 & n291;
  assign n311 = P2ZZZ5 & n290;
  assign n312 = ~n310 & ~n311;
  assign TXWRD13_P = n309 | ~n312;
  assign n314 = ~VZZZE & VYBB0;
  assign n315 = ~RYZ & n314;
  assign n316 = ~RYZ & ~n314;
  assign n317 = V1ZZZ5 & n315;
  assign n318 = V1ZZZ4 & n316;
  assign V1ZZZ4_P = n317 | n318;
  assign n320 = PZZZE & PYBB0;
  assign n321 = ~RYZ & n320;
  assign n322 = ~RYZ & ~n320;
  assign n323 = PYBB2 & n321;
  assign n324 = P2ZZZ1 & n322;
  assign P2ZZZ1_P = n323 | n324;
  assign n326 = INZZZE & INYBB0;
  assign n327 = ~RYZ & n326;
  assign n328 = ~RYZ & ~n326;
  assign n329 = INYBB3 & n327;
  assign n330 = I2ZZZ2 & n328;
  assign I2ZZZ2_P = n329 | n330;
  assign n332 = ~INFIN & PFIN;
  assign n333 = TXWRD1 & n283;
  assign n334 = TXWRD0 & n284;
  assign n335 = V1ZZZ0 & VFIN;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~n333 & n336;
  assign n338 = P1ZZZ0 & n332;
  assign n339 = n241 & ~n337;
  assign n340 = INFIN & I1ZZZ0;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~n338 & n341;
  assign TXWRD0_P = ~RYZ & ~n342;
  assign n344 = B & ~QPR4;
  assign n345 = ~QPR4 & CBT2;
  assign n346 = QPR3 & n344;
  assign n347 = ~QPR3 & ~n345;
  assign n348 = ~n346 & ~n347;
  assign n349 = QPR0 & ~QPR1;
  assign n350 = QPR2 & n349;
  assign n351 = ~n348 & n350;
  assign n352 = ~TXMESS_N & n351;
  assign n353 = ~A & ~n352;
  assign A_P = ~RYZ & ~n353;
  assign n355 = V2ZZZ2 & n236;
  assign n356 = V2ZZZ1 & n237;
  assign V2ZZZ1_P = n355 | n356;
  assign n358 = TXWRD9 & n283;
  assign n359 = TXWRD8 & n284;
  assign n360 = V2ZZZ0 & VFIN;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n358 & n361;
  assign n363 = n280 & ~n362;
  assign n364 = P2ZZZ0 & n290;
  assign n365 = I2ZZZ0 & n291;
  assign n366 = ~n364 & ~n365;
  assign TXWRD8_P = n363 | ~n366;
  assign n368 = QPR3 & n246;
  assign n369 = QPR2 & QPR3;
  assign n370 = ~QPR4 & n369;
  assign n371 = n249 & n370;
  assign n372 = QPR4 & ~n368;
  assign n373 = ~RYZ & n372;
  assign QPR4_P = n371 | n373;
  assign n375 = XZ320 & XZ323;
  assign n376 = n255 & n375;
  assign n377 = XZ322 & XZ323;
  assign n378 = n256 & ~n377;
  assign n379 = n260 & ~n378;
  assign n380 = XZ324 & ~n379;
  assign n381 = ~XZ324 & n376;
  assign n382 = n256 & n381;
  assign XZ324_P = n380 | n382;
  assign n384 = PYBB4 & n268;
  assign n385 = P1ZZZ3 & n269;
  assign P1ZZZ3_P = n384 | n385;
  assign n387 = INYBB5 & n274;
  assign n388 = I1ZZZ4 & n275;
  assign I1ZZZ4_P = n387 | n388;
  assign n390 = V1ZZZ4 & n315;
  assign n391 = V1ZZZ3 & n316;
  assign V1ZZZ3_P = n390 | n391;
  assign n393 = ~AXZ0 & ~AXZ1;
  assign n394 = A & ~n393;
  assign n395 = ~QPR0 & SLAD1;
  assign n396 = QPR0 & SLAD0;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~QPR0 & SLAD3;
  assign n399 = QPR0 & SLAD2;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~QPR1 & QPR2;
  assign n402 = ~n397 & n401;
  assign n403 = QPR1 & ~QPR2;
  assign n404 = ~n400 & n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = TXWRD0 & ~n281;
  assign n407 = ~QPR3 & n281;
  assign n408 = ~QPR4 & n407;
  assign n409 = ~n405 & n408;
  assign n410 = ~n406 & ~n409;
  assign n411 = ~n394 & n410;
  assign n412 = ~TXMESS_N & ~n411;
  assign n413 = AXZ1 & ESRSUM;
  assign n414 = AXZ0 & ~MMERR;
  assign n415 = ~n413 & ~n414;
  assign n416 = AXZ0 & MMERR;
  assign n417 = AXZ1 & ~ESRSUM;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~TXMESS_N & ~n415;
  assign n420 = ~COMPPAR & n419;
  assign n421 = COMPPAR & ~n418;
  assign n422 = ~n298 & ~n421;
  assign n423 = ~n420 & n422;
  assign n424 = ~n394 & ~n410;
  assign n425 = ~TXMESS_N & n424;
  assign n426 = ~COMPPAR & n425;
  assign n427 = A & ~n423;
  assign n428 = COMPPAR & ~n412;
  assign n429 = ~n427 & ~n428;
  assign n430 = ~n426 & n429;
  assign COMPPAR_P = ~RYZ & ~n430;
  assign n432 = OFS1 & OFS2;
  assign OFS1_P = PSYNC & ~ICLR;
  assign n434 = XZFS & ~ICLR;
  assign n435 = ~OFS1_P & ~n434;
  assign n436 = PSRW & ~n435;
  assign XZFS_P = ~n432 & n436;
  assign n438 = PYBB5 & n321;
  assign n439 = P2ZZZ4 & n322;
  assign P2ZZZ4_P = n438 | n439;
  assign n441 = INYBB4 & n327;
  assign n442 = I2ZZZ3 & n328;
  assign I2ZZZ3_P = n441 | n442;
  assign n444 = XZ323 & XZ324;
  assign n445 = n255 & n444;
  assign n446 = ~XZ160_N & n445;
  assign n447 = n256 & ~n445;
  assign n448 = ~XZ320_P & ~n447;
  assign n449 = XZ160_N & ~n448;
  assign n450 = n257 & n446;
  assign XZ160_F = n449 | n450;
  assign n452 = ~CBT0 & ~CBT1;
  assign n453 = CBT2 & ~n452;
  assign n454 = ~QPR3 & ~n453;
  assign n455 = ~TXMESS_N & n350;
  assign n456 = ~QPR4 & n455;
  assign n457 = ~n454 & n456;
  assign n458 = n350 & n453;
  assign n459 = ~B & n458;
  assign n460 = ~QPR3 & n459;
  assign n461 = ~QPR4 & n460;
  assign n462 = ~TXMESS_N & n461;
  assign n463 = B & ~n457;
  assign n464 = ~n462 & ~n463;
  assign B_P = ~RYZ & ~n464;
  assign n466 = TXWRD8 & n283;
  assign n467 = TXWRD7 & n284;
  assign n468 = V1ZZZ7 & VFIN;
  assign n469 = ~n467 & ~n468;
  assign n470 = ~n466 & n469;
  assign n471 = P1ZZZ7 & n332;
  assign n472 = INFIN & I1ZZZ7;
  assign n473 = n241 & ~n470;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n471 & n474;
  assign TXWRD7_P = ~RYZ & ~n475;
  assign n477 = PYBB7 & n268;
  assign n478 = P1ZZZ6 & n269;
  assign P1ZZZ6_P = n477 | n478;
  assign n480 = V2ZZZ5 & n236;
  assign n481 = V2ZZZ4 & n237;
  assign V2ZZZ4_P = n480 | n481;
  assign n483 = INYBB6 & n274;
  assign n484 = I1ZZZ5 & n275;
  assign I1ZZZ5_P = n483 | n484;
  assign n486 = ~PFIN & VFIN;
  assign n487 = ~PFIN & n284;
  assign n488 = V2ZZZ7 & n486;
  assign n489 = TXWRD15 & n487;
  assign n490 = PFIN & P2ZZZ7;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~n488 & n491;
  assign n493 = n279 & ~n492;
  assign n494 = I2ZZZ7 & n291;
  assign TXWRD15_P = n493 | n494;
  assign n496 = V1ZZZ7 & n315;
  assign n497 = V1ZZZ6 & n316;
  assign V1ZZZ6_P = n496 | n497;
  assign n499 = n256 & ~n446;
  assign n500 = ~XZ320_P & ~n499;
  assign n501 = XZ161 & ~n500;
  assign n502 = ~XZ161 & n446;
  assign n503 = n257 & n502;
  assign XZ161_P = n501 | n503;
  assign n505 = ~SLAD2 & ~SLAD3;
  assign n506 = PSYNC & n505;
  assign n507 = XZFS & n506;
  assign n508 = RXZ0 & RXZ1;
  assign n509 = ~XZ160_N & SLAD0;
  assign n510 = XZ160_N & ~SLAD0;
  assign n511 = ~n509 & ~n510;
  assign n512 = XZ161 & SLAD1;
  assign n513 = ~XZ161 & ~SLAD1;
  assign n514 = ~n512 & ~n513;
  assign n515 = XZ162 & SLAD2;
  assign n516 = ~XZ162 & ~SLAD2;
  assign n517 = ~n515 & ~n516;
  assign n518 = XZ163 & SLAD3;
  assign n519 = ~XZ163 & ~SLAD3;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n517 & ~n520;
  assign n522 = ENWIN & XZ324;
  assign n523 = n376 & n522;
  assign n524 = n521 & n523;
  assign n525 = ~n514 & n524;
  assign n526 = ~n511 & n525;
  assign n527 = ~SLAD0 & ~SLAD1;
  assign n528 = n507 & n527;
  assign n529 = RPTWIN & ~n508;
  assign n530 = ~n526 & ~n529;
  assign n531 = ~n528 & n530;
  assign RPTWIN_P = ~RYZ & ~n531;
  assign n533 = PYBB4 & n321;
  assign n534 = P2ZZZ3 & n322;
  assign P2ZZZ3_P = n533 | n534;
  assign n536 = ~A & ~n351;
  assign n537 = ~TXMESS_N & ~n536;
  assign n538 = AXZ0 & ~n537;
  assign n539 = ~AXZ0 & n537;
  assign n540 = ~n538 & ~n539;
  assign AXZ0_P = ~RYZ & ~n540;
  assign n542 = INYBB5 & n327;
  assign n543 = I2ZZZ4 & n328;
  assign I2ZZZ4_P = n542 | n543;
  assign n545 = ~PFIN & n283;
  assign n546 = V1ZZZ2 & n486;
  assign n547 = TXWRD3 & n545;
  assign n548 = TXWRD2 & n487;
  assign n549 = PFIN & P1ZZZ2;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n547 & n550;
  assign n552 = ~n546 & n551;
  assign n553 = I1ZZZ2 & n291;
  assign n554 = n279 & ~n552;
  assign TXWRD2_P = n553 | n554;
  assign n556 = CBT2 & n452;
  assign n557 = ~QPR4 & ~n556;
  assign n558 = ~QPR3 & n350;
  assign n559 = ~TXMESS_N & n558;
  assign n560 = ~n557 & n559;
  assign n561 = C & ~n560;
  assign n562 = ~C & n560;
  assign n563 = ~n561 & ~n562;
  assign C_P = ~RYZ & ~n563;
  assign n565 = PYBB6 & n268;
  assign n566 = P1ZZZ5 & n269;
  assign P1ZZZ5_P = n565 | n566;
  assign n568 = V2ZZZ4 & n236;
  assign n569 = V2ZZZ3 & n237;
  assign V2ZZZ3_P = n568 | n569;
  assign n571 = INYBB7 & n274;
  assign n572 = I1ZZZ6 & n275;
  assign I1ZZZ6_P = n571 | n572;
  assign OFS2_P = OFS1 & ~ICLR;
  assign n575 = OFS2 & OFS2_P;
  assign n576 = XZFR1 & ~ICLR;
  assign FSESR_P = n575 | n576;
  assign n578 = V1ZZZ6 & n315;
  assign n579 = V1ZZZ5 & n316;
  assign V1ZZZ5_P = n578 | n579;
  assign n581 = XZ161 & XZ320;
  assign n582 = n446 & n581;
  assign n583 = ~XZ161 & n256;
  assign n584 = n500 & ~n583;
  assign n585 = ~XZ162 & n582;
  assign n586 = n256 & n585;
  assign n587 = XZ162 & ~n584;
  assign XZ162_P = n586 | n587;
  assign n589 = TXWRD11 & n283;
  assign n590 = TXWRD10 & n284;
  assign n591 = V2ZZZ2 & VFIN;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n589 & n592;
  assign n594 = INFIN & I2ZZZ2;
  assign n595 = n241 & ~n593;
  assign n596 = P2ZZZ2 & n332;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n594 & n597;
  assign TXWRD10_P = ~RYZ & ~n598;
  assign n600 = PYBB1 & n268;
  assign n601 = P1ZZZ0 & n269;
  assign P1ZZZ0_P = n600 | n601;
  assign n603 = PYBB7 & n321;
  assign n604 = P2ZZZ6 & n322;
  assign P2ZZZ6_P = n603 | n604;
  assign n606 = AXZ0 & n537;
  assign n607 = ~AXZ1 & n606;
  assign n608 = AXZ1 & ~n606;
  assign n609 = ~n607 & ~n608;
  assign AXZ1_P = ~RYZ & ~n609;
  assign n611 = INYBB6 & n327;
  assign n612 = I2ZZZ5 & n328;
  assign I2ZZZ5_P = n611 | n612;
  assign n614 = V1ZZZ1 & n486;
  assign n615 = TXWRD2 & n545;
  assign n616 = TXWRD1 & n487;
  assign n617 = PFIN & P1ZZZ1;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n615 & n618;
  assign n620 = ~n614 & n619;
  assign n621 = n279 & ~n620;
  assign n622 = I1ZZZ1 & n291;
  assign TXWRD1_P = n621 | n622;
  assign n624 = INYBB8 & n274;
  assign n625 = I1ZZZ7 & n275;
  assign I1ZZZ7_P = n624 | n625;
  assign n627 = V2ZZZ1 & n486;
  assign n628 = TXWRD10 & n545;
  assign n629 = TXWRD9 & n487;
  assign n630 = PFIN & P2ZZZ1;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n628 & n631;
  assign n633 = ~n627 & n632;
  assign n634 = n279 & ~n633;
  assign n635 = I2ZZZ1 & n291;
  assign TXWRD9_P = n634 | n635;
  assign n637 = XZFS & OFS1_P;
  assign n638 = ENWIN & ~ICLR;
  assign n639 = ~n637 & ~n638;
  assign n640 = PSRW & ~n639;
  assign ENWIN_P = ~n432 & n640;
  assign n642 = V1ZZZ1 & n315;
  assign n643 = V1ZZZ0 & n316;
  assign V1ZZZ0_P = n642 | n643;
  assign n645 = V2ZZZ7 & n236;
  assign n646 = V2ZZZ6 & n237;
  assign V2ZZZ6_P = n645 | n646;
  assign n648 = XZ161 & XZ162;
  assign n649 = n256 & ~n648;
  assign n650 = n500 & ~n649;
  assign n651 = XZ162 & n582;
  assign n652 = ~XZ163 & n651;
  assign n653 = n256 & n652;
  assign n654 = XZ163 & ~n650;
  assign XZ163_P = n653 | n654;
  assign n656 = PYBB6 & n321;
  assign n657 = P2ZZZ5 & n322;
  assign P2ZZZ5_P = n656 | n657;
  assign n659 = INYBB1 & n274;
  assign n660 = I1ZZZ0 & n275;
  assign I1ZZZ0_P = n659 | n660;
  assign n662 = INYBB7 & n327;
  assign n663 = I2ZZZ6 & n328;
  assign I2ZZZ6_P = n662 | n663;
  assign n665 = QPR0 & ~RYZ;
  assign n666 = n243 & n665;
  assign n667 = ~QPR0 & ~TXMESS_F;
  assign QPR0_P = n666 | n667;
  assign n669 = PYBB8 & n268;
  assign n670 = P1ZZZ7 & n269;
  assign P1ZZZ7_P = n669 | n670;
  assign n672 = TXWRD5 & n283;
  assign n673 = TXWRD4 & n284;
  assign n674 = V1ZZZ4 & VFIN;
  assign n675 = ~n673 & ~n674;
  assign n676 = ~n672 & n675;
  assign n677 = n280 & ~n676;
  assign n678 = P1ZZZ4 & n290;
  assign n679 = I1ZZZ4 & n291;
  assign n680 = ~n678 & ~n679;
  assign TXWRD4_P = n677 | ~n680;
  assign n682 = XZ162 & ~SLAD2;
  assign n683 = XZ163 & ~SLAD3;
  assign n684 = ~n682 & ~n683;
  assign n685 = XZ320 & n684;
  assign n686 = XZ161 & ~SLAD1;
  assign n687 = ENWIN & ~n686;
  assign n688 = n446 & n687;
  assign n689 = n685 & n688;
  assign n690 = ~XZ160_N & ~SLAD0;
  assign n691 = n445 & ~n690;
  assign n692 = n687 & n691;
  assign n693 = XZ163 & ~n682;
  assign n694 = XZ320 & n693;
  assign n695 = n685 & n691;
  assign n696 = XZ161 & n695;
  assign n697 = ENWIN & n696;
  assign n698 = XZ162 & ~n683;
  assign n699 = XZ320 & n698;
  assign n700 = ~XZFS & ~n685;
  assign n701 = SLAD0 & ~n689;
  assign n702 = ~n507 & ~n692;
  assign n703 = ~PSYNC & ~n684;
  assign n704 = SLAD3 & ~n694;
  assign n705 = SLAD1 & ~n697;
  assign n706 = SLAD2 & ~n699;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~n704 & n707;
  assign n709 = ~n703 & n708;
  assign n710 = ~n702 & n709;
  assign n711 = ~n701 & n710;
  assign n712 = ~n700 & n711;
  assign n713 = ~ICLR & ~n712;
  assign n714 = ~XZ320_P & ~n713;
  assign n715 = ~RPTWIN & ~n526;
  assign n716 = ~ICLR & ~n715;
  assign n717 = ~SLAD0 & n637;
  assign n718 = ~SLAD1 & n717;
  assign n719 = ~SLAD2 & n718;
  assign n720 = ~SLAD3 & n719;
  assign n721 = ~n716 & ~n720;
  assign n722 = RXZ0 & ~RPTWIN;
  assign n723 = ~n714 & n722;
  assign n724 = ~RXZ0 & ~n721;
  assign RXZ0_P = n723 | n724;
  assign n726 = V2ZZZ6 & n236;
  assign n727 = V2ZZZ5 & n237;
  assign V2ZZZ5_P = n726 | n727;
  assign SBUFF = ~TXMESS_N | RPTWIN;
  assign n730 = VYBB1 & n315;
  assign n731 = V1ZZZ7 & n316;
  assign V1ZZZ7_P = n730 | n731;
  assign n733 = PYBB1 & n321;
  assign n734 = P2ZZZ0 & n322;
  assign P2ZZZ0_P = n733 | n734;
  assign n736 = TXWRD13 & n283;
  assign n737 = TXWRD12 & n284;
  assign n738 = V2ZZZ4 & VFIN;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = INFIN & I2ZZZ4;
  assign n742 = n241 & ~n740;
  assign n743 = P2ZZZ4 & n332;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n741 & n744;
  assign TXWRD12_P = ~RYZ & ~n745;
  assign n747 = INYBB8 & n327;
  assign n748 = I2ZZZ7 & n328;
  assign I2ZZZ7_P = n747 | n748;
  assign n750 = PYBB3 & n268;
  assign n751 = P1ZZZ2 & n269;
  assign P1ZZZ2_P = n750 | n751;
  assign n753 = V2ZZZ1 & n236;
  assign n754 = V2ZZZ0 & n237;
  assign V2ZZZ0_P = n753 | n754;
  assign n756 = INYBB2 & n274;
  assign n757 = I1ZZZ1 & n275;
  assign I1ZZZ1_P = n756 | n757;
  assign n759 = QPR1 & ~n244;
  assign n760 = ~RYZ & n759;
  assign n761 = ~TXMESS_F & n349;
  assign QPR1_P = n760 | n761;
  assign n763 = XZ321 & XZ320_P;
  assign n764 = ~XZ321 & n257;
  assign XZ321_P = n763 | n764;
  assign n766 = TXWRD4 & n283;
  assign n767 = TXWRD3 & n284;
  assign n768 = V1ZZZ3 & VFIN;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n766 & n769;
  assign n771 = n280 & ~n770;
  assign n772 = P1ZZZ3 & n290;
  assign n773 = I1ZZZ3 & n291;
  assign n774 = ~n772 & ~n773;
  assign TXWRD3_P = n771 | ~n774;
  assign n776 = ~RXZ0 & ~ICLR;
  assign n777 = ~RPTWIN & ~n714;
  assign n778 = ~n776 & ~n777;
  assign n779 = RXZ0 & ~RXZ1;
  assign n780 = ~n721 & n779;
  assign n781 = RXZ1 & ~n778;
  assign RXZ1_P = n780 | n781;
  assign n783 = V1ZZZ3 & n315;
  assign n784 = V1ZZZ2 & n316;
  assign V1ZZZ2_P = n783 | n784;
  assign n786 = ~XZ161 & XZ160_N;
  assign n787 = ~XZ162 & n786;
  assign n788 = ~XZ163 & n787;
  assign n789 = n445 & n788;
  assign n790 = n256 & ~n789;
  assign n791 = ~XZ320_P & ~n790;
  assign n792 = XZFR0 & ~n791;
  assign n793 = ~XZFR0 & n789;
  assign n794 = n257 & n793;
  assign XZFR0_P = n792 | n794;
  assign n796 = ~RPTWIN & n281;
  assign n797 = ~n394 & n796;
  assign n798 = SBUFF & ~n797;
  assign n799 = RXZ0 & ~ESRSUM;
  assign n800 = ~RXZ1 & n799;
  assign n801 = ~RXZ0 & ESRSUM;
  assign n802 = RXZ1 & n801;
  assign n803 = ~n800 & ~n802;
  assign n804 = AXZ0 & ~COMPPAR;
  assign n805 = ~AXZ0 & ESRSUM;
  assign n806 = ~n804 & ~n805;
  assign n807 = ~AXZ1 & n414;
  assign n808 = AXZ1 & ~n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n394 & n406;
  assign n811 = A & ~n809;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~QPR3 & ~n405;
  assign n814 = ~QPR4 & n813;
  assign n815 = ~n798 & n814;
  assign n816 = RPTEN & RPTWIN;
  assign n817 = ~n803 & n816;
  assign n818 = ~RPTWIN & ~n812;
  assign n819 = ~TXMESS_N & n818;
  assign n820 = ~n817 & ~n819;
  assign n821 = ~n815 & n820;
  assign TD_P = ~RYZ & ~n821;
  assign n823 = INYBB1 & n327;
  assign n824 = I2ZZZ0 & n328;
  assign I2ZZZ0_P = n823 | n824;
  assign n826 = PYBB8 & n321;
  assign n827 = P2ZZZ7 & n322;
  assign P2ZZZ7_P = n826 | n827;
  assign n829 = TXWRD12 & n283;
  assign n830 = TXWRD11 & n284;
  assign n831 = V2ZZZ3 & VFIN;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n829 & n832;
  assign n834 = INFIN & I2ZZZ3;
  assign n835 = n241 & ~n833;
  assign n836 = P2ZZZ3 & n332;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~n834 & n837;
  assign TXWRD11_P = ~RYZ & ~n838;
  assign n840 = PYBB2 & n268;
  assign n841 = P1ZZZ1 & n269;
  assign P1ZZZ1_P = n840 | n841;
  assign n843 = INYBB3 & n274;
  assign n844 = I1ZZZ2 & n275;
  assign I1ZZZ2_P = n843 | n844;
  assign RYZ_P = ICLR | n299;
  assign n847 = ~QPR2 & n249;
  assign n848 = QPR2 & ~n245;
  assign n849 = ~RYZ & n848;
  assign QPR2_P = n847 | n849;
  assign n851 = XZ321 & ~XZ322;
  assign n852 = n257 & n851;
  assign n853 = XZ322 & ~n260;
  assign XZ322_P = n852 | n853;
  assign n855 = VYBB1 & n236;
  assign n856 = V2ZZZ7 & n237;
  assign V2ZZZ7_P = n855 | n856;
  assign n858 = TXWRD7 & n283;
  assign n859 = TXWRD6 & n284;
  assign n860 = V1ZZZ6 & VFIN;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n858 & n861;
  assign n863 = n280 & ~n862;
  assign n864 = P1ZZZ6 & n290;
  assign n865 = I1ZZZ6 & n291;
  assign n866 = ~n864 & ~n865;
  assign TXWRD6_P = n863 | ~n866;
  assign n868 = V1ZZZ2 & n315;
  assign n869 = V1ZZZ1 & n316;
  assign V1ZZZ1_P = n868 | n869;
  assign n871 = ~XZFR0 & n256;
  assign n872 = n791 & ~n871;
  assign n873 = XZFR0 & ~XZFR1;
  assign n874 = n257 & n873;
  assign n875 = n789 & n874;
  assign n876 = XZFR1 & ~n872;
  assign XZFR1_P = n875 | n876;
  assign n878 = TXWRD15 & n283;
  assign n879 = TXWRD14 & n284;
  assign n880 = V2ZZZ6 & VFIN;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n878 & n881;
  assign n883 = n280 & ~n882;
  assign n884 = I2ZZZ6 & n291;
  assign n885 = P2ZZZ6 & n290;
  assign n886 = ~n884 & ~n885;
  assign TXWRD14_P = n883 | ~n886;
  assign n888 = PYBB3 & n321;
  assign n889 = P2ZZZ2 & n322;
  assign P2ZZZ2_P = n888 | n889;
  assign n891 = INYBB2 & n327;
  assign n892 = I2ZZZ1 & n328;
  assign I2ZZZ1_P = n891 | n892;
endmodule


