// Benchmark "dalu" written by ABC on Tue May 16 16:07:48 2017

module dalu ( 
    inA10, inA11, inA12, inA13, inA14, inA15, inB10, inB11, inB12, inB13,
    inB14, inB15, inC10, inC11, inC12, inC13, inC14, inC15, inD10, inD11,
    inD12, inD13, inD14, inD15, inA0, inA1, inA2, inA3, inA4, inA5, inA6,
    inA7, inA8, inA9, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7, inB8,
    inB9, inC0, inC1, inC2, inC3, inC4, inC5, inC6, inC7, inC8, inC9, inD0,
    inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, inD9, sh0, sh1, sh2,
    musel1, musel2, musel3, musel4, opsel0, opsel1, opsel2, opsel3,
    O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15  );
  input  inA10, inA11, inA12, inA13, inA14, inA15, inB10, inB11, inB12,
    inB13, inB14, inB15, inC10, inC11, inC12, inC13, inC14, inC15, inD10,
    inD11, inD12, inD13, inD14, inD15, inA0, inA1, inA2, inA3, inA4, inA5,
    inA6, inA7, inA8, inA9, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7,
    inB8, inB9, inC0, inC1, inC2, inC3, inC4, inC5, inC6, inC7, inC8, inC9,
    inD0, inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, inD9, sh0, sh1,
    sh2, musel1, musel2, musel3, musel4, opsel0, opsel1, opsel2, opsel3;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830;
  assign n92 = inC0 & musel2;
  assign n93 = musel1 & ~musel2;
  assign n94 = inA0 & n93;
  assign n95 = ~musel1 & n92;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~musel3 & ~n96;
  assign n98 = musel4 & n97;
  assign n99 = inC15 & musel2;
  assign n100 = inA15 & n93;
  assign n101 = ~musel1 & n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = ~musel3 & ~n102;
  assign n104 = musel4 & n103;
  assign n105 = ~n98 & n104;
  assign n106 = n98 & ~n104;
  assign n107 = ~n105 & ~n106;
  assign n108 = n104 & n107;
  assign n109 = ~n104 & ~n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = opsel2 & ~n110;
  assign n112 = ~opsel0 & ~opsel1;
  assign n113 = n111 & n112;
  assign n114 = musel3 & ~musel4;
  assign n115 = inD4 & musel2;
  assign n116 = ~musel1 & musel2;
  assign n117 = ~n93 & ~n116;
  assign n118 = ~inB4 & ~n115;
  assign n119 = ~inB4 & ~musel1;
  assign n120 = ~n115 & n117;
  assign n121 = ~musel1 & n117;
  assign n122 = ~n120 & ~n121;
  assign n123 = ~n119 & n122;
  assign n124 = ~n118 & n123;
  assign n125 = ~musel1 & ~musel2;
  assign n126 = ~musel3 & n125;
  assign n127 = musel4 & n126;
  assign n128 = inD4 & n127;
  assign n129 = n114 & n124;
  assign n130 = ~n128 & ~n129;
  assign n131 = inD0 & musel2;
  assign n132 = ~inB0 & ~n131;
  assign n133 = ~inB0 & ~musel1;
  assign n134 = n117 & ~n131;
  assign n135 = ~n121 & ~n134;
  assign n136 = ~n133 & n135;
  assign n137 = ~n132 & n136;
  assign n138 = inD0 & n127;
  assign n139 = n114 & n137;
  assign n140 = ~n138 & ~n139;
  assign n141 = sh2 & ~n130;
  assign n142 = ~sh2 & ~n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = inD8 & musel2;
  assign n145 = ~inB8 & ~n144;
  assign n146 = ~inB8 & ~musel1;
  assign n147 = n117 & ~n144;
  assign n148 = ~n121 & ~n147;
  assign n149 = ~n146 & n148;
  assign n150 = ~n145 & n149;
  assign n151 = inD8 & n127;
  assign n152 = n114 & n150;
  assign n153 = ~n151 & ~n152;
  assign n154 = inD2 & musel2;
  assign n155 = ~inB2 & ~n154;
  assign n156 = ~inB2 & ~musel1;
  assign n157 = n117 & ~n154;
  assign n158 = ~n121 & ~n157;
  assign n159 = ~n156 & n158;
  assign n160 = ~n155 & n159;
  assign n161 = inD2 & n127;
  assign n162 = n114 & n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = sh2 & ~n153;
  assign n165 = ~sh2 & ~n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = ~sh1 & n143;
  assign n168 = n143 & n166;
  assign n169 = sh1 & n166;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n167 & n170;
  assign n172 = inD5 & musel2;
  assign n173 = ~inB5 & ~n172;
  assign n174 = ~inB5 & ~musel1;
  assign n175 = n117 & ~n172;
  assign n176 = ~n121 & ~n175;
  assign n177 = ~n174 & n176;
  assign n178 = ~n173 & n177;
  assign n179 = inD5 & n127;
  assign n180 = n114 & n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = inD1 & musel2;
  assign n183 = ~inB1 & ~n182;
  assign n184 = ~inB1 & ~musel1;
  assign n185 = n117 & ~n182;
  assign n186 = ~n121 & ~n185;
  assign n187 = ~n184 & n186;
  assign n188 = ~n183 & n187;
  assign n189 = inD1 & n127;
  assign n190 = n114 & n188;
  assign n191 = ~n189 & ~n190;
  assign n192 = sh2 & ~n181;
  assign n193 = ~sh2 & ~n191;
  assign n194 = ~n192 & ~n193;
  assign n195 = inD3 & musel2;
  assign n196 = ~inB3 & ~n195;
  assign n197 = ~inB3 & ~musel1;
  assign n198 = n117 & ~n195;
  assign n199 = ~n121 & ~n198;
  assign n200 = ~n197 & n199;
  assign n201 = ~n196 & n200;
  assign n202 = inD3 & n127;
  assign n203 = n114 & n201;
  assign n204 = ~n202 & ~n203;
  assign n205 = sh2 & ~n140;
  assign n206 = ~sh2 & ~n204;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~sh1 & n194;
  assign n209 = n194 & n207;
  assign n210 = sh1 & n207;
  assign n211 = ~n209 & ~n210;
  assign n212 = ~n208 & n211;
  assign n213 = ~sh0 & n171;
  assign n214 = sh0 & n212;
  assign n215 = ~n213 & ~n214;
  assign n216 = ~opsel2 & n110;
  assign n217 = n110 & n215;
  assign n218 = opsel2 & n215;
  assign n219 = ~n217 & ~n218;
  assign n220 = ~n216 & n219;
  assign n221 = ~n113 & ~n220;
  assign n222 = n112 & ~n113;
  assign n223 = ~n221 & ~n222;
  assign n224 = opsel0 & opsel1;
  assign n225 = ~n112 & ~n224;
  assign n226 = opsel2 & opsel3;
  assign n227 = opsel1 & ~opsel2;
  assign n228 = ~opsel1 & ~opsel3;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~opsel0 & n229;
  assign n231 = ~n226 & n230;
  assign n232 = ~inA0 & ~n92;
  assign n233 = ~inA0 & ~musel1;
  assign n234 = ~n92 & n117;
  assign n235 = ~n121 & ~n234;
  assign n236 = ~n233 & n235;
  assign n237 = ~n232 & n236;
  assign n238 = ~musel4 & n237;
  assign n239 = musel3 & n238;
  assign n240 = inC0 & musel4;
  assign n241 = ~musel3 & n240;
  assign n242 = ~musel2 & n241;
  assign n243 = ~musel1 & n242;
  assign n244 = ~n239 & ~n243;
  assign n245 = ~n231 & ~n244;
  assign n246 = n231 & n244;
  assign n247 = ~n245 & ~n246;
  assign n248 = musel2 & ~musel3;
  assign n249 = inB0 & n248;
  assign n250 = ~musel2 & musel3;
  assign n251 = inD0 & n250;
  assign n252 = ~musel1 & n249;
  assign n253 = ~musel1 & n251;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~inA0 & ~inC0;
  assign n256 = ~inA0 & ~musel2;
  assign n257 = ~inC0 & musel2;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~n255 & n258;
  assign n260 = ~musel3 & n259;
  assign n261 = musel1 & n260;
  assign n262 = n254 & ~n261;
  assign n263 = ~musel4 & ~n262;
  assign n264 = n247 & n263;
  assign n265 = ~n247 & ~n263;
  assign n266 = ~n264 & ~n265;
  assign n267 = opsel1 & ~opsel3;
  assign n268 = opsel2 & n267;
  assign n269 = ~opsel1 & ~opsel2;
  assign n270 = opsel3 & n269;
  assign n271 = ~n268 & ~n270;
  assign n272 = ~opsel0 & ~n271;
  assign n273 = n266 & n272;
  assign n274 = n266 & ~n273;
  assign n275 = n272 & ~n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = n225 & n276;
  assign n278 = n112 & ~n215;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~opsel2 & ~n279;
  assign n281 = opsel3 & n280;
  assign n282 = ~opsel3 & n223;
  assign O0 = n281 | n282;
  assign n284 = n104 & ~n107;
  assign n285 = inC1 & musel2;
  assign n286 = inA1 & n93;
  assign n287 = ~musel1 & n285;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~musel3 & ~n288;
  assign n290 = musel4 & n289;
  assign n291 = n104 & ~n290;
  assign n292 = ~n104 & n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = ~n284 & ~n293;
  assign n295 = n284 & n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = opsel2 & ~n296;
  assign n298 = n112 & n297;
  assign n299 = inD9 & musel2;
  assign n300 = ~inB9 & ~n299;
  assign n301 = ~inB9 & ~musel1;
  assign n302 = n117 & ~n299;
  assign n303 = ~n121 & ~n302;
  assign n304 = ~n301 & n303;
  assign n305 = ~n300 & n304;
  assign n306 = inD9 & n127;
  assign n307 = n114 & n305;
  assign n308 = ~n306 & ~n307;
  assign n309 = sh2 & ~n308;
  assign n310 = ~n206 & ~n309;
  assign n311 = n194 & n310;
  assign n312 = sh1 & n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = ~n208 & n313;
  assign n315 = inD6 & musel2;
  assign n316 = ~inB6 & ~n315;
  assign n317 = ~inB6 & ~musel1;
  assign n318 = n117 & ~n315;
  assign n319 = ~n121 & ~n318;
  assign n320 = ~n317 & n319;
  assign n321 = ~n316 & n320;
  assign n322 = inD6 & n127;
  assign n323 = n114 & n321;
  assign n324 = ~n322 & ~n323;
  assign n325 = sh2 & ~n324;
  assign n326 = ~n165 & ~n325;
  assign n327 = sh2 & ~n191;
  assign n328 = ~sh2 & ~n130;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~sh1 & n326;
  assign n331 = n326 & n329;
  assign n332 = sh1 & n329;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n330 & n333;
  assign n335 = ~sh0 & n314;
  assign n336 = sh0 & n334;
  assign n337 = ~n335 & ~n336;
  assign n338 = ~opsel2 & n296;
  assign n339 = n296 & n337;
  assign n340 = opsel2 & n337;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~n338 & n341;
  assign n343 = ~n298 & ~n342;
  assign n344 = n112 & ~n298;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~inA1 & ~n285;
  assign n347 = ~inA1 & ~musel1;
  assign n348 = n117 & ~n285;
  assign n349 = ~n121 & ~n348;
  assign n350 = ~n347 & n349;
  assign n351 = ~n346 & n350;
  assign n352 = ~musel4 & n351;
  assign n353 = musel3 & n352;
  assign n354 = inC1 & musel4;
  assign n355 = ~musel3 & n354;
  assign n356 = ~musel2 & n355;
  assign n357 = ~musel1 & n356;
  assign n358 = ~n353 & ~n357;
  assign n359 = ~n231 & ~n358;
  assign n360 = n231 & n358;
  assign n361 = ~n359 & ~n360;
  assign n362 = inB1 & n248;
  assign n363 = inD1 & n250;
  assign n364 = ~musel1 & n362;
  assign n365 = ~musel1 & n363;
  assign n366 = ~n364 & ~n365;
  assign n367 = ~inA1 & ~inC1;
  assign n368 = ~inA1 & ~musel2;
  assign n369 = ~inC1 & musel2;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~n367 & n370;
  assign n372 = ~musel3 & n371;
  assign n373 = musel1 & n372;
  assign n374 = n366 & ~n373;
  assign n375 = ~musel4 & ~n374;
  assign n376 = ~n361 & ~n375;
  assign n377 = n361 & n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = n247 & ~n263;
  assign n380 = n272 & ~n379;
  assign n381 = ~n247 & n263;
  assign n382 = n378 & n380;
  assign n383 = n378 & n381;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n272 & ~n381;
  assign n386 = ~n379 & ~n385;
  assign n387 = n378 & n384;
  assign n388 = n384 & n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = n225 & n389;
  assign n391 = n112 & ~n337;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~opsel2 & ~n392;
  assign n394 = opsel3 & n393;
  assign n395 = ~opsel3 & n345;
  assign O1 = n394 | n395;
  assign n397 = n104 & ~n293;
  assign n398 = ~n107 & n397;
  assign n399 = inC2 & musel2;
  assign n400 = inA2 & n93;
  assign n401 = ~musel1 & n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~musel3 & ~n402;
  assign n404 = musel4 & n403;
  assign n405 = n104 & ~n404;
  assign n406 = ~n104 & n404;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n398 & ~n407;
  assign n409 = n398 & n407;
  assign n410 = ~n408 & ~n409;
  assign n411 = opsel2 & ~n410;
  assign n412 = n112 & n411;
  assign n413 = inD10 & musel2;
  assign n414 = ~inB10 & ~n413;
  assign n415 = ~inB10 & ~musel1;
  assign n416 = n117 & ~n413;
  assign n417 = ~n121 & ~n416;
  assign n418 = ~n415 & n417;
  assign n419 = ~n414 & n418;
  assign n420 = inD10 & n127;
  assign n421 = n114 & n419;
  assign n422 = ~n420 & ~n421;
  assign n423 = sh2 & ~n422;
  assign n424 = ~n328 & ~n423;
  assign n425 = n326 & n424;
  assign n426 = sh1 & n424;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n330 & n427;
  assign n429 = inD7 & musel2;
  assign n430 = ~inB7 & ~n429;
  assign n431 = ~inB7 & ~musel1;
  assign n432 = n117 & ~n429;
  assign n433 = ~n121 & ~n432;
  assign n434 = ~n431 & n433;
  assign n435 = ~n430 & n434;
  assign n436 = inD7 & n127;
  assign n437 = n114 & n435;
  assign n438 = ~n436 & ~n437;
  assign n439 = sh2 & ~n438;
  assign n440 = ~n206 & ~n439;
  assign n441 = sh2 & ~n163;
  assign n442 = ~sh2 & ~n181;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~sh1 & n440;
  assign n445 = n440 & n443;
  assign n446 = sh1 & n443;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n444 & n447;
  assign n449 = ~sh0 & n428;
  assign n450 = sh0 & n448;
  assign n451 = ~n449 & ~n450;
  assign n452 = ~opsel2 & n410;
  assign n453 = n410 & n451;
  assign n454 = opsel2 & n451;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~n452 & n455;
  assign n457 = ~n412 & ~n456;
  assign n458 = n112 & ~n412;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~inA2 & ~n399;
  assign n461 = ~inA2 & ~musel1;
  assign n462 = n117 & ~n399;
  assign n463 = ~n121 & ~n462;
  assign n464 = ~n461 & n463;
  assign n465 = ~n460 & n464;
  assign n466 = ~musel4 & n465;
  assign n467 = musel3 & n466;
  assign n468 = inC2 & musel4;
  assign n469 = ~musel3 & n468;
  assign n470 = ~musel2 & n469;
  assign n471 = ~musel1 & n470;
  assign n472 = ~n467 & ~n471;
  assign n473 = ~n231 & ~n472;
  assign n474 = n231 & n472;
  assign n475 = ~n473 & ~n474;
  assign n476 = inB2 & n248;
  assign n477 = inD2 & n250;
  assign n478 = ~musel1 & n476;
  assign n479 = ~musel1 & n477;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~inA2 & ~inC2;
  assign n482 = ~inA2 & ~musel2;
  assign n483 = ~inC2 & musel2;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n481 & n484;
  assign n486 = ~musel3 & n485;
  assign n487 = musel1 & n486;
  assign n488 = n480 & ~n487;
  assign n489 = ~musel4 & ~n488;
  assign n490 = ~n475 & ~n489;
  assign n491 = n475 & n489;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n380 & ~n381;
  assign n494 = n361 & ~n375;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n361 & n375;
  assign n497 = n492 & n495;
  assign n498 = n492 & n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n379 & n381;
  assign n501 = ~n380 & ~n500;
  assign n502 = ~n496 & n501;
  assign n503 = ~n494 & ~n502;
  assign n504 = n492 & n499;
  assign n505 = n499 & n503;
  assign n506 = ~n504 & ~n505;
  assign n507 = n225 & n506;
  assign n508 = n112 & ~n451;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~opsel2 & ~n509;
  assign n511 = opsel3 & n510;
  assign n512 = ~opsel3 & n459;
  assign O2 = n511 | n512;
  assign n514 = ~n293 & ~n407;
  assign n515 = ~n107 & n514;
  assign n516 = n104 & n515;
  assign n517 = inC3 & musel2;
  assign n518 = inA3 & n93;
  assign n519 = ~musel1 & n517;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~musel3 & ~n520;
  assign n522 = musel4 & n521;
  assign n523 = n104 & ~n522;
  assign n524 = ~n104 & n522;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n516 & ~n525;
  assign n527 = n516 & n525;
  assign n528 = ~n526 & ~n527;
  assign n529 = opsel2 & ~n528;
  assign n530 = n112 & n529;
  assign n531 = inD11 & musel2;
  assign n532 = ~inB11 & ~n531;
  assign n533 = ~inB11 & ~musel1;
  assign n534 = n117 & ~n531;
  assign n535 = ~n121 & ~n534;
  assign n536 = ~n533 & n535;
  assign n537 = ~n532 & n536;
  assign n538 = inD11 & n127;
  assign n539 = n114 & n537;
  assign n540 = ~n538 & ~n539;
  assign n541 = sh2 & ~n540;
  assign n542 = ~n442 & ~n541;
  assign n543 = n440 & n542;
  assign n544 = sh1 & n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n444 & n545;
  assign n547 = ~n164 & ~n328;
  assign n548 = sh2 & ~n204;
  assign n549 = ~sh2 & ~n324;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~sh1 & n547;
  assign n552 = n547 & n550;
  assign n553 = sh1 & n550;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~n551 & n554;
  assign n556 = ~sh0 & n546;
  assign n557 = sh0 & n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~opsel2 & n528;
  assign n560 = n528 & n558;
  assign n561 = opsel2 & n558;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n559 & n562;
  assign n564 = ~n530 & ~n563;
  assign n565 = n112 & ~n530;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~inA3 & ~n517;
  assign n568 = ~inA3 & ~musel1;
  assign n569 = n117 & ~n517;
  assign n570 = ~n121 & ~n569;
  assign n571 = ~n568 & n570;
  assign n572 = ~n567 & n571;
  assign n573 = ~musel4 & n572;
  assign n574 = musel3 & n573;
  assign n575 = inC3 & musel4;
  assign n576 = ~musel3 & n575;
  assign n577 = ~musel2 & n576;
  assign n578 = ~musel1 & n577;
  assign n579 = ~n574 & ~n578;
  assign n580 = ~n231 & ~n579;
  assign n581 = n231 & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = inB3 & n248;
  assign n584 = inD3 & n250;
  assign n585 = ~musel1 & n583;
  assign n586 = ~musel1 & n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~inA3 & ~inC3;
  assign n589 = ~inA3 & ~musel2;
  assign n590 = ~inC3 & musel2;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n588 & n591;
  assign n593 = ~musel3 & n592;
  assign n594 = musel1 & n593;
  assign n595 = n587 & ~n594;
  assign n596 = ~musel4 & ~n595;
  assign n597 = ~n582 & ~n596;
  assign n598 = n582 & n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n495 & ~n496;
  assign n601 = n475 & ~n489;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n475 & n489;
  assign n604 = n599 & n602;
  assign n605 = n599 & n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n503 & ~n603;
  assign n608 = ~n601 & ~n607;
  assign n609 = n606 & n608;
  assign n610 = n599 & n606;
  assign n611 = ~n609 & ~n610;
  assign n612 = n225 & n611;
  assign n613 = n112 & ~n558;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~opsel2 & ~n614;
  assign n616 = opsel3 & n615;
  assign n617 = ~opsel3 & n566;
  assign O3 = n616 | n617;
  assign n619 = ~n407 & ~n525;
  assign n620 = ~n293 & n619;
  assign n621 = ~n107 & n620;
  assign n622 = n104 & n621;
  assign n623 = inC4 & musel2;
  assign n624 = inA4 & n93;
  assign n625 = ~musel1 & n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = ~musel3 & ~n626;
  assign n628 = musel4 & n627;
  assign n629 = n104 & ~n628;
  assign n630 = ~n104 & n628;
  assign n631 = ~n629 & ~n630;
  assign n632 = n622 & n631;
  assign n633 = ~n622 & ~n631;
  assign n634 = ~n632 & ~n633;
  assign n635 = opsel2 & ~n634;
  assign n636 = n112 & n635;
  assign n637 = inD12 & musel2;
  assign n638 = ~inB12 & ~n637;
  assign n639 = ~inB12 & ~musel1;
  assign n640 = n117 & ~n637;
  assign n641 = ~n121 & ~n640;
  assign n642 = ~n639 & n641;
  assign n643 = ~n638 & n642;
  assign n644 = inD12 & n127;
  assign n645 = n114 & n643;
  assign n646 = ~n644 & ~n645;
  assign n647 = sh2 & ~n646;
  assign n648 = ~n549 & ~n647;
  assign n649 = n547 & n648;
  assign n650 = sh1 & n648;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n551 & n651;
  assign n653 = ~n309 & ~n442;
  assign n654 = ~sh2 & ~n438;
  assign n655 = ~n141 & ~n654;
  assign n656 = ~sh1 & n653;
  assign n657 = n653 & n655;
  assign n658 = sh1 & n655;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n656 & n659;
  assign n661 = ~sh0 & n652;
  assign n662 = sh0 & n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~opsel2 & n634;
  assign n665 = n634 & n663;
  assign n666 = opsel2 & n663;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n664 & n667;
  assign n669 = ~n636 & ~n668;
  assign n670 = n112 & ~n636;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~opsel2 & opsel3;
  assign n673 = opsel0 & ~opsel1;
  assign n674 = ~opsel0 & opsel1;
  assign n675 = ~n673 & ~n674;
  assign n676 = ~n247 & ~n361;
  assign n677 = ~n247 & n375;
  assign n678 = n263 & ~n361;
  assign n679 = n263 & n375;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~n677 & n680;
  assign n682 = ~n676 & n681;
  assign n683 = ~n475 & ~n582;
  assign n684 = ~n475 & n596;
  assign n685 = n489 & ~n582;
  assign n686 = n489 & n596;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n684 & n687;
  assign n689 = ~n683 & n688;
  assign n690 = ~n682 & ~n689;
  assign n691 = ~n381 & ~n496;
  assign n692 = n494 & ~n496;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~n475 & n693;
  assign n695 = n489 & n693;
  assign n696 = ~n694 & ~n695;
  assign n697 = n582 & ~n596;
  assign n698 = ~n603 & n696;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n582 & n596;
  assign n701 = ~n699 & ~n700;
  assign n702 = n272 & n690;
  assign n703 = n701 & ~n702;
  assign n704 = ~inA4 & ~n623;
  assign n705 = ~inA4 & ~musel1;
  assign n706 = n117 & ~n623;
  assign n707 = ~n121 & ~n706;
  assign n708 = ~n705 & n707;
  assign n709 = ~n704 & n708;
  assign n710 = ~musel4 & n709;
  assign n711 = musel3 & n710;
  assign n712 = inC4 & musel4;
  assign n713 = ~musel3 & n712;
  assign n714 = ~musel2 & n713;
  assign n715 = ~musel1 & n714;
  assign n716 = ~n711 & ~n715;
  assign n717 = ~n231 & ~n716;
  assign n718 = n231 & n716;
  assign n719 = ~n717 & ~n718;
  assign n720 = inB4 & n248;
  assign n721 = inD4 & n250;
  assign n722 = ~musel1 & n720;
  assign n723 = ~musel1 & n721;
  assign n724 = ~n722 & ~n723;
  assign n725 = ~inA4 & ~inC4;
  assign n726 = ~inA4 & ~musel2;
  assign n727 = ~inC4 & musel2;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n725 & n728;
  assign n730 = ~musel3 & n729;
  assign n731 = musel1 & n730;
  assign n732 = n724 & ~n731;
  assign n733 = ~musel4 & ~n732;
  assign n734 = n719 & n733;
  assign n735 = ~n719 & ~n733;
  assign n736 = ~n734 & ~n735;
  assign n737 = n703 & ~n736;
  assign n738 = ~n703 & n736;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n112 & n675;
  assign n741 = n663 & n675;
  assign n742 = ~n112 & n739;
  assign n743 = n663 & n739;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n741 & n744;
  assign n746 = ~n740 & n745;
  assign n747 = ~opsel3 & n671;
  assign n748 = n672 & n746;
  assign O4 = n747 | n748;
  assign n750 = n622 & ~n631;
  assign n751 = inC5 & musel2;
  assign n752 = inA5 & n93;
  assign n753 = ~musel1 & n751;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~musel3 & ~n754;
  assign n756 = musel4 & n755;
  assign n757 = n104 & ~n756;
  assign n758 = ~n104 & n756;
  assign n759 = ~n757 & ~n758;
  assign n760 = ~n750 & ~n759;
  assign n761 = n750 & n759;
  assign n762 = ~n760 & ~n761;
  assign n763 = opsel2 & ~n762;
  assign n764 = n112 & n763;
  assign n765 = inD13 & musel2;
  assign n766 = ~inB13 & ~n765;
  assign n767 = ~inB13 & ~musel1;
  assign n768 = n117 & ~n765;
  assign n769 = ~n121 & ~n768;
  assign n770 = ~n767 & n769;
  assign n771 = ~n766 & n770;
  assign n772 = inD13 & n127;
  assign n773 = n114 & n771;
  assign n774 = ~n772 & ~n773;
  assign n775 = sh2 & ~n774;
  assign n776 = ~n654 & ~n775;
  assign n777 = n653 & n776;
  assign n778 = sh1 & n776;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~n656 & n779;
  assign n781 = ~n423 & ~n549;
  assign n782 = ~sh2 & ~n153;
  assign n783 = ~n192 & ~n782;
  assign n784 = ~sh1 & n781;
  assign n785 = n781 & n783;
  assign n786 = sh1 & n783;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~n784 & n787;
  assign n789 = ~sh0 & n780;
  assign n790 = sh0 & n788;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~opsel2 & n762;
  assign n793 = n762 & n791;
  assign n794 = opsel2 & n791;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n792 & n795;
  assign n797 = ~n764 & ~n796;
  assign n798 = n112 & ~n764;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~inA5 & ~n751;
  assign n801 = ~inA5 & ~musel1;
  assign n802 = n117 & ~n751;
  assign n803 = ~n121 & ~n802;
  assign n804 = ~n801 & n803;
  assign n805 = ~n800 & n804;
  assign n806 = ~musel4 & n805;
  assign n807 = musel3 & n806;
  assign n808 = inC5 & musel4;
  assign n809 = ~musel3 & n808;
  assign n810 = ~musel2 & n809;
  assign n811 = ~musel1 & n810;
  assign n812 = ~n807 & ~n811;
  assign n813 = ~n231 & ~n812;
  assign n814 = n231 & n812;
  assign n815 = ~n813 & ~n814;
  assign n816 = inB5 & n248;
  assign n817 = inD5 & n250;
  assign n818 = ~musel1 & n816;
  assign n819 = ~musel1 & n817;
  assign n820 = ~n818 & ~n819;
  assign n821 = ~inA5 & ~inC5;
  assign n822 = ~inA5 & ~musel2;
  assign n823 = ~inC5 & musel2;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n821 & n824;
  assign n826 = ~musel3 & n825;
  assign n827 = musel1 & n826;
  assign n828 = n820 & ~n827;
  assign n829 = ~musel4 & ~n828;
  assign n830 = ~n815 & ~n829;
  assign n831 = n815 & n829;
  assign n832 = ~n830 & ~n831;
  assign n833 = n719 & ~n733;
  assign n834 = ~n703 & ~n833;
  assign n835 = ~n719 & n733;
  assign n836 = n832 & n834;
  assign n837 = n832 & n835;
  assign n838 = ~n836 & ~n837;
  assign n839 = n703 & ~n835;
  assign n840 = ~n833 & ~n839;
  assign n841 = n832 & n838;
  assign n842 = n838 & n840;
  assign n843 = ~n841 & ~n842;
  assign n844 = n225 & n843;
  assign n845 = n112 & ~n791;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~opsel2 & ~n846;
  assign n848 = opsel3 & n847;
  assign n849 = ~opsel3 & n799;
  assign O5 = n848 | n849;
  assign n851 = n622 & ~n759;
  assign n852 = ~n631 & n851;
  assign n853 = inC6 & musel2;
  assign n854 = inA6 & n93;
  assign n855 = ~musel1 & n853;
  assign n856 = ~n854 & ~n855;
  assign n857 = ~musel3 & ~n856;
  assign n858 = musel4 & n857;
  assign n859 = n104 & ~n858;
  assign n860 = ~n104 & n858;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n852 & ~n861;
  assign n863 = n852 & n861;
  assign n864 = ~n862 & ~n863;
  assign n865 = opsel2 & ~n864;
  assign n866 = n112 & n865;
  assign n867 = inD14 & musel2;
  assign n868 = ~inB14 & ~n867;
  assign n869 = ~inB14 & ~musel1;
  assign n870 = n117 & ~n867;
  assign n871 = ~n121 & ~n870;
  assign n872 = ~n869 & n871;
  assign n873 = ~n868 & n872;
  assign n874 = inD14 & n127;
  assign n875 = n114 & n873;
  assign n876 = ~n874 & ~n875;
  assign n877 = sh2 & ~n876;
  assign n878 = ~n782 & ~n877;
  assign n879 = n781 & n878;
  assign n880 = sh1 & n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n784 & n881;
  assign n883 = ~n541 & ~n654;
  assign n884 = ~sh2 & ~n308;
  assign n885 = ~n325 & ~n884;
  assign n886 = ~sh1 & n883;
  assign n887 = n883 & n885;
  assign n888 = sh1 & n885;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n886 & n889;
  assign n891 = ~sh0 & n882;
  assign n892 = sh0 & n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~opsel2 & n864;
  assign n895 = n864 & n893;
  assign n896 = opsel2 & n893;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n894 & n897;
  assign n899 = ~n866 & ~n898;
  assign n900 = n112 & ~n866;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~inA6 & ~n853;
  assign n903 = ~inA6 & ~musel1;
  assign n904 = n117 & ~n853;
  assign n905 = ~n121 & ~n904;
  assign n906 = ~n903 & n905;
  assign n907 = ~n902 & n906;
  assign n908 = ~musel4 & n907;
  assign n909 = musel3 & n908;
  assign n910 = inC6 & musel4;
  assign n911 = ~musel3 & n910;
  assign n912 = ~musel2 & n911;
  assign n913 = ~musel1 & n912;
  assign n914 = ~n909 & ~n913;
  assign n915 = ~n231 & ~n914;
  assign n916 = n231 & n914;
  assign n917 = ~n915 & ~n916;
  assign n918 = inB6 & n248;
  assign n919 = inD6 & n250;
  assign n920 = ~musel1 & n918;
  assign n921 = ~musel1 & n919;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~inA6 & ~inC6;
  assign n924 = ~inA6 & ~musel2;
  assign n925 = ~inC6 & musel2;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n923 & n926;
  assign n928 = ~musel3 & n927;
  assign n929 = musel1 & n928;
  assign n930 = n922 & ~n929;
  assign n931 = ~musel4 & ~n930;
  assign n932 = ~n917 & ~n931;
  assign n933 = n917 & n931;
  assign n934 = ~n932 & ~n933;
  assign n935 = ~n834 & ~n835;
  assign n936 = n815 & ~n829;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n815 & n829;
  assign n939 = n934 & n937;
  assign n940 = n934 & n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n840 & ~n938;
  assign n943 = ~n936 & ~n942;
  assign n944 = n934 & n941;
  assign n945 = n941 & n943;
  assign n946 = ~n944 & ~n945;
  assign n947 = n225 & n946;
  assign n948 = n112 & ~n893;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~opsel2 & ~n949;
  assign n951 = opsel3 & n950;
  assign n952 = ~opsel3 & n901;
  assign O6 = n951 | n952;
  assign n954 = ~n759 & ~n861;
  assign n955 = ~n631 & n954;
  assign n956 = n622 & n955;
  assign n957 = inC7 & musel2;
  assign n958 = inA7 & n93;
  assign n959 = ~musel1 & n957;
  assign n960 = ~n958 & ~n959;
  assign n961 = ~musel3 & ~n960;
  assign n962 = musel4 & n961;
  assign n963 = n104 & ~n962;
  assign n964 = ~n104 & n962;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n956 & ~n965;
  assign n967 = n956 & n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = opsel2 & ~n968;
  assign n970 = n112 & n969;
  assign n971 = inD15 & musel2;
  assign n972 = ~inB15 & ~n971;
  assign n973 = ~inB15 & ~musel1;
  assign n974 = n117 & ~n971;
  assign n975 = ~n121 & ~n974;
  assign n976 = ~n973 & n975;
  assign n977 = ~n972 & n976;
  assign n978 = inD15 & n126;
  assign n979 = musel4 & n978;
  assign n980 = n114 & n977;
  assign n981 = ~n979 & ~n980;
  assign n982 = sh2 & ~n981;
  assign n983 = ~n884 & ~n982;
  assign n984 = n883 & n983;
  assign n985 = sh1 & n983;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n886 & n986;
  assign n988 = ~n647 & ~n782;
  assign n989 = ~sh2 & ~n422;
  assign n990 = ~n439 & ~n989;
  assign n991 = ~sh1 & n988;
  assign n992 = n988 & n990;
  assign n993 = sh1 & n990;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~n991 & n994;
  assign n996 = ~sh0 & n987;
  assign n997 = sh0 & n995;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~opsel2 & n968;
  assign n1000 = n968 & n998;
  assign n1001 = opsel2 & n998;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~n999 & n1002;
  assign n1004 = ~n970 & ~n1003;
  assign n1005 = n112 & ~n970;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~inA7 & ~n957;
  assign n1008 = ~inA7 & ~musel1;
  assign n1009 = n117 & ~n957;
  assign n1010 = ~n121 & ~n1009;
  assign n1011 = ~n1008 & n1010;
  assign n1012 = ~n1007 & n1011;
  assign n1013 = ~musel4 & n1012;
  assign n1014 = musel3 & n1013;
  assign n1015 = inC7 & musel4;
  assign n1016 = ~musel3 & n1015;
  assign n1017 = ~musel2 & n1016;
  assign n1018 = ~musel1 & n1017;
  assign n1019 = ~n1014 & ~n1018;
  assign n1020 = ~n231 & ~n1019;
  assign n1021 = n231 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = inB7 & n248;
  assign n1024 = inD7 & n250;
  assign n1025 = ~musel1 & n1023;
  assign n1026 = ~musel1 & n1024;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~inA7 & ~inC7;
  assign n1029 = ~inA7 & ~musel2;
  assign n1030 = ~inC7 & musel2;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = ~n1028 & n1031;
  assign n1033 = ~musel3 & n1032;
  assign n1034 = musel1 & n1033;
  assign n1035 = n1027 & ~n1034;
  assign n1036 = ~musel4 & ~n1035;
  assign n1037 = ~n1022 & ~n1036;
  assign n1038 = n1022 & n1036;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = n833 & ~n835;
  assign n1041 = ~n839 & ~n1040;
  assign n1042 = ~n936 & n1041;
  assign n1043 = ~n938 & ~n1042;
  assign n1044 = n917 & ~n931;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~n917 & n931;
  assign n1047 = n1039 & n1045;
  assign n1048 = n1039 & n1046;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = n840 & ~n936;
  assign n1051 = ~n936 & n938;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = ~n1046 & n1052;
  assign n1054 = ~n1044 & ~n1053;
  assign n1055 = n1049 & n1054;
  assign n1056 = n1039 & n1049;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = n225 & n1057;
  assign n1059 = n112 & ~n998;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = ~opsel2 & ~n1060;
  assign n1062 = opsel3 & n1061;
  assign n1063 = ~opsel3 & n1006;
  assign O7 = n1062 | n1063;
  assign n1065 = inC8 & musel2;
  assign n1066 = inA8 & n93;
  assign n1067 = ~musel1 & n1065;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~musel3 & ~n1068;
  assign n1070 = musel4 & n1069;
  assign n1071 = n104 & ~n1070;
  assign n1072 = ~n104 & n1070;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = inC9 & musel2;
  assign n1075 = inA9 & n93;
  assign n1076 = ~musel1 & n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~musel3 & ~n1077;
  assign n1079 = musel4 & n1078;
  assign n1080 = n104 & ~n1079;
  assign n1081 = ~n104 & n1079;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = inC10 & musel2;
  assign n1084 = inA10 & n93;
  assign n1085 = ~musel1 & n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~musel3 & ~n1086;
  assign n1088 = musel4 & n1087;
  assign n1089 = n104 & ~n1088;
  assign n1090 = ~n104 & n1088;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = inC11 & musel2;
  assign n1093 = inA11 & n93;
  assign n1094 = ~musel1 & n1092;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~musel3 & ~n1095;
  assign n1097 = musel4 & n1096;
  assign n1098 = n104 & ~n1097;
  assign n1099 = ~n104 & n1097;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n1091 & ~n1100;
  assign n1102 = ~n1082 & n1101;
  assign n1103 = ~n1073 & n1102;
  assign n1104 = n621 & n1103;
  assign n1105 = n104 & n1104;
  assign n1106 = n1073 & n1105;
  assign n1107 = ~n1073 & ~n1105;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = opsel2 & ~n1108;
  assign n1110 = n112 & n1109;
  assign n1111 = ~n982 & ~n989;
  assign n1112 = n988 & n1111;
  assign n1113 = sh1 & n1111;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = ~n991 & n1114;
  assign n1116 = ~n775 & ~n884;
  assign n1117 = ~sh2 & ~n540;
  assign n1118 = ~n164 & ~n1117;
  assign n1119 = ~sh1 & n1116;
  assign n1120 = n1116 & n1118;
  assign n1121 = sh1 & n1118;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~n1119 & n1122;
  assign n1124 = ~sh0 & n1115;
  assign n1125 = sh0 & n1123;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~opsel2 & n1108;
  assign n1128 = n1108 & n1126;
  assign n1129 = opsel2 & n1126;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1127 & n1130;
  assign n1132 = ~n1110 & ~n1131;
  assign n1133 = n112 & ~n1110;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n719 & ~n815;
  assign n1136 = ~n719 & n829;
  assign n1137 = n733 & ~n815;
  assign n1138 = n733 & n829;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1136 & n1139;
  assign n1141 = ~n1135 & n1140;
  assign n1142 = ~n917 & ~n1022;
  assign n1143 = ~n917 & n1036;
  assign n1144 = n931 & ~n1022;
  assign n1145 = n931 & n1036;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1143 & n1146;
  assign n1148 = ~n1142 & n1147;
  assign n1149 = ~n1141 & ~n1148;
  assign n1150 = ~n835 & ~n938;
  assign n1151 = n936 & ~n938;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n917 & n1152;
  assign n1154 = n931 & n1152;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = n1022 & ~n1036;
  assign n1157 = ~n1046 & n1155;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = ~n1022 & n1036;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n703 & n1149;
  assign n1162 = n1160 & ~n1161;
  assign n1163 = ~inA8 & ~n1065;
  assign n1164 = ~inA8 & ~musel1;
  assign n1165 = n117 & ~n1065;
  assign n1166 = ~n121 & ~n1165;
  assign n1167 = ~n1164 & n1166;
  assign n1168 = ~n1163 & n1167;
  assign n1169 = ~musel4 & n1168;
  assign n1170 = musel3 & n1169;
  assign n1171 = inC8 & musel4;
  assign n1172 = ~musel3 & n1171;
  assign n1173 = ~musel2 & n1172;
  assign n1174 = ~musel1 & n1173;
  assign n1175 = ~n1170 & ~n1174;
  assign n1176 = ~n231 & ~n1175;
  assign n1177 = n231 & n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = inB8 & n248;
  assign n1180 = inD8 & n250;
  assign n1181 = ~musel1 & n1179;
  assign n1182 = ~musel1 & n1180;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~inA8 & ~inC8;
  assign n1185 = ~inA8 & ~musel2;
  assign n1186 = ~inC8 & musel2;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = ~n1184 & n1187;
  assign n1189 = ~musel3 & n1188;
  assign n1190 = musel1 & n1189;
  assign n1191 = n1183 & ~n1190;
  assign n1192 = ~musel4 & ~n1191;
  assign n1193 = n1178 & n1192;
  assign n1194 = ~n1178 & ~n1192;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1162 & ~n1195;
  assign n1197 = ~n1162 & n1195;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = n675 & n1126;
  assign n1200 = ~n112 & n1198;
  assign n1201 = n1126 & n1198;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1199 & n1202;
  assign n1204 = ~n740 & n1203;
  assign n1205 = ~opsel3 & n1134;
  assign n1206 = n672 & n1204;
  assign O8 = n1205 | n1206;
  assign n1208 = ~n1073 & n1105;
  assign n1209 = ~n1082 & ~n1208;
  assign n1210 = n1082 & n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = opsel2 & ~n1211;
  assign n1213 = n112 & n1212;
  assign n1214 = ~n982 & ~n1117;
  assign n1215 = n1116 & n1214;
  assign n1216 = sh1 & n1214;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~n1119 & n1217;
  assign n1219 = ~n877 & ~n989;
  assign n1220 = ~sh2 & ~n646;
  assign n1221 = ~n309 & ~n1220;
  assign n1222 = ~sh1 & n1219;
  assign n1223 = n1219 & n1221;
  assign n1224 = sh1 & n1221;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = ~n1222 & n1225;
  assign n1227 = ~sh0 & n1218;
  assign n1228 = sh0 & n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~opsel2 & n1211;
  assign n1231 = n1211 & n1229;
  assign n1232 = opsel2 & n1229;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1230 & n1233;
  assign n1235 = ~n1213 & ~n1234;
  assign n1236 = n112 & ~n1213;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~inA9 & ~n1074;
  assign n1239 = ~inA9 & ~musel1;
  assign n1240 = n117 & ~n1074;
  assign n1241 = ~n121 & ~n1240;
  assign n1242 = ~n1239 & n1241;
  assign n1243 = ~n1238 & n1242;
  assign n1244 = ~musel4 & n1243;
  assign n1245 = musel3 & n1244;
  assign n1246 = inC9 & musel4;
  assign n1247 = ~musel3 & n1246;
  assign n1248 = ~musel2 & n1247;
  assign n1249 = ~musel1 & n1248;
  assign n1250 = ~n1245 & ~n1249;
  assign n1251 = ~n231 & ~n1250;
  assign n1252 = n231 & n1250;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = inB9 & n248;
  assign n1255 = inD9 & n250;
  assign n1256 = ~musel1 & n1254;
  assign n1257 = ~musel1 & n1255;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~inA9 & ~inC9;
  assign n1260 = ~inA9 & ~musel2;
  assign n1261 = ~inC9 & musel2;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~n1259 & n1262;
  assign n1264 = ~musel3 & n1263;
  assign n1265 = musel1 & n1264;
  assign n1266 = n1258 & ~n1265;
  assign n1267 = ~musel4 & ~n1266;
  assign n1268 = ~n1253 & ~n1267;
  assign n1269 = n1253 & n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = n1178 & ~n1192;
  assign n1272 = ~n1162 & ~n1271;
  assign n1273 = ~n1178 & n1192;
  assign n1274 = n1270 & n1272;
  assign n1275 = n1270 & n1273;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1162 & ~n1273;
  assign n1278 = ~n1271 & ~n1277;
  assign n1279 = n1270 & n1276;
  assign n1280 = n1276 & n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = n225 & n1281;
  assign n1283 = n112 & ~n1229;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = ~opsel2 & ~n1284;
  assign n1286 = opsel3 & n1285;
  assign n1287 = ~opsel3 & n1237;
  assign O9 = n1286 | n1287;
  assign n1289 = ~n1082 & n1105;
  assign n1290 = ~n1073 & n1289;
  assign n1291 = ~n1091 & ~n1290;
  assign n1292 = n1091 & n1290;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = opsel2 & ~n1293;
  assign n1295 = n112 & n1294;
  assign n1296 = ~n982 & ~n1220;
  assign n1297 = n1219 & n1296;
  assign n1298 = sh1 & n1296;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = ~n1222 & n1299;
  assign n1301 = ~sh2 & ~n774;
  assign n1302 = ~n423 & ~n1301;
  assign n1303 = ~sh1 & n1214;
  assign n1304 = n1214 & n1302;
  assign n1305 = sh1 & n1302;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n1303 & n1306;
  assign n1308 = ~sh0 & n1300;
  assign n1309 = sh0 & n1307;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~opsel2 & n1293;
  assign n1312 = n1293 & n1310;
  assign n1313 = opsel2 & n1310;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1311 & n1314;
  assign n1316 = ~n1295 & ~n1315;
  assign n1317 = n112 & ~n1295;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~inA10 & ~n1083;
  assign n1320 = ~inA10 & ~musel1;
  assign n1321 = n117 & ~n1083;
  assign n1322 = ~n121 & ~n1321;
  assign n1323 = ~n1320 & n1322;
  assign n1324 = ~n1319 & n1323;
  assign n1325 = ~musel4 & n1324;
  assign n1326 = musel3 & n1325;
  assign n1327 = inC10 & musel4;
  assign n1328 = ~musel3 & n1327;
  assign n1329 = ~musel2 & n1328;
  assign n1330 = ~musel1 & n1329;
  assign n1331 = ~n1326 & ~n1330;
  assign n1332 = ~n231 & ~n1331;
  assign n1333 = n231 & n1331;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = inB10 & n248;
  assign n1336 = inD10 & n250;
  assign n1337 = ~musel1 & n1335;
  assign n1338 = ~musel1 & n1336;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~inA10 & ~inC10;
  assign n1341 = ~inA10 & ~musel2;
  assign n1342 = ~inC10 & musel2;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1340 & n1343;
  assign n1345 = ~musel3 & n1344;
  assign n1346 = musel1 & n1345;
  assign n1347 = n1339 & ~n1346;
  assign n1348 = ~musel4 & ~n1347;
  assign n1349 = n1334 & n1348;
  assign n1350 = ~n1334 & ~n1348;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1272 & ~n1273;
  assign n1353 = n1253 & ~n1267;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = ~n1253 & n1267;
  assign n1356 = n1351 & n1354;
  assign n1357 = n1351 & n1355;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~n1278 & ~n1355;
  assign n1360 = ~n1353 & ~n1359;
  assign n1361 = n1351 & n1358;
  assign n1362 = n1358 & n1360;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n225 & n1363;
  assign n1365 = n112 & ~n1310;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~opsel2 & ~n1366;
  assign n1368 = opsel3 & n1367;
  assign n1369 = ~opsel3 & n1318;
  assign O10 = n1368 | n1369;
  assign n1371 = ~n1082 & ~n1091;
  assign n1372 = ~n1073 & n1371;
  assign n1373 = n1105 & n1372;
  assign n1374 = ~n1100 & ~n1373;
  assign n1375 = n1100 & n1373;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = opsel2 & ~n1376;
  assign n1378 = n112 & n1377;
  assign n1379 = sh0 & sh1;
  assign n1380 = ~sh2 & ~n876;
  assign n1381 = ~sh2 & ~n1380;
  assign n1382 = n540 & ~n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = sh1 & ~n774;
  assign n1385 = n540 & ~n1384;
  assign n1386 = sh1 & ~n1384;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = sh0 & ~sh1;
  assign n1389 = ~sh0 & n1387;
  assign n1390 = ~n646 & n1388;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n982 & n1391;
  assign n1393 = n1379 & n1391;
  assign n1394 = sh2 & ~n982;
  assign n1395 = sh2 & n1379;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1393 & n1396;
  assign n1398 = ~n1392 & n1397;
  assign n1399 = n1379 & n1383;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = ~opsel2 & n1376;
  assign n1402 = n1376 & n1400;
  assign n1403 = opsel2 & n1400;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1401 & n1404;
  assign n1406 = ~n1378 & ~n1405;
  assign n1407 = n112 & ~n1378;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~inA11 & ~n1092;
  assign n1410 = ~inA11 & ~musel1;
  assign n1411 = n117 & ~n1092;
  assign n1412 = ~n121 & ~n1411;
  assign n1413 = ~n1410 & n1412;
  assign n1414 = ~n1409 & n1413;
  assign n1415 = ~musel4 & n1414;
  assign n1416 = musel3 & n1415;
  assign n1417 = inC11 & musel4;
  assign n1418 = ~musel3 & n1417;
  assign n1419 = ~musel2 & n1418;
  assign n1420 = ~musel1 & n1419;
  assign n1421 = ~n1416 & ~n1420;
  assign n1422 = ~n231 & ~n1421;
  assign n1423 = n231 & n1421;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = inB11 & n248;
  assign n1426 = inD11 & n250;
  assign n1427 = ~musel1 & n1425;
  assign n1428 = ~musel1 & n1426;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~inA11 & ~inC11;
  assign n1431 = ~inA11 & ~musel2;
  assign n1432 = ~inC11 & musel2;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = ~musel3 & n1434;
  assign n1436 = musel1 & n1435;
  assign n1437 = n1429 & ~n1436;
  assign n1438 = ~musel4 & ~n1437;
  assign n1439 = n1424 & n1438;
  assign n1440 = ~n1424 & ~n1438;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n1271 & ~n1273;
  assign n1443 = ~n1277 & ~n1442;
  assign n1444 = ~n1353 & n1443;
  assign n1445 = ~n1355 & ~n1444;
  assign n1446 = n1334 & ~n1348;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1334 & n1348;
  assign n1449 = n1441 & n1447;
  assign n1450 = n1441 & n1448;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = n1278 & ~n1353;
  assign n1453 = ~n1353 & n1355;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1448 & n1454;
  assign n1456 = ~n1446 & ~n1455;
  assign n1457 = n1451 & n1456;
  assign n1458 = n1441 & n1451;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = n225 & n1459;
  assign n1461 = n112 & ~n1400;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~opsel2 & ~n1462;
  assign n1464 = opsel3 & n1463;
  assign n1465 = ~opsel3 & n1408;
  assign O11 = n1464 | n1465;
  assign n1467 = ~n861 & ~n965;
  assign n1468 = ~n759 & n1467;
  assign n1469 = ~n631 & n1468;
  assign n1470 = n1103 & n1469;
  assign n1471 = n104 & n1470;
  assign n1472 = n621 & n1471;
  assign n1473 = inC12 & musel2;
  assign n1474 = inA12 & n93;
  assign n1475 = ~musel1 & n1473;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~musel3 & ~n1476;
  assign n1478 = musel4 & n1477;
  assign n1479 = n104 & ~n1478;
  assign n1480 = ~n104 & n1478;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = n1472 & n1481;
  assign n1483 = ~n1472 & ~n1481;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = opsel2 & ~n1484;
  assign n1486 = n112 & n1485;
  assign n1487 = ~n981 & n1379;
  assign n1488 = ~n774 & n1388;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = sh1 & ~n876;
  assign n1491 = ~sh1 & ~n646;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n1489 & n1492;
  assign n1494 = sh0 & n1489;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = n646 & n1379;
  assign n1497 = n981 & ~n1379;
  assign n1498 = n646 & n981;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1496 & n1499;
  assign n1501 = ~sh2 & n1495;
  assign n1502 = sh2 & n1500;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~opsel2 & n1484;
  assign n1505 = n1484 & n1503;
  assign n1506 = opsel2 & n1503;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1504 & n1507;
  assign n1509 = ~n1486 & ~n1508;
  assign n1510 = n112 & ~n1486;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1253 & n1273;
  assign n1513 = n1267 & n1273;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1355 & n1514;
  assign n1516 = ~n1446 & ~n1515;
  assign n1517 = ~n1448 & ~n1516;
  assign n1518 = n1424 & ~n1438;
  assign n1519 = ~n1438 & n1517;
  assign n1520 = ~n1438 & n1518;
  assign n1521 = n1424 & n1517;
  assign n1522 = n1424 & n1518;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1520 & n1523;
  assign n1525 = ~n1519 & n1524;
  assign n1526 = ~n1178 & ~n1253;
  assign n1527 = ~n1178 & n1267;
  assign n1528 = n1192 & ~n1253;
  assign n1529 = n1192 & n1267;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1527 & n1530;
  assign n1532 = ~n1526 & n1531;
  assign n1533 = ~n1334 & ~n1424;
  assign n1534 = ~n1334 & n1438;
  assign n1535 = n1348 & ~n1424;
  assign n1536 = n1348 & n1438;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1534 & n1537;
  assign n1539 = ~n1533 & n1538;
  assign n1540 = ~n1162 & ~n1539;
  assign n1541 = ~n1532 & n1540;
  assign n1542 = ~n1525 & ~n1541;
  assign n1543 = ~inA12 & ~n1473;
  assign n1544 = ~inA12 & ~musel1;
  assign n1545 = n117 & ~n1473;
  assign n1546 = ~n121 & ~n1545;
  assign n1547 = ~n1544 & n1546;
  assign n1548 = ~n1543 & n1547;
  assign n1549 = ~musel4 & n1548;
  assign n1550 = musel3 & n1549;
  assign n1551 = inC12 & musel4;
  assign n1552 = ~musel3 & n1551;
  assign n1553 = ~musel2 & n1552;
  assign n1554 = ~musel1 & n1553;
  assign n1555 = ~n1550 & ~n1554;
  assign n1556 = ~n231 & ~n1555;
  assign n1557 = n231 & n1555;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = inB12 & n248;
  assign n1560 = inD12 & n250;
  assign n1561 = ~musel1 & n1559;
  assign n1562 = ~musel1 & n1560;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = ~inA12 & ~inC12;
  assign n1565 = ~inA12 & ~musel2;
  assign n1566 = ~inC12 & musel2;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1564 & n1567;
  assign n1569 = ~musel3 & n1568;
  assign n1570 = musel1 & n1569;
  assign n1571 = n1563 & ~n1570;
  assign n1572 = ~musel4 & ~n1571;
  assign n1573 = n1558 & n1572;
  assign n1574 = ~n1558 & ~n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = n1542 & ~n1575;
  assign n1577 = ~n1542 & n1575;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = n675 & n1503;
  assign n1580 = ~n112 & n1578;
  assign n1581 = n1503 & n1578;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~n1579 & n1582;
  assign n1584 = ~n740 & n1583;
  assign n1585 = ~opsel3 & n1511;
  assign n1586 = n672 & n1584;
  assign O12 = n1585 | n1586;
  assign n1588 = n1472 & ~n1481;
  assign n1589 = inC13 & musel2;
  assign n1590 = inA13 & n93;
  assign n1591 = ~musel1 & n1589;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~musel3 & ~n1592;
  assign n1594 = musel4 & n1593;
  assign n1595 = n104 & ~n1594;
  assign n1596 = ~n104 & n1594;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1588 & ~n1597;
  assign n1599 = n1588 & n1597;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = opsel2 & ~n1600;
  assign n1602 = n112 & n1601;
  assign n1603 = sh0 & sh2;
  assign n1604 = ~sh1 & ~sh2;
  assign n1605 = sh1 & ~n1603;
  assign n1606 = ~sh1 & sh2;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = sh0 & ~n876;
  assign n1609 = ~sh0 & ~n774;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = ~n1604 & n1607;
  assign n1612 = n981 & ~n1604;
  assign n1613 = n1607 & n1610;
  assign n1614 = n981 & n1610;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = ~n1611 & n1616;
  assign n1618 = n1384 & n1603;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~opsel2 & n1600;
  assign n1621 = n1600 & n1619;
  assign n1622 = opsel2 & n1619;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n1620 & n1623;
  assign n1625 = ~n1602 & ~n1624;
  assign n1626 = n112 & ~n1602;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~inA13 & ~n1589;
  assign n1629 = ~inA13 & ~musel1;
  assign n1630 = n117 & ~n1589;
  assign n1631 = ~n121 & ~n1630;
  assign n1632 = ~n1629 & n1631;
  assign n1633 = ~n1628 & n1632;
  assign n1634 = ~musel4 & n1633;
  assign n1635 = musel3 & n1634;
  assign n1636 = inC13 & musel4;
  assign n1637 = ~musel3 & n1636;
  assign n1638 = ~musel2 & n1637;
  assign n1639 = ~musel1 & n1638;
  assign n1640 = ~n1635 & ~n1639;
  assign n1641 = ~n231 & ~n1640;
  assign n1642 = n231 & n1640;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = inB13 & n248;
  assign n1645 = inD13 & n250;
  assign n1646 = ~musel1 & n1644;
  assign n1647 = ~musel1 & n1645;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~inA13 & ~inC13;
  assign n1650 = ~inA13 & ~musel2;
  assign n1651 = ~inC13 & musel2;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = ~n1649 & n1652;
  assign n1654 = ~musel3 & n1653;
  assign n1655 = musel1 & n1654;
  assign n1656 = n1648 & ~n1655;
  assign n1657 = ~musel4 & ~n1656;
  assign n1658 = ~n1643 & ~n1657;
  assign n1659 = n1643 & n1657;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = n1558 & ~n1572;
  assign n1662 = ~n1542 & ~n1661;
  assign n1663 = ~n1558 & n1572;
  assign n1664 = n1660 & n1662;
  assign n1665 = n1660 & n1663;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = n1542 & ~n1663;
  assign n1668 = ~n1661 & ~n1667;
  assign n1669 = n1660 & n1666;
  assign n1670 = n1666 & n1668;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = n225 & n1671;
  assign n1673 = n112 & ~n1619;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~opsel2 & ~n1674;
  assign n1676 = opsel3 & n1675;
  assign n1677 = ~opsel3 & n1627;
  assign O13 = n1676 | n1677;
  assign n1679 = n1472 & ~n1597;
  assign n1680 = ~n1481 & n1679;
  assign n1681 = inC14 & musel2;
  assign n1682 = inA14 & n93;
  assign n1683 = ~musel1 & n1681;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = ~musel3 & ~n1684;
  assign n1686 = musel4 & n1685;
  assign n1687 = ~n104 & n1686;
  assign n1688 = n104 & ~n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1680 & ~n1689;
  assign n1691 = n1680 & n1689;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = opsel2 & ~n1692;
  assign n1694 = n112 & n1693;
  assign n1695 = ~sh0 & ~sh2;
  assign n1696 = sh1 & ~sh2;
  assign n1697 = ~n1379 & ~n1696;
  assign n1698 = ~n1695 & n1697;
  assign n1699 = ~n1696 & ~n1698;
  assign n1700 = ~n981 & ~n1699;
  assign n1701 = ~n876 & n1699;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~opsel2 & n1692;
  assign n1704 = n1692 & n1702;
  assign n1705 = opsel2 & n1702;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1703 & n1706;
  assign n1708 = ~n1694 & ~n1707;
  assign n1709 = n112 & ~n1694;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~inA14 & ~n1681;
  assign n1712 = ~inA14 & ~musel1;
  assign n1713 = n117 & ~n1681;
  assign n1714 = ~n121 & ~n1713;
  assign n1715 = ~n1712 & n1714;
  assign n1716 = ~n1711 & n1715;
  assign n1717 = ~musel4 & n1716;
  assign n1718 = musel3 & n1717;
  assign n1719 = inC14 & musel4;
  assign n1720 = ~musel3 & n1719;
  assign n1721 = ~musel2 & n1720;
  assign n1722 = ~musel1 & n1721;
  assign n1723 = ~n1718 & ~n1722;
  assign n1724 = ~n231 & ~n1723;
  assign n1725 = n231 & n1723;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = inB14 & n248;
  assign n1728 = inD14 & n250;
  assign n1729 = ~musel1 & n1727;
  assign n1730 = ~musel1 & n1728;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = ~inA14 & ~inC14;
  assign n1733 = ~inA14 & ~musel2;
  assign n1734 = ~inC14 & musel2;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = ~n1732 & n1735;
  assign n1737 = ~musel3 & n1736;
  assign n1738 = musel1 & n1737;
  assign n1739 = n1731 & ~n1738;
  assign n1740 = ~musel4 & ~n1739;
  assign n1741 = ~n1726 & ~n1740;
  assign n1742 = n1726 & n1740;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = ~n1662 & ~n1663;
  assign n1745 = n1643 & ~n1657;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n1643 & n1657;
  assign n1748 = n1743 & n1746;
  assign n1749 = n1743 & n1747;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = ~n1668 & ~n1747;
  assign n1752 = ~n1745 & ~n1751;
  assign n1753 = n1743 & n1750;
  assign n1754 = n1750 & n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = n225 & n1755;
  assign n1757 = n112 & ~n1702;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~opsel2 & ~n1758;
  assign n1760 = opsel3 & n1759;
  assign n1761 = ~opsel3 & n1710;
  assign O14 = n1760 | n1761;
  assign n1763 = ~n1597 & ~n1689;
  assign n1764 = ~n1481 & n1763;
  assign n1765 = n1472 & n1764;
  assign n1766 = opsel2 & n112;
  assign n1767 = n1765 & n1766;
  assign n1768 = opsel2 & ~n981;
  assign n1769 = ~opsel2 & n1765;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1767 & n1770;
  assign n1772 = n112 & ~n1767;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~inA15 & ~n99;
  assign n1775 = ~inA15 & ~musel1;
  assign n1776 = ~n99 & n117;
  assign n1777 = ~n121 & ~n1776;
  assign n1778 = ~n1775 & n1777;
  assign n1779 = ~n1774 & n1778;
  assign n1780 = ~musel4 & n1779;
  assign n1781 = musel3 & n1780;
  assign n1782 = inC15 & musel4;
  assign n1783 = ~musel3 & n1782;
  assign n1784 = ~musel2 & n1783;
  assign n1785 = ~musel1 & n1784;
  assign n1786 = ~n1781 & ~n1785;
  assign n1787 = ~n231 & ~n1786;
  assign n1788 = n231 & n1786;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = inB15 & n248;
  assign n1791 = inD15 & n250;
  assign n1792 = ~musel1 & n1790;
  assign n1793 = ~musel1 & n1791;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = ~inA15 & ~inC15;
  assign n1796 = ~inA15 & ~musel2;
  assign n1797 = ~inC15 & musel2;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = ~n1795 & n1798;
  assign n1800 = ~musel3 & n1799;
  assign n1801 = musel1 & n1800;
  assign n1802 = n1794 & ~n1801;
  assign n1803 = ~musel4 & ~n1802;
  assign n1804 = ~n1789 & ~n1803;
  assign n1805 = n1789 & n1803;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = n1661 & ~n1663;
  assign n1808 = ~n1667 & ~n1807;
  assign n1809 = ~n1745 & n1808;
  assign n1810 = ~n1747 & ~n1809;
  assign n1811 = n1726 & ~n1740;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = ~n1726 & n1740;
  assign n1814 = n1806 & n1812;
  assign n1815 = n1806 & n1813;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = n1668 & ~n1745;
  assign n1818 = ~n1745 & n1747;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~n1813 & n1819;
  assign n1821 = ~n1811 & ~n1820;
  assign n1822 = n1816 & n1821;
  assign n1823 = n1806 & n1816;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = n225 & n1824;
  assign n1826 = n112 & ~n981;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = ~opsel2 & ~n1827;
  assign n1829 = opsel3 & n1828;
  assign n1830 = ~opsel3 & n1773;
  assign O15 = n1829 | n1830;
endmodule


