// Benchmark "pair" written by ABC on Tue May 16 16:07:51 2017

module pair ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, c0, c1, c2, c3, c4,
    c5, d0, d1, d2, d3, d4, d5, e0, e1, e2, e3, e4, e5, f0, f1, f2, f3, f4,
    f5, g0, g1, g2, g3, g4, g5, h0, h1, h2, h3, h4, h5, i0, i1, i2, i3, i4,
    i5, j0, j1, j2, j3, j4, j5, k0, k1, k2, k3, k4, k5, l0, l1, l2, l3, l4,
    l5, m0, m1, m2, m3, m4, m5, n0, n1, n2, n3, n4, n5, o0, o1, o2, o3, o4,
    o5, p0, p1, p2, p3, p4, p5, q0, q1, q2, q3, q4, q5, r0, r1, r2, r3, r4,
    r5, s0, s1, s2, s3, s4, t0, t1, t2, t3, t4, u0, u1, u2, u3, u4, v0, v1,
    v2, v3, v4, w0, w1, w2, w3, w4, x0, x1, x2, x3, x4, y0, y1, y2, y3, y4,
    z0, z1, z2, z3, z4,
    h10, x10, i10, y10, j10, k10, l10, m10, n10, a6, a7, a8, a9, b6, b7,
    b8, b9, c6, c7, c8, c9, d6, d7, d8, d9, e6, e7, e8, e9, f6, f7, f8, f9,
    g6, g7, g8, g9, h6, h7, h8, h9, i6, i7, i8, i9, j6, j7, j8, j9, k6, k7,
    k8, k9, l6, l7, l8, l9, m6, m7, m8, m9, n6, n7, n8, n9, o10, o6, o7,
    o8, o9, p6, p7, p8, p9, q6, q7, q8, q9, r6, r7, r8, r9, s5, s6, s7, s8,
    s9, t5, t6, t7, t8, t9, u5, u6, u7, u8, u9, v5, v6, v7, v8, v9, w5, w6,
    w7, w8, w9, x5, x6, x7, x8, x9, y5, y6, y7, y8, y9, z5, z6, z7, z8, z9,
    p10, a10, q10, b10, r10, c10, s10, d10, t10, e10, u10, f10, v10, g10,
    w10  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, c0, c1, c2,
    c3, c4, c5, d0, d1, d2, d3, d4, d5, e0, e1, e2, e3, e4, e5, f0, f1, f2,
    f3, f4, f5, g0, g1, g2, g3, g4, g5, h0, h1, h2, h3, h4, h5, i0, i1, i2,
    i3, i4, i5, j0, j1, j2, j3, j4, j5, k0, k1, k2, k3, k4, k5, l0, l1, l2,
    l3, l4, l5, m0, m1, m2, m3, m4, m5, n0, n1, n2, n3, n4, n5, o0, o1, o2,
    o3, o4, o5, p0, p1, p2, p3, p4, p5, q0, q1, q2, q3, q4, q5, r0, r1, r2,
    r3, r4, r5, s0, s1, s2, s3, s4, t0, t1, t2, t3, t4, u0, u1, u2, u3, u4,
    v0, v1, v2, v3, v4, w0, w1, w2, w3, w4, x0, x1, x2, x3, x4, y0, y1, y2,
    y3, y4, z0, z1, z2, z3, z4;
  output h10, x10, i10, y10, j10, k10, l10, m10, n10, a6, a7, a8, a9, b6, b7,
    b8, b9, c6, c7, c8, c9, d6, d7, d8, d9, e6, e7, e8, e9, f6, f7, f8, f9,
    g6, g7, g8, g9, h6, h7, h8, h9, i6, i7, i8, i9, j6, j7, j8, j9, k6, k7,
    k8, k9, l6, l7, l8, l9, m6, m7, m8, m9, n6, n7, n8, n9, o10, o6, o7,
    o8, o9, p6, p7, p8, p9, q6, q7, q8, q9, r6, r7, r8, r9, s5, s6, s7, s8,
    s9, t5, t6, t7, t8, t9, u5, u6, u7, u8, u9, v5, v6, v7, v8, v9, w5, w6,
    w7, w8, w9, x5, x6, x7, x8, x9, y5, y6, y7, y8, y9, z5, z6, z7, z8, z9,
    p10, a10, q10, b10, r10, c10, s10, d10, t10, e10, u10, f10, v10, g10,
    w10;
  wire n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n337, n338, n339, n340, n342, n343, n344, n345, n346, n347,
    n349, n350, n351, n352, n353, n354, n356, n357, n358, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n374, n375,
    n376, n377, n378, n379, n380, n382, n383, n384, n385, n386, n387, n388,
    n390, n391, n392, n393, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n652, n653, n654, n655, n656, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n711, n712, n713, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n727, n728,
    n729, n730, n731, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n768,
    n769, n770, n771, n772, n773, n774, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n814, n815, n816, n817, n818, n819, n820,
    n821, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n837, n838, n839, n840, n841, n842, n843, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n857, n858, n859, n860,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n920, n921, n922, n923, n924,
    n926, n927, n928, n929, n930, n931, n932, n934, n935, n936, n937, n938,
    n939, n940, n941, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n959, n960, n961, n962, n963, n964,
    n965, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1013, n1014,
    n1015, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1035, n1036, n1037,
    n1038, n1040, n1041, n1042, n1043, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1087, n1088, n1089, n1090, n1091, n1093,
    n1094, n1095, n1097, n1098, n1099, n1100, n1101, n1102, n1104, n1105,
    n1106, n1107, n1109, n1110, n1111, n1113, n1114, n1115, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1163,
    n1164, n1165, n1166, n1167, n1168, n1170, n1171, n1172, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1184, n1185, n1186,
    n1187, n1188, n1190, n1191, n1192, n1194, n1195, n1196, n1197, n1198,
    n1199, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1209, n1210,
    n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1235, n1236, n1237, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1293, n1294, n1295, n1296, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1390, n1391, n1392, n1393, n1394, n1395, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1535, n1536,
    n1537, n1538, n1540, n1541, n1542, n1544, n1545, n1546, n1548, n1549,
    n1550, n1551, n1552, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1592,
    n1593, n1594, n1595, n1597, n1598, n1599, n1600, n1601, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1642, n1643, n1644, n1645, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1680,
    n1681, n1682, n1683, n1684, n1685, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1716, n1717, n1718, n1719, n1720, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1744, n1745, n1746, n1748,
    n1749, n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1761, n1762, n1763, n1764, n1765, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1791, n1792, n1793,
    n1794, n1795, n1796, n1798, n1799, n1800, n1801, n1802, n1804, n1805,
    n1806, n1807, n1809, n1810, n1811;
  assign n311 = l5 & ~m5;
  assign n312 = n5 & n311;
  assign n313 = ~z & ~n312;
  assign n314 = n5 & n313;
  assign n315 = ~b0 & m5;
  assign n316 = ~b0 & ~n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~c0 & ~n314;
  assign n319 = ~c0 & ~l5;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~n317 & ~n320;
  assign n322 = ~z & ~q5;
  assign n323 = ~r5 & n322;
  assign n324 = ~z & ~p5;
  assign n325 = ~r5 & n324;
  assign n326 = ~q5 & n324;
  assign n327 = ~n325 & ~n326;
  assign n328 = ~n323 & n327;
  assign n329 = q5 & ~n328;
  assign n330 = n321 & n329;
  assign n331 = r5 & ~n328;
  assign n332 = n317 & n331;
  assign n333 = p5 & ~n328;
  assign n334 = n320 & n333;
  assign n335 = ~n332 & ~n334;
  assign x10 = n330 | ~n335;
  assign n337 = n321 & n331;
  assign n338 = n317 & n333;
  assign n339 = n320 & n329;
  assign n340 = ~n338 & ~n339;
  assign y10 = n337 | ~n340;
  assign n342 = g5 & ~i5;
  assign n343 = o5 & n342;
  assign n344 = a5 & ~b5;
  assign n345 = n343 & n344;
  assign n346 = ~d5 & n344;
  assign n347 = ~n345 & n346;
  assign j10 = e5 | n347;
  assign n349 = ~e5 & ~n345;
  assign n350 = n343 & n349;
  assign n351 = ~d5 & ~n350;
  assign n352 = n313 & ~n344;
  assign n353 = ~n351 & n352;
  assign n354 = ~d5 & ~n351;
  assign k10 = n353 | n354;
  assign n356 = n313 & j10;
  assign n357 = ~n343 & n356;
  assign n358 = ~e5 & j10;
  assign l10 = n357 | n358;
  assign n360 = d4 & e4;
  assign n361 = f4 & n360;
  assign n362 = ~j0 & q5;
  assign n363 = ~n361 & ~n362;
  assign n364 = i4 & ~n363;
  assign n365 = ~j0 & ~p5;
  assign n366 = ~n364 & n365;
  assign n367 = g4 & ~n366;
  assign n368 = p4 & n367;
  assign n369 = n311 & n313;
  assign n370 = ~z & n5;
  assign n371 = ~z & m5;
  assign n372 = ~n369 & ~n371;
  assign v10 = ~n370 & n372;
  assign n374 = n313 & ~n369;
  assign n375 = ~v10 & ~n374;
  assign n376 = ~z & ~h5;
  assign n377 = n368 & n376;
  assign n378 = ~z & h5;
  assign n379 = ~n368 & n378;
  assign n380 = ~n375 & ~n379;
  assign o10 = n377 | ~n380;
  assign n382 = ~h5 & o10;
  assign n383 = ~f5 & ~g5;
  assign n384 = ~n375 & n383;
  assign n385 = n382 & n384;
  assign n386 = f5 & ~n375;
  assign n387 = ~n382 & n386;
  assign n388 = ~z & ~n387;
  assign m10 = n385 | ~n388;
  assign n390 = ~z & g5;
  assign n391 = ~n382 & n390;
  assign n392 = f5 & ~m10;
  assign n393 = ~n375 & ~n392;
  assign n10 = n391 | ~n393;
  assign n395 = o0 & r5;
  assign n396 = n0 & p5;
  assign n397 = m5 & p0;
  assign n398 = t0 & w4;
  assign n399 = r4 & u0;
  assign n400 = m4 & q0;
  assign n401 = h4 & r0;
  assign n402 = d4 & s0;
  assign n403 = k0 & q3;
  assign n404 = l0 & m3;
  assign n405 = f3 & m0;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n403 & n406;
  assign n408 = ~n402 & n407;
  assign n409 = ~n401 & n408;
  assign n410 = ~n400 & n409;
  assign n411 = ~n399 & n410;
  assign n412 = ~n398 & n411;
  assign n413 = ~n397 & n412;
  assign n414 = ~n396 & n413;
  assign a6 = n395 | ~n414;
  assign n416 = ~x0 & ~y0;
  assign n417 = ~z0 & n416;
  assign n418 = ~a1 & n417;
  assign n419 = ~b1 & n418;
  assign n420 = ~c1 & n419;
  assign n421 = l1 & ~m1;
  assign n422 = n1 & n421;
  assign n423 = ~b & ~n422;
  assign n424 = n421 & n423;
  assign n425 = ~b & n1;
  assign n426 = ~b & m1;
  assign n427 = ~n424 & ~n426;
  assign v6 = ~n425 & n427;
  assign n429 = ~d1 & ~w0;
  assign n430 = v6 & n429;
  assign n431 = n420 & n430;
  assign n432 = ~n424 & ~n431;
  assign n433 = ~v0 & ~n424;
  assign n434 = ~n432 & ~n433;
  assign n435 = ~b & ~n434;
  assign n436 = ~h & ~p1;
  assign n437 = ~q1 & n436;
  assign n438 = ~n420 & n437;
  assign n439 = ~r1 & n437;
  assign n440 = ~n417 & n436;
  assign n441 = ~h & ~n416;
  assign n442 = ~h & ~v6;
  assign n443 = ~h & ~w0;
  assign n444 = ~h & v0;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n442 & n445;
  assign n447 = ~n441 & n446;
  assign n448 = ~n440 & n447;
  assign n449 = ~n439 & n448;
  assign n450 = ~n438 & n449;
  assign n451 = j1 & ~k1;
  assign n452 = o1 & n451;
  assign n453 = e1 & ~f1;
  assign n454 = n452 & n453;
  assign n455 = ~h1 & n453;
  assign n456 = ~n454 & n455;
  assign n6 = i1 | n456;
  assign n458 = ~g1 & ~n6;
  assign n459 = ~i & n458;
  assign n460 = s1 & ~n459;
  assign n461 = n450 & n460;
  assign n462 = ~s1 & n459;
  assign n463 = n450 & n462;
  assign n464 = ~n461 & ~n463;
  assign n465 = ~b & n434;
  assign n466 = t1 & n464;
  assign n467 = n435 & n466;
  assign n468 = ~t1 & ~n464;
  assign n469 = n435 & n468;
  assign n470 = x2 & n465;
  assign n471 = ~n469 & ~n470;
  assign a7 = n467 | ~n471;
  assign n473 = q2 & r2;
  assign n474 = m1 & ~n1;
  assign n475 = ~b & l1;
  assign n476 = ~b & ~n474;
  assign n477 = ~n475 & ~n476;
  assign n478 = n474 & ~n477;
  assign n479 = ~j & n478;
  assign n480 = ~p1 & ~q1;
  assign n481 = ~n473 & n480;
  assign n482 = ~n473 & ~n479;
  assign n483 = ~s2 & ~n479;
  assign n484 = ~p1 & ~s2;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~n482 & n485;
  assign n487 = ~n481 & n486;
  assign n488 = ~g & ~v6;
  assign n489 = ~g & n458;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~q2 & ~r2;
  assign n492 = ~q1 & ~n487;
  assign n493 = ~n491 & n492;
  assign n494 = ~n479 & ~n491;
  assign n495 = s2 & ~n487;
  assign n496 = ~p1 & s2;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n494 & n497;
  assign n499 = ~n493 & n498;
  assign n500 = ~i1 & ~n454;
  assign n501 = n452 & n500;
  assign n502 = ~h1 & ~n501;
  assign n503 = n458 & n502;
  assign n504 = ~v0 & ~n503;
  assign n505 = n431 & n504;
  assign n506 = ~r1 & n478;
  assign n507 = v0 & n478;
  assign n508 = ~f & ~n507;
  assign n509 = ~n506 & n508;
  assign n510 = ~n505 & n509;
  assign n511 = ~n487 & n490;
  assign n512 = ~n490 & ~n499;
  assign n513 = ~n510 & ~n512;
  assign n514 = ~n511 & n513;
  assign n515 = n477 & n490;
  assign n516 = ~t2 & ~n477;
  assign n517 = n514 & n516;
  assign n518 = t2 & ~n477;
  assign n519 = ~n514 & n518;
  assign n520 = ~n515 & ~n519;
  assign a8 = n517 | ~n520;
  assign n522 = f3 & g3;
  assign n523 = m5 & ~n5;
  assign n524 = ~z & l5;
  assign n525 = ~z & ~n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = n523 & ~n526;
  assign n528 = ~h0 & n527;
  assign n529 = ~p5 & ~q5;
  assign n530 = ~n522 & n529;
  assign n531 = ~n522 & ~n528;
  assign n532 = ~h3 & ~n528;
  assign n533 = ~h3 & ~p5;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n531 & n534;
  assign n536 = ~n530 & n535;
  assign n537 = ~c5 & ~j10;
  assign n538 = ~e0 & ~v10;
  assign n539 = ~e0 & n537;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~f3 & ~g3;
  assign n542 = ~q5 & ~n536;
  assign n543 = ~n541 & n542;
  assign n544 = ~n528 & ~n541;
  assign n545 = h3 & ~n536;
  assign n546 = ~p5 & n536;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n544 & n547;
  assign n549 = ~n543 & n548;
  assign n550 = ~t4 & ~u4;
  assign n551 = ~v4 & n550;
  assign n552 = ~w4 & n551;
  assign n553 = ~x4 & n552;
  assign n554 = ~y4 & n553;
  assign n555 = ~s4 & ~z4;
  assign n556 = n554 & n555;
  assign n557 = ~r4 & v10;
  assign n558 = n351 & n537;
  assign n559 = n557 & ~n558;
  assign n560 = n556 & n559;
  assign n561 = ~j5 & k5;
  assign n562 = ~r5 & n561;
  assign n563 = ~j5 & r4;
  assign n564 = k5 & n563;
  assign n565 = ~d0 & ~n564;
  assign n566 = ~n562 & n565;
  assign n567 = ~n560 & n566;
  assign n568 = ~n536 & n540;
  assign n569 = ~n540 & ~n549;
  assign n570 = ~n567 & ~n569;
  assign n571 = ~n568 & n570;
  assign n572 = i3 & n540;
  assign n573 = n571 & n572;
  assign n574 = h0 & ~n567;
  assign n575 = ~i3 & ~n540;
  assign n576 = n571 & n575;
  assign n577 = ~n574 & ~n576;
  assign n578 = ~n573 & n577;
  assign n579 = n540 & ~n578;
  assign n580 = ~n540 & ~n578;
  assign n581 = j3 & n580;
  assign n582 = k3 & n579;
  assign n583 = ~n581 & ~n582;
  assign n584 = p3 & n540;
  assign n585 = ~n583 & n584;
  assign n586 = ~p3 & ~n540;
  assign n587 = ~n583 & n586;
  assign n588 = h0 & ~n578;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n585 & n589;
  assign n591 = q3 & n540;
  assign n592 = ~n590 & n591;
  assign n593 = ~q3 & ~n540;
  assign n594 = ~n590 & n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = ~r3 & ~s3;
  assign n597 = ~n540 & n596;
  assign n598 = ~n595 & n597;
  assign n599 = r3 & s3;
  assign n600 = n540 & n599;
  assign n601 = ~n595 & n600;
  assign n602 = ~n598 & ~n601;
  assign n603 = n526 & n540;
  assign n604 = t3 & ~n526;
  assign n605 = n602 & n604;
  assign n606 = ~t3 & ~n526;
  assign n607 = ~n602 & n606;
  assign n608 = ~n603 & ~n607;
  assign a9 = n605 | ~n608;
  assign n610 = p3 & q3;
  assign n611 = r3 & n610;
  assign n612 = s3 & n611;
  assign n613 = t3 & n612;
  assign n614 = n3 & ~o3;
  assign n615 = ~p3 & n614;
  assign n616 = ~q3 & n615;
  assign n617 = ~r3 & n616;
  assign n618 = ~s3 & n617;
  assign n619 = ~t3 & n618;
  assign n620 = q0 & n368;
  assign n621 = m0 & n613;
  assign n622 = k0 & n619;
  assign n623 = s0 & n567;
  assign n624 = n0 & q5;
  assign n625 = n5 & p0;
  assign n626 = l5 & u0;
  assign n627 = t0 & v4;
  assign n628 = g4 & r0;
  assign n629 = l0 & l3;
  assign n630 = ~n628 & ~n629;
  assign n631 = ~n627 & n630;
  assign n632 = ~n626 & n631;
  assign n633 = ~n625 & n632;
  assign n634 = ~n624 & n633;
  assign n635 = o0 & n526;
  assign n636 = n634 & ~n635;
  assign n637 = ~n623 & n636;
  assign n638 = ~n622 & n637;
  assign n639 = ~n621 & n638;
  assign b6 = n620 | ~n639;
  assign n641 = ~t1 & ~n459;
  assign n642 = t1 & n459;
  assign n643 = ~n464 & ~n642;
  assign n644 = ~n641 & n643;
  assign n645 = ~u1 & n435;
  assign n646 = n644 & n645;
  assign n647 = y2 & n465;
  assign n648 = u1 & n435;
  assign n649 = ~n644 & n648;
  assign n650 = ~n647 & ~n649;
  assign b7 = n646 | ~n650;
  assign n652 = ~w2 & ~x2;
  assign n653 = ~y2 & n652;
  assign n654 = ~z2 & n653;
  assign n655 = ~n477 & n654;
  assign n656 = n477 & ~n490;
  assign b8 = n655 | n656;
  assign n658 = ~n369 & ~n556;
  assign n659 = ~n369 & ~v10;
  assign n660 = ~n557 & ~n659;
  assign n661 = ~n658 & n660;
  assign n662 = ~z & ~n661;
  assign n663 = ~f0 & ~p5;
  assign n664 = ~q5 & n663;
  assign n665 = ~n554 & n664;
  assign n666 = ~r5 & n664;
  assign n667 = ~n551 & n663;
  assign n668 = ~f0 & ~n557;
  assign n669 = ~f0 & ~n550;
  assign n670 = ~f0 & ~s4;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n668 & n671;
  assign n673 = ~n667 & n672;
  assign n674 = ~n666 & n673;
  assign n675 = ~n665 & n674;
  assign n676 = ~z & n661;
  assign n677 = ~u3 & n675;
  assign n678 = n662 & n677;
  assign n679 = l3 & n676;
  assign n680 = u3 & ~n675;
  assign n681 = n662 & n680;
  assign n682 = ~n679 & ~n681;
  assign b9 = n678 | ~n682;
  assign n684 = r1 & n478;
  assign n685 = n503 & ~n684;
  assign n686 = r1 & v0;
  assign n687 = n478 & n686;
  assign n688 = v6 & n503;
  assign n689 = n423 & ~n688;
  assign n690 = ~n687 & n689;
  assign n691 = v0 & n690;
  assign n692 = n685 & n691;
  assign n693 = ~v0 & n690;
  assign n694 = ~n685 & n693;
  assign c6 = n692 | n694;
  assign n696 = u1 & ~n459;
  assign n697 = n644 & n696;
  assign n698 = ~u1 & n459;
  assign n699 = n644 & n698;
  assign n700 = k & n450;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n697 & n701;
  assign n703 = v1 & ~n434;
  assign n704 = n702 & n703;
  assign n705 = ~v1 & ~n434;
  assign n706 = ~n702 & n705;
  assign n707 = z2 & n434;
  assign n708 = ~b & ~n707;
  assign n709 = ~n706 & n708;
  assign c7 = n704 | ~n709;
  assign n711 = w2 & x2;
  assign n712 = y2 & n711;
  assign n713 = z2 & n712;
  assign c8 = ~n477 & n713;
  assign n715 = ~g0 & n537;
  assign n716 = u3 & n675;
  assign n717 = ~n715 & n716;
  assign n718 = n677 & n715;
  assign n719 = ~n717 & ~n718;
  assign n720 = v3 & n719;
  assign n721 = n662 & n720;
  assign n722 = ~v3 & ~n719;
  assign n723 = n662 & n722;
  assign n724 = m3 & n676;
  assign n725 = ~n723 & ~n724;
  assign c9 = n721 | ~n725;
  assign n727 = v0 & ~n685;
  assign n728 = w0 & n690;
  assign n729 = ~n727 & n728;
  assign n730 = ~w0 & n690;
  assign n731 = n727 & n730;
  assign d6 = n729 | n731;
  assign n733 = ~v1 & ~n459;
  assign n734 = v1 & n459;
  assign n735 = ~n702 & ~n734;
  assign n736 = ~n733 & n735;
  assign n737 = ~w1 & ~n434;
  assign n738 = n736 & n737;
  assign n739 = w1 & ~n434;
  assign n740 = ~n736 & n739;
  assign n741 = a3 & n434;
  assign n742 = ~b & ~n741;
  assign n743 = ~n740 & n742;
  assign d7 = n738 | ~n743;
  assign n745 = t2 & n490;
  assign n746 = n514 & n745;
  assign n747 = j & ~n510;
  assign n748 = ~t2 & ~n490;
  assign n749 = n514 & n748;
  assign n750 = ~n747 & ~n749;
  assign n751 = ~n746 & n750;
  assign n752 = ~w2 & ~n477;
  assign n753 = ~n751 & n752;
  assign n754 = w2 & ~n477;
  assign n755 = n751 & n754;
  assign d8 = n753 | n755;
  assign n757 = ~v3 & ~n715;
  assign n758 = v3 & n715;
  assign n759 = ~n719 & ~n758;
  assign n760 = ~n757 & n759;
  assign n761 = ~w3 & n662;
  assign n762 = n760 & n761;
  assign n763 = n3 & n676;
  assign n764 = w3 & n662;
  assign n765 = ~n760 & n764;
  assign n766 = ~n763 & ~n765;
  assign d9 = n762 | ~n766;
  assign n768 = w0 & ~x0;
  assign n769 = ~d6 & n768;
  assign n770 = n690 & n769;
  assign n771 = x0 & d6;
  assign n772 = ~w0 & x0;
  assign n773 = n690 & n772;
  assign n774 = ~n771 & ~n773;
  assign e6 = n770 | ~n774;
  assign n776 = w1 & ~n459;
  assign n777 = n736 & n776;
  assign n778 = ~w1 & n459;
  assign n779 = n736 & n778;
  assign n780 = ~n777 & ~n779;
  assign n781 = x1 & ~n434;
  assign n782 = n780 & n781;
  assign n783 = ~x1 & ~n434;
  assign n784 = ~n780 & n783;
  assign n785 = b3 & n434;
  assign n786 = ~b & ~n785;
  assign n787 = ~n784 & n786;
  assign e7 = n782 | ~n787;
  assign n789 = n490 & ~n751;
  assign n790 = ~n490 & ~n751;
  assign n791 = ~w2 & n790;
  assign n792 = w2 & n789;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~x2 & ~n477;
  assign n795 = ~n793 & n794;
  assign n796 = x2 & ~n477;
  assign n797 = n793 & n796;
  assign e8 = n795 | n797;
  assign n799 = w3 & ~n715;
  assign n800 = n760 & n799;
  assign n801 = ~w3 & n715;
  assign n802 = n760 & n801;
  assign n803 = i0 & n675;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n800 & n804;
  assign n806 = ~x3 & ~n805;
  assign n807 = x3 & ~n661;
  assign n808 = n805 & n807;
  assign n809 = ~n661 & n806;
  assign n810 = o3 & n661;
  assign n811 = ~z & ~n810;
  assign n812 = ~n809 & n811;
  assign e9 = n808 | ~n812;
  assign n814 = w0 & x0;
  assign n815 = y0 & n814;
  assign n816 = n727 & n815;
  assign n817 = x0 & ~e6;
  assign n818 = n690 & n817;
  assign n819 = ~n816 & n818;
  assign n820 = y0 & n690;
  assign n821 = ~n816 & n820;
  assign f6 = n819 | n821;
  assign n823 = x1 & ~n459;
  assign n824 = ~n780 & n823;
  assign n825 = ~x1 & n459;
  assign n826 = ~n780 & n825;
  assign n827 = k & ~n702;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n824 & n828;
  assign n830 = y1 & n829;
  assign n831 = n435 & n830;
  assign n832 = ~y1 & ~n829;
  assign n833 = n435 & n832;
  assign n834 = c3 & n465;
  assign n835 = ~n833 & ~n834;
  assign f7 = n831 | ~n835;
  assign n837 = n711 & n789;
  assign n838 = n652 & n790;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~y2 & ~n477;
  assign n841 = ~n839 & n840;
  assign n842 = y2 & ~n477;
  assign n843 = n839 & n842;
  assign f8 = n841 | n843;
  assign n845 = x3 & ~n715;
  assign n846 = ~n805 & n845;
  assign n847 = n715 & n806;
  assign n848 = ~n846 & ~n847;
  assign n849 = y3 & ~n661;
  assign n850 = n848 & n849;
  assign n851 = ~y3 & ~n661;
  assign n852 = ~n848 & n851;
  assign n853 = p3 & n661;
  assign n854 = ~z & ~n853;
  assign n855 = ~n852 & n854;
  assign f9 = n850 | ~n855;
  assign n857 = z0 & n690;
  assign n858 = ~n816 & n857;
  assign n859 = ~z0 & n690;
  assign n860 = n816 & n859;
  assign g6 = n858 | n860;
  assign n862 = ~y1 & n459;
  assign n863 = y1 & z1;
  assign n864 = ~n459 & n863;
  assign n865 = ~n829 & n864;
  assign n866 = ~z1 & ~n829;
  assign n867 = n862 & n866;
  assign n868 = ~n865 & ~n867;
  assign n869 = y1 & ~n459;
  assign n870 = ~n434 & n869;
  assign n871 = ~n829 & n870;
  assign n872 = n868 & n871;
  assign n873 = z1 & ~n434;
  assign n874 = n868 & n873;
  assign n875 = ~n862 & n874;
  assign n876 = ~n434 & n459;
  assign n877 = ~n868 & n876;
  assign n878 = n829 & n873;
  assign n879 = d3 & n434;
  assign n880 = ~b & ~n879;
  assign n881 = ~n878 & n880;
  assign n882 = ~n877 & n881;
  assign n883 = ~n875 & n882;
  assign g7 = n872 | ~n883;
  assign n885 = x2 & y2;
  assign n886 = ~z2 & n885;
  assign n887 = n490 & n886;
  assign n888 = ~n793 & n887;
  assign n889 = ~y2 & ~z2;
  assign n890 = e8 & n889;
  assign n891 = ~n490 & n890;
  assign n892 = ~n793 & n891;
  assign n893 = z2 & ~e8;
  assign n894 = ~n477 & n893;
  assign n895 = ~n490 & n894;
  assign n896 = z2 & ~n477;
  assign n897 = n793 & n896;
  assign n898 = ~y2 & z2;
  assign n899 = n490 & n898;
  assign n900 = y2 & z2;
  assign n901 = e8 & n900;
  assign n902 = ~n515 & ~n901;
  assign n903 = ~n899 & n902;
  assign n904 = ~n897 & n903;
  assign n905 = ~n895 & n904;
  assign n906 = ~n892 & n905;
  assign g8 = n888 | ~n906;
  assign n908 = ~y3 & ~n715;
  assign n909 = y3 & n715;
  assign n910 = ~n848 & ~n909;
  assign n911 = ~n908 & n910;
  assign n912 = ~z3 & ~n661;
  assign n913 = n911 & n912;
  assign n914 = z3 & ~n661;
  assign n915 = ~n911 & n914;
  assign n916 = q3 & n661;
  assign n917 = ~z & ~n916;
  assign n918 = ~n915 & n917;
  assign g9 = n913 | ~n918;
  assign n920 = z0 & n816;
  assign n921 = a1 & n690;
  assign n922 = ~n920 & n921;
  assign n923 = ~a1 & n690;
  assign n924 = n920 & n923;
  assign h6 = n922 | n924;
  assign n926 = a2 & ~n434;
  assign n927 = n868 & n926;
  assign n928 = ~a2 & ~n434;
  assign n929 = ~n868 & n928;
  assign n930 = e3 & n434;
  assign n931 = ~b & ~n930;
  assign n932 = ~n929 & n931;
  assign h7 = n927 | ~n932;
  assign n934 = u2 & n790;
  assign n935 = v2 & n789;
  assign n936 = ~n934 & ~n935;
  assign n937 = a3 & ~n477;
  assign n938 = n936 & n937;
  assign n939 = ~a3 & ~n477;
  assign n940 = ~n936 & n939;
  assign n941 = ~n515 & ~n940;
  assign h8 = n938 | ~n941;
  assign n943 = ~y3 & ~z3;
  assign n944 = ~n848 & n943;
  assign n945 = n806 & n944;
  assign n946 = y3 & z3;
  assign n947 = ~n715 & n946;
  assign n948 = ~n848 & n947;
  assign n949 = i0 & ~n805;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n945 & n950;
  assign n952 = a4 & n951;
  assign n953 = n662 & n952;
  assign n954 = ~a4 & ~n951;
  assign n955 = n662 & n954;
  assign n956 = r3 & n676;
  assign n957 = ~n955 & ~n956;
  assign h9 = n953 | ~n957;
  assign n959 = a1 & ~b1;
  assign n960 = ~h6 & n959;
  assign n961 = n690 & n960;
  assign n962 = b1 & h6;
  assign n963 = ~a1 & b1;
  assign n964 = n690 & n963;
  assign n965 = ~n962 & ~n964;
  assign i6 = n961 | ~n965;
  assign i7 = b | ~b2;
  assign n968 = a3 & n490;
  assign n969 = ~n936 & n968;
  assign n970 = ~a3 & ~n490;
  assign n971 = ~n936 & n970;
  assign n972 = j & ~n751;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n969 & n973;
  assign n975 = b3 & ~n477;
  assign n976 = n974 & n975;
  assign n977 = ~b3 & ~n477;
  assign n978 = ~n974 & n977;
  assign n979 = ~n515 & ~n978;
  assign i8 = n976 | ~n979;
  assign n981 = ~a4 & n715;
  assign n982 = a4 & b4;
  assign n983 = ~n715 & n982;
  assign n984 = ~n951 & n983;
  assign n985 = ~b4 & ~n951;
  assign n986 = n981 & n985;
  assign n987 = ~n984 & ~n986;
  assign n988 = a4 & ~n661;
  assign n989 = ~n715 & n988;
  assign n990 = ~n951 & n989;
  assign n991 = n987 & n990;
  assign n992 = b4 & ~n661;
  assign n993 = n987 & n992;
  assign n994 = ~n981 & n993;
  assign n995 = ~n661 & n715;
  assign n996 = ~n987 & n995;
  assign n997 = n951 & n992;
  assign n998 = s3 & n661;
  assign n999 = ~z & ~n998;
  assign n1000 = ~n997 & n999;
  assign n1001 = ~n996 & n1000;
  assign n1002 = ~n994 & n1001;
  assign i9 = n991 | ~n1002;
  assign n1004 = a1 & b1;
  assign n1005 = c1 & n1004;
  assign n1006 = n920 & n1005;
  assign n1007 = b1 & ~i6;
  assign n1008 = n690 & n1007;
  assign n1009 = ~n1006 & n1008;
  assign n1010 = c1 & n690;
  assign n1011 = ~n1006 & n1010;
  assign j6 = n1009 | n1011;
  assign n1013 = b2 & ~c2;
  assign n1014 = ~b2 & c2;
  assign n1015 = ~b & ~n1014;
  assign j7 = n1013 | ~n1015;
  assign n1017 = b3 & n490;
  assign n1018 = ~n974 & n1017;
  assign n1019 = ~b3 & ~n490;
  assign n1020 = ~n974 & n1019;
  assign n1021 = ~n1018 & ~n1020;
  assign n1022 = ~c3 & ~n477;
  assign n1023 = ~n1021 & n1022;
  assign n1024 = c3 & ~n477;
  assign n1025 = n1021 & n1024;
  assign j8 = n1023 | n1025;
  assign n1027 = c4 & ~n661;
  assign n1028 = n987 & n1027;
  assign n1029 = ~c4 & ~n661;
  assign n1030 = ~n987 & n1029;
  assign n1031 = t3 & n661;
  assign n1032 = ~z & ~n1031;
  assign n1033 = ~n1030 & n1032;
  assign j9 = n1028 | ~n1033;
  assign n1035 = d1 & n690;
  assign n1036 = ~n1006 & n1035;
  assign n1037 = ~d1 & n690;
  assign n1038 = n1006 & n1037;
  assign k6 = n1036 | n1038;
  assign n1040 = b2 & c2;
  assign n1041 = ~d2 & n1040;
  assign n1042 = d2 & ~n1040;
  assign n1043 = ~b & ~n1042;
  assign k7 = n1041 | ~n1043;
  assign n1045 = c3 & d3;
  assign n1046 = ~c3 & ~d3;
  assign n1047 = ~n490 & n1046;
  assign n1048 = ~n1021 & n1047;
  assign n1049 = n490 & ~n1021;
  assign n1050 = n1045 & n1049;
  assign n1051 = ~n1048 & ~n1050;
  assign n1052 = c3 & n490;
  assign n1053 = ~n1021 & n1052;
  assign n1054 = ~n1045 & n1053;
  assign n1055 = d3 & ~j8;
  assign n1056 = ~n477 & n1055;
  assign n1057 = n1051 & n1056;
  assign n1058 = d3 & n490;
  assign n1059 = ~n1045 & n1058;
  assign n1060 = j8 & n1045;
  assign n1061 = j8 & ~n1051;
  assign n1062 = ~n515 & ~n1061;
  assign n1063 = ~n1060 & n1062;
  assign n1064 = ~n1059 & n1063;
  assign n1065 = ~n1057 & n1064;
  assign k8 = n1054 | ~n1065;
  assign k9 = z | ~d4;
  assign n1068 = d2 & n1040;
  assign n1069 = ~l & q1;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = g2 & ~n1070;
  assign n1072 = ~l & ~p1;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = e2 & ~n1073;
  assign n1075 = n2 & n1074;
  assign n1076 = ~n423 & ~n477;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1074 & n1077;
  assign n1079 = n1071 & n1078;
  assign n1080 = ~n1072 & n1078;
  assign n1081 = e2 & n1078;
  assign n1082 = s1 & ~n1077;
  assign n1083 = ~b & ~n1082;
  assign n1084 = ~n1081 & n1083;
  assign n1085 = ~n1080 & n1084;
  assign l7 = n1079 | ~n1085;
  assign n1087 = e3 & ~n477;
  assign n1088 = n1051 & n1087;
  assign n1089 = ~e3 & ~n477;
  assign n1090 = ~n1051 & n1089;
  assign n1091 = ~n515 & ~n1090;
  assign l8 = n1088 | ~n1091;
  assign n1093 = d4 & ~e4;
  assign n1094 = ~d4 & e4;
  assign n1095 = ~z & ~n1094;
  assign l9 = n1093 | ~n1095;
  assign n1097 = ~f2 & n1077;
  assign n1098 = n1074 & n1097;
  assign n1099 = f2 & n1078;
  assign n1100 = t1 & ~n1077;
  assign n1101 = ~b & ~n1100;
  assign n1102 = ~n1099 & n1101;
  assign m7 = n1098 | ~n1102;
  assign n1104 = ~f3 & ~n526;
  assign n1105 = ~n567 & n1104;
  assign n1106 = f3 & ~n526;
  assign n1107 = n567 & n1106;
  assign m8 = n1105 | n1107;
  assign n1109 = ~f4 & n360;
  assign n1110 = f4 & ~n360;
  assign n1111 = ~z & ~n1110;
  assign m9 = n1109 | ~n1111;
  assign n1113 = g2 & n1070;
  assign n1114 = ~g2 & ~n1070;
  assign n1115 = ~b & ~n1114;
  assign n7 = n1113 | ~n1115;
  assign n1117 = ~f3 & n540;
  assign n1118 = f3 & ~n540;
  assign n1119 = ~n567 & ~n1118;
  assign n1120 = ~n1117 & n1119;
  assign n1121 = g3 & ~n526;
  assign n1122 = ~n1120 & n1121;
  assign n1123 = ~g3 & ~n526;
  assign n1124 = n1120 & n1123;
  assign n8 = n1122 | n1124;
  assign n1126 = ~n313 & ~n526;
  assign n1127 = ~n368 & ~n1126;
  assign n1128 = ~n367 & n1127;
  assign n1129 = n364 & n1128;
  assign n1130 = ~n365 & n1128;
  assign n1131 = g4 & n1128;
  assign n1132 = u3 & ~n1127;
  assign n1133 = ~z & ~n1132;
  assign n1134 = ~n1131 & n1133;
  assign n1135 = ~n1130 & n1134;
  assign n9 = n1129 | ~n1135;
  assign n1137 = n423 & ~n453;
  assign n1138 = ~n502 & n1137;
  assign n1139 = ~h1 & ~n502;
  assign o6 = n1138 | n1139;
  assign n1141 = f2 & n1074;
  assign n1142 = ~h2 & n1077;
  assign n1143 = n1141 & n1142;
  assign n1144 = h2 & n1077;
  assign n1145 = ~n1141 & n1144;
  assign n1146 = u1 & ~n1077;
  assign n1147 = ~b & ~n1146;
  assign n1148 = ~n1145 & n1147;
  assign o7 = n1143 | ~n1148;
  assign n1150 = n540 & ~n567;
  assign n1151 = n522 & n1150;
  assign n1152 = ~n540 & ~n567;
  assign n1153 = n541 & n1152;
  assign n1154 = q5 & ~n567;
  assign n1155 = n528 & n1154;
  assign n1156 = ~n1153 & ~n1155;
  assign n1157 = ~n1151 & n1156;
  assign n1158 = ~h3 & ~n526;
  assign n1159 = ~n1157 & n1158;
  assign n1160 = h3 & ~n526;
  assign n1161 = n1157 & n1160;
  assign o8 = n1159 | n1161;
  assign n1163 = ~h4 & n367;
  assign n1164 = n1127 & n1163;
  assign n1165 = h4 & n1128;
  assign n1166 = v3 & ~n1127;
  assign n1167 = ~z & ~n1166;
  assign n1168 = ~n1165 & n1167;
  assign o9 = n1164 | ~n1168;
  assign n1170 = n423 & n6;
  assign n1171 = ~n452 & n1170;
  assign n1172 = ~i1 & n6;
  assign p6 = n1171 | n1172;
  assign n1174 = h2 & i2;
  assign n1175 = n1141 & n1174;
  assign n1176 = n1144 & ~n1175;
  assign n1177 = n1141 & n1176;
  assign n1178 = i2 & n1077;
  assign n1179 = ~n1175 & n1178;
  assign n1180 = v1 & ~n1077;
  assign n1181 = ~b & ~n1180;
  assign n1182 = ~n1179 & n1181;
  assign p7 = n1177 | ~n1182;
  assign n1184 = ~i3 & ~n526;
  assign n1185 = n571 & n1184;
  assign n1186 = i3 & ~n526;
  assign n1187 = ~n571 & n1186;
  assign n1188 = ~n603 & ~n1187;
  assign p8 = n1185 | ~n1188;
  assign n1190 = i4 & n363;
  assign n1191 = ~i4 & ~n363;
  assign n1192 = ~z & ~n1191;
  assign p9 = n1190 | ~n1192;
  assign n1194 = j1 & n423;
  assign n1195 = n1077 & n1194;
  assign n1196 = n421 & ~n477;
  assign n1197 = ~j1 & n423;
  assign n1198 = ~n1077 & n1197;
  assign n1199 = ~n1196 & ~n1198;
  assign q6 = n1195 | ~n1199;
  assign n1201 = j2 & n1077;
  assign n1202 = ~n1175 & n1201;
  assign n1203 = ~j2 & n1077;
  assign n1204 = n1175 & n1203;
  assign n1205 = w1 & ~n1077;
  assign n1206 = ~b & ~n1205;
  assign n1207 = ~n1204 & n1206;
  assign q7 = n1202 | ~n1207;
  assign n1209 = ~l3 & ~m3;
  assign n1210 = ~n3 & n1209;
  assign n1211 = ~o3 & n1210;
  assign n1212 = ~n526 & n1211;
  assign n1213 = n526 & ~n540;
  assign q8 = n1212 | n1213;
  assign n1215 = h4 & n367;
  assign n1216 = ~j4 & n1127;
  assign n1217 = n1215 & n1216;
  assign n1218 = j4 & n1127;
  assign n1219 = ~n1215 & n1218;
  assign n1220 = w3 & ~n1127;
  assign n1221 = ~z & ~n1220;
  assign n1222 = ~n1219 & n1221;
  assign q9 = n1217 | ~n1222;
  assign n1224 = j2 & n1175;
  assign n1225 = ~l & ~n1224;
  assign n1226 = k2 & ~n1225;
  assign n1227 = n1077 & ~n1226;
  assign n1228 = ~n1225 & n1227;
  assign n1229 = k2 & n1077;
  assign n1230 = ~n1226 & n1229;
  assign n1231 = x1 & ~n1077;
  assign n1232 = ~b & ~n1231;
  assign n1233 = ~n1230 & n1232;
  assign r7 = n1228 | ~n1233;
  assign n1235 = l3 & m3;
  assign n1236 = n3 & n1235;
  assign n1237 = o3 & n1236;
  assign r8 = ~n526 & n1237;
  assign n1239 = j4 & k4;
  assign n1240 = n1215 & n1239;
  assign n1241 = n1218 & ~n1240;
  assign n1242 = n1215 & n1241;
  assign n1243 = k4 & n1127;
  assign n1244 = ~n1240 & n1243;
  assign n1245 = x3 & ~n1127;
  assign n1246 = ~z & ~n1245;
  assign n1247 = ~n1244 & n1246;
  assign r9 = n1242 | ~n1247;
  assign n1249 = m & e3;
  assign n1250 = n & a3;
  assign n1251 = o & t2;
  assign n1252 = s & o2;
  assign n1253 = t & j2;
  assign n1254 = u & g2;
  assign n1255 = p & a2;
  assign n1256 = q & x1;
  assign n1257 = r & u1;
  assign n1258 = v & d1;
  assign n1259 = w & y0;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1257 & n1260;
  assign n1262 = ~n1256 & n1261;
  assign n1263 = ~n1255 & n1262;
  assign n1264 = ~n1254 & n1263;
  assign n1265 = ~n1253 & n1264;
  assign n1266 = ~n1252 & n1265;
  assign n1267 = ~n1251 & n1266;
  assign n1268 = ~n1250 & n1267;
  assign s5 = n1249 | ~n1268;
  assign n1270 = e3 & n1045;
  assign n1271 = y2 & ~z2;
  assign n1272 = ~a3 & n1271;
  assign n1273 = ~b3 & n1272;
  assign n1274 = ~c3 & n1273;
  assign n1275 = ~d3 & n1274;
  assign n1276 = ~e3 & n1275;
  assign n1277 = n453 & ~n1276;
  assign n1278 = n423 & n477;
  assign n1279 = n453 & n1278;
  assign n1280 = n478 & ~n1270;
  assign n1281 = n478 & ~n1277;
  assign n1282 = ~n424 & ~n1281;
  assign n1283 = ~n1280 & n1282;
  assign s6 = n1279 | ~n1283;
  assign n1285 = l2 & n1077;
  assign n1286 = ~n1226 & n1285;
  assign n1287 = ~l2 & n1077;
  assign n1288 = n1226 & n1287;
  assign n1289 = y1 & ~n1077;
  assign n1290 = ~b & ~n1289;
  assign n1291 = ~n1288 & n1290;
  assign s7 = n1286 | ~n1291;
  assign n1293 = ~l3 & ~n526;
  assign n1294 = ~n578 & n1293;
  assign n1295 = l3 & ~n526;
  assign n1296 = n578 & n1295;
  assign s8 = n1294 | n1296;
  assign n1298 = l4 & n1127;
  assign n1299 = ~n1240 & n1298;
  assign n1300 = ~l4 & n1127;
  assign n1301 = n1240 & n1300;
  assign n1302 = y3 & ~n1127;
  assign n1303 = ~z & ~n1302;
  assign n1304 = ~n1301 & n1303;
  assign s9 = n1299 | ~n1304;
  assign n1306 = m & d3;
  assign n1307 = n & z2;
  assign n1308 = o & s2;
  assign n1309 = s & m2;
  assign n1310 = t & i2;
  assign n1311 = u & d2;
  assign n1312 = p & z1;
  assign n1313 = q & w1;
  assign n1314 = r & t1;
  assign n1315 = v & c1;
  assign n1316 = w & x0;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~n1314 & n1317;
  assign n1319 = ~n1313 & n1318;
  assign n1320 = ~n1312 & n1319;
  assign n1321 = ~n1311 & n1320;
  assign n1322 = ~n1310 & n1321;
  assign n1323 = ~n1309 & n1322;
  assign n1324 = ~n1308 & n1323;
  assign n1325 = ~n1307 & n1324;
  assign t5 = n1306 | ~n1325;
  assign n1327 = n1 & n423;
  assign n1328 = d1 & v6;
  assign n1329 = n1006 & n1328;
  assign n1330 = n423 & n1329;
  assign n1331 = d1 & ~r1;
  assign n1332 = v6 & n1331;
  assign n1333 = n423 & n1332;
  assign n1334 = c & v6;
  assign n1335 = n423 & n1334;
  assign n1336 = ~n1278 & ~n1327;
  assign n1337 = ~n1281 & n1336;
  assign n1338 = ~n1335 & n1337;
  assign n1339 = ~n1333 & n1338;
  assign t6 = n1330 | ~n1339;
  assign n1341 = l2 & n1226;
  assign n1342 = ~m2 & n1077;
  assign n1343 = n1341 & n1342;
  assign n1344 = m2 & n1077;
  assign n1345 = ~n1341 & n1344;
  assign n1346 = z1 & ~n1077;
  assign n1347 = ~b & ~n1346;
  assign n1348 = ~n1345 & n1347;
  assign t7 = n1343 | ~n1348;
  assign n1350 = ~l3 & n580;
  assign n1351 = l3 & n579;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~m3 & ~n526;
  assign n1354 = ~n1352 & n1353;
  assign n1355 = m3 & ~n526;
  assign n1356 = n1352 & n1355;
  assign t8 = n1354 | n1356;
  assign n1358 = l4 & n1240;
  assign n1359 = ~j0 & ~n1358;
  assign n1360 = m4 & ~n1359;
  assign n1361 = n1127 & ~n1360;
  assign n1362 = ~n1359 & n1361;
  assign n1363 = m4 & n1127;
  assign n1364 = ~n1360 & n1363;
  assign n1365 = z3 & ~n1127;
  assign n1366 = ~z & ~n1365;
  assign n1367 = ~n1364 & n1366;
  assign t9 = n1362 | ~n1367;
  assign n1369 = m & c3;
  assign n1370 = n & y2;
  assign n1371 = o & r2;
  assign n1372 = s & l2;
  assign n1373 = t & h2;
  assign n1374 = u & c2;
  assign n1375 = p & y1;
  assign n1376 = q & v1;
  assign n1377 = r & s1;
  assign n1378 = v & b1;
  assign n1379 = w & w0;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~n1377 & n1380;
  assign n1382 = ~n1376 & n1381;
  assign n1383 = ~n1375 & n1382;
  assign n1384 = ~n1374 & n1383;
  assign n1385 = ~n1373 & n1384;
  assign n1386 = ~n1372 & n1385;
  assign n1387 = ~n1371 & n1386;
  assign n1388 = ~n1370 & n1387;
  assign u5 = n1369 | ~n1388;
  assign n1390 = ~m1 & ~v6;
  assign n1391 = n423 & n1390;
  assign n1392 = l1 & ~s6;
  assign n1393 = n423 & n1392;
  assign n1394 = n478 & n1276;
  assign n1395 = ~n1393 & ~n1394;
  assign u6 = n1391 | ~n1395;
  assign n1397 = f2 & h2;
  assign n1398 = i2 & n1397;
  assign n1399 = j2 & n1398;
  assign n1400 = k2 & n1399;
  assign n1401 = l2 & n1400;
  assign n1402 = m2 & n1401;
  assign n1403 = o2 & n1402;
  assign n1404 = n1077 & n1403;
  assign n1405 = b & f2;
  assign n1406 = h2 & n1405;
  assign n1407 = i2 & n1406;
  assign n1408 = j2 & n1407;
  assign n1409 = k2 & n1408;
  assign n1410 = l2 & n1409;
  assign n1411 = m2 & n1410;
  assign n1412 = o2 & n1411;
  assign u7 = n1404 | n1412;
  assign n1414 = n579 & n1235;
  assign n1415 = n580 & n1209;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n3 & ~n526;
  assign n1418 = ~n1416 & n1417;
  assign n1419 = n3 & ~n526;
  assign n1420 = n1416 & n1419;
  assign u8 = n1418 | n1420;
  assign n1422 = n4 & n1127;
  assign n1423 = ~n1360 & n1422;
  assign n1424 = ~n4 & n1127;
  assign n1425 = n1360 & n1424;
  assign n1426 = a4 & ~n1127;
  assign n1427 = ~z & ~n1426;
  assign n1428 = ~n1425 & n1427;
  assign u9 = n1423 | ~n1428;
  assign n1430 = m & b3;
  assign n1431 = n & x2;
  assign n1432 = o & q2;
  assign n1433 = s & k2;
  assign n1434 = t & f2;
  assign n1435 = u & b2;
  assign n1436 = q & r1;
  assign n1437 = p & p1;
  assign n1438 = r & m1;
  assign n1439 = v & a1;
  assign n1440 = w & v0;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~n1438 & n1441;
  assign n1443 = ~n1437 & n1442;
  assign n1444 = ~n1436 & n1443;
  assign n1445 = ~n1435 & n1444;
  assign n1446 = ~n1434 & n1445;
  assign n1447 = ~n1433 & n1446;
  assign n1448 = ~n1432 & n1447;
  assign n1449 = ~n1431 & n1448;
  assign v5 = n1430 | ~n1449;
  assign n1451 = m2 & n1341;
  assign n1452 = ~o2 & n1077;
  assign n1453 = n1451 & n1452;
  assign n1454 = o2 & n1077;
  assign n1455 = ~n1451 & n1454;
  assign n1456 = a2 & ~n1077;
  assign n1457 = ~b & ~n1456;
  assign n1458 = ~n1455 & n1457;
  assign v7 = n1453 | ~n1458;
  assign n1460 = m3 & n3;
  assign n1461 = ~o3 & n1460;
  assign n1462 = n540 & n1461;
  assign n1463 = ~n1352 & n1462;
  assign n1464 = ~n3 & ~o3;
  assign n1465 = t8 & n1464;
  assign n1466 = ~n540 & n1465;
  assign n1467 = ~n1352 & n1466;
  assign n1468 = o3 & ~t8;
  assign n1469 = ~n526 & n1468;
  assign n1470 = ~n540 & n1469;
  assign n1471 = o3 & ~n526;
  assign n1472 = n1352 & n1471;
  assign n1473 = ~n3 & o3;
  assign n1474 = n540 & n1473;
  assign n1475 = n3 & o3;
  assign n1476 = t8 & n1475;
  assign n1477 = ~n603 & ~n1476;
  assign n1478 = ~n1474 & n1477;
  assign n1479 = ~n1472 & n1478;
  assign n1480 = ~n1470 & n1479;
  assign n1481 = ~n1467 & n1480;
  assign v8 = n1463 | ~n1481;
  assign n1483 = n4 & n1360;
  assign n1484 = ~o4 & n1127;
  assign n1485 = n1483 & n1484;
  assign n1486 = o4 & n1127;
  assign n1487 = ~n1483 & n1486;
  assign n1488 = b4 & ~n1127;
  assign n1489 = ~z & ~n1488;
  assign n1490 = ~n1487 & n1489;
  assign v9 = n1485 | ~n1490;
  assign n1492 = o & n1270;
  assign n1493 = s & n1075;
  assign n1494 = m & n1276;
  assign n1495 = u & n510;
  assign n1496 = n & w2;
  assign n1497 = t & e2;
  assign n1498 = p & q1;
  assign n1499 = r & n1;
  assign n1500 = w & l1;
  assign n1501 = v & z0;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1499 & n1502;
  assign n1504 = ~n1498 & n1503;
  assign n1505 = ~n1497 & n1504;
  assign n1506 = ~n1496 & n1505;
  assign n1507 = q & n477;
  assign n1508 = n1506 & ~n1507;
  assign n1509 = ~n1495 & n1508;
  assign n1510 = ~n1494 & n1509;
  assign n1511 = ~n1493 & n1510;
  assign w5 = n1492 | ~n1511;
  assign n1513 = ~e & ~n1327;
  assign n1514 = ~e & ~l1;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~d & m1;
  assign n1517 = ~d & ~n1327;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1515 & ~n1518;
  assign n1520 = ~b & ~q1;
  assign n1521 = ~r1 & n1520;
  assign n1522 = ~b & ~p1;
  assign n1523 = ~r1 & n1522;
  assign n1524 = ~q1 & n1522;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1521 & n1525;
  assign n1527 = r1 & ~n1526;
  assign n1528 = n1519 & n1527;
  assign n1529 = p1 & ~n1526;
  assign n1530 = n1518 & n1529;
  assign n1531 = q1 & ~n1526;
  assign n1532 = n1515 & n1531;
  assign n1533 = ~n1530 & ~n1532;
  assign y6 = n1528 | ~n1533;
  assign n1535 = n1519 & n1531;
  assign n1536 = n1518 & n1527;
  assign n1537 = n1515 & n1529;
  assign n1538 = ~n1536 & ~n1537;
  assign x6 = n1535 | ~n1538;
  assign n1540 = ~p1 & n1518;
  assign n1541 = n1515 & n1540;
  assign n1542 = ~y6 & ~x6;
  assign w6 = n1541 | n1542;
  assign n1544 = j1 & n1075;
  assign n1545 = ~a & n1544;
  assign n1546 = p2 & ~n1544;
  assign w7 = n1545 | n1546;
  assign n1548 = p3 & ~n526;
  assign n1549 = n583 & n1548;
  assign n1550 = ~p3 & ~n526;
  assign n1551 = ~n583 & n1550;
  assign n1552 = ~n603 & ~n1551;
  assign w8 = n1549 | ~n1552;
  assign n1554 = h4 & j4;
  assign n1555 = k4 & n1554;
  assign n1556 = l4 & n1555;
  assign n1557 = m4 & n1556;
  assign n1558 = n4 & n1557;
  assign n1559 = o4 & n1558;
  assign n1560 = q4 & n1559;
  assign n1561 = n1127 & n1560;
  assign n1562 = z & h4;
  assign n1563 = j4 & n1562;
  assign n1564 = k4 & n1563;
  assign n1565 = l4 & n1564;
  assign n1566 = m4 & n1565;
  assign n1567 = n4 & n1566;
  assign n1568 = o4 & n1567;
  assign n1569 = q4 & n1568;
  assign w9 = n1561 | n1569;
  assign n1571 = t0 & z4;
  assign n1572 = u0 & u4;
  assign n1573 = q0 & q4;
  assign n1574 = l4 & r0;
  assign n1575 = i4 & s0;
  assign n1576 = c4 & n0;
  assign n1577 = o0 & z3;
  assign n1578 = p0 & w3;
  assign n1579 = k0 & t3;
  assign n1580 = l0 & p3;
  assign n1581 = i3 & m0;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~n1579 & n1582;
  assign n1584 = ~n1578 & n1583;
  assign n1585 = ~n1577 & n1584;
  assign n1586 = ~n1576 & n1585;
  assign n1587 = ~n1575 & n1586;
  assign n1588 = ~n1574 & n1587;
  assign n1589 = ~n1573 & n1588;
  assign n1590 = ~n1572 & n1589;
  assign x5 = n1571 | ~n1590;
  assign n1592 = ~q2 & ~n477;
  assign n1593 = ~n510 & n1592;
  assign n1594 = q2 & ~n477;
  assign n1595 = n510 & n1594;
  assign x7 = n1593 | n1595;
  assign n1597 = q3 & ~n526;
  assign n1598 = n590 & n1597;
  assign n1599 = ~q3 & ~n526;
  assign n1600 = ~n590 & n1599;
  assign n1601 = ~n603 & ~n1600;
  assign x8 = n1598 | ~n1601;
  assign n1603 = o4 & n1483;
  assign n1604 = ~q4 & n1127;
  assign n1605 = n1603 & n1604;
  assign n1606 = q4 & n1127;
  assign n1607 = ~n1603 & n1606;
  assign n1608 = c4 & ~n1127;
  assign n1609 = ~z & ~n1608;
  assign n1610 = ~n1607 & n1609;
  assign x9 = n1605 | ~n1610;
  assign n1612 = t0 & y4;
  assign n1613 = t4 & u0;
  assign n1614 = o4 & q0;
  assign n1615 = k4 & r0;
  assign n1616 = f4 & s0;
  assign n1617 = b4 & n0;
  assign n1618 = o0 & y3;
  assign n1619 = p0 & v3;
  assign n1620 = k0 & s3;
  assign n1621 = l0 & o3;
  assign n1622 = h3 & m0;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n1620 & n1623;
  assign n1625 = ~n1619 & n1624;
  assign n1626 = ~n1618 & n1625;
  assign n1627 = ~n1617 & n1626;
  assign n1628 = ~n1616 & n1627;
  assign n1629 = ~n1615 & n1628;
  assign n1630 = ~n1614 & n1629;
  assign n1631 = ~n1613 & n1630;
  assign y5 = n1612 | ~n1631;
  assign n1633 = ~q2 & n490;
  assign n1634 = q2 & ~n490;
  assign n1635 = ~n510 & ~n1634;
  assign n1636 = ~n1633 & n1635;
  assign n1637 = r2 & ~n477;
  assign n1638 = ~n1636 & n1637;
  assign n1639 = ~r2 & ~n477;
  assign n1640 = n1636 & n1639;
  assign y7 = n1638 | n1640;
  assign n1642 = ~r3 & ~n526;
  assign n1643 = ~n595 & n1642;
  assign n1644 = r3 & ~n526;
  assign n1645 = n595 & n1644;
  assign y8 = n1643 | n1645;
  assign n1647 = r5 & n527;
  assign n1648 = n558 & ~n1647;
  assign n1649 = r4 & r5;
  assign n1650 = n527 & n1649;
  assign n1651 = v10 & n558;
  assign n1652 = n313 & ~n1651;
  assign n1653 = ~n1650 & n1652;
  assign n1654 = r4 & n1653;
  assign n1655 = n1648 & n1654;
  assign n1656 = ~r4 & n1653;
  assign n1657 = ~n1648 & n1656;
  assign y9 = n1655 | n1657;
  assign n1659 = t0 & x4;
  assign n1660 = s4 & u0;
  assign n1661 = n4 & q0;
  assign n1662 = j4 & r0;
  assign n1663 = e4 & s0;
  assign n1664 = a4 & n0;
  assign n1665 = o0 & x3;
  assign n1666 = p0 & u3;
  assign n1667 = k0 & r3;
  assign n1668 = l0 & n3;
  assign n1669 = g3 & m0;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = ~n1667 & n1670;
  assign n1672 = ~n1666 & n1671;
  assign n1673 = ~n1665 & n1672;
  assign n1674 = ~n1664 & n1673;
  assign n1675 = ~n1663 & n1674;
  assign n1676 = ~n1662 & n1675;
  assign n1677 = ~n1661 & n1676;
  assign n1678 = ~n1660 & n1677;
  assign z5 = n1659 | ~n1678;
  assign n1680 = ~s1 & n450;
  assign n1681 = n435 & n1680;
  assign n1682 = w2 & n465;
  assign n1683 = s1 & ~n450;
  assign n1684 = n435 & n1683;
  assign n1685 = ~n1682 & ~n1684;
  assign z6 = n1681 | ~n1685;
  assign n1687 = n490 & ~n510;
  assign n1688 = n473 & n1687;
  assign n1689 = ~n490 & ~n510;
  assign n1690 = n491 & n1689;
  assign n1691 = q1 & ~n510;
  assign n1692 = n479 & n1691;
  assign n1693 = ~n1690 & ~n1692;
  assign n1694 = ~n1688 & n1693;
  assign n1695 = ~s2 & ~n477;
  assign n1696 = ~n1694 & n1695;
  assign n1697 = s2 & ~n477;
  assign n1698 = n1694 & n1697;
  assign z7 = n1696 | n1698;
  assign n1700 = r3 & n540;
  assign n1701 = ~n595 & n1700;
  assign n1702 = n602 & n1701;
  assign n1703 = s3 & ~y8;
  assign n1704 = ~n526 & n1703;
  assign n1705 = n602 & n1704;
  assign n1706 = s3 & n540;
  assign n1707 = n602 & n1706;
  assign n1708 = s3 & ~n526;
  assign n1709 = n595 & n1708;
  assign n1710 = ~n602 & y8;
  assign n1711 = ~n603 & ~n1710;
  assign n1712 = ~n1709 & n1711;
  assign n1713 = ~n1707 & n1712;
  assign n1714 = ~n1705 & n1713;
  assign z8 = n1702 | ~n1714;
  assign n1716 = r4 & ~n1648;
  assign n1717 = s4 & n1653;
  assign n1718 = ~n1716 & n1717;
  assign n1719 = ~s4 & n1653;
  assign n1720 = n1716 & n1719;
  assign z9 = n1718 | n1720;
  assign n1722 = s4 & ~t4;
  assign n1723 = ~z9 & n1722;
  assign n1724 = n1653 & n1723;
  assign n1725 = t4 & z9;
  assign n1726 = ~s4 & t4;
  assign n1727 = n1653 & n1726;
  assign n1728 = ~n1725 & ~n1727;
  assign a10 = n1724 | ~n1728;
  assign n1730 = ~j5 & ~k5;
  assign n1731 = n527 & n1730;
  assign n1732 = ~z & j5;
  assign n1733 = ~n527 & n1732;
  assign q10 = n1731 | n1733;
  assign n1735 = s4 & t4;
  assign n1736 = u4 & n1735;
  assign n1737 = n1716 & n1736;
  assign n1738 = t4 & ~a10;
  assign n1739 = n1653 & n1738;
  assign n1740 = ~n1737 & n1739;
  assign n1741 = u4 & n1653;
  assign n1742 = ~n1737 & n1741;
  assign b10 = n1740 | n1742;
  assign n1744 = j5 & ~k5;
  assign n1745 = n527 & n1744;
  assign n1746 = k5 & q10;
  assign r10 = n1745 | n1746;
  assign n1748 = v4 & n1653;
  assign n1749 = ~n1737 & n1748;
  assign n1750 = ~v4 & n1653;
  assign n1751 = n1737 & n1750;
  assign c10 = n1749 | n1751;
  assign n1753 = n344 & ~n619;
  assign n1754 = n313 & n526;
  assign n1755 = n344 & n1754;
  assign n1756 = n527 & ~n1753;
  assign n1757 = n527 & ~n613;
  assign n1758 = ~n369 & ~n1757;
  assign n1759 = ~n1756 & n1758;
  assign s10 = n1755 | ~n1759;
  assign n1761 = v4 & n1737;
  assign n1762 = w4 & n1653;
  assign n1763 = ~n1761 & n1762;
  assign n1764 = ~w4 & n1653;
  assign n1765 = n1761 & n1764;
  assign d10 = n1763 | n1765;
  assign n1767 = w4 & x4;
  assign n1768 = y4 & n1767;
  assign n1769 = n1761 & n1768;
  assign n1770 = z4 & v10;
  assign n1771 = n1769 & n1770;
  assign n1772 = n313 & n1771;
  assign n1773 = ~r5 & z4;
  assign n1774 = v10 & n1773;
  assign n1775 = n313 & n1774;
  assign n1776 = a0 & v10;
  assign n1777 = n313 & n1776;
  assign n1778 = ~n314 & ~n1754;
  assign n1779 = ~n1756 & n1778;
  assign n1780 = ~n1777 & n1779;
  assign n1781 = ~n1775 & n1780;
  assign t10 = n1772 | ~n1781;
  assign n1783 = w4 & ~x4;
  assign n1784 = ~d10 & n1783;
  assign n1785 = n1653 & n1784;
  assign n1786 = x4 & d10;
  assign n1787 = ~w4 & x4;
  assign n1788 = n1653 & n1787;
  assign n1789 = ~n1786 & ~n1788;
  assign e10 = n1785 | ~n1789;
  assign n1791 = ~m5 & ~v10;
  assign n1792 = n313 & n1791;
  assign n1793 = l5 & ~s10;
  assign n1794 = n313 & n1793;
  assign n1795 = n527 & n619;
  assign n1796 = ~n1794 & ~n1795;
  assign u10 = n1792 | ~n1796;
  assign n1798 = x4 & ~e10;
  assign n1799 = n1653 & n1798;
  assign n1800 = ~n1769 & n1799;
  assign n1801 = y4 & n1653;
  assign n1802 = ~n1769 & n1801;
  assign f10 = n1800 | n1802;
  assign n1804 = z4 & n1653;
  assign n1805 = ~n1769 & n1804;
  assign n1806 = ~z4 & n1653;
  assign n1807 = n1769 & n1806;
  assign g10 = n1805 | n1807;
  assign n1809 = ~p5 & n317;
  assign n1810 = n320 & n1809;
  assign n1811 = ~x10 & ~y10;
  assign w10 = n1810 | n1811;
  assign h10 = y;
  assign i10 = a5;
  assign l6 = a;
  assign m6 = e1;
  assign r6 = j1;
  assign p10 = g5;
endmodule


