// Benchmark "k2" written by ABC on Tue May 16 16:07:51 2017

module k2 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, r0, s0,
    z0, z1, a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2,
    i1, i2, j1, j2, k1, k2, l1, l2, m1, n1, o1, p1, q1, r1, s1, t0, t1, u0,
    u1, v0, v1, w0, w1, x0, x1, y0, y1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0, p0, q0, r0, s0;
  output z0, z1, a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1,
    h2, i1, i2, j1, j2, k1, k2, l1, l2, m1, n1, o1, p1, q1, r1, s1, t0, t1,
    u0, u1, v0, v1, w0, w1, x0, x1, y0, y1;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n365, n366, n367, n368, n369, n370,
    n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n633, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n857, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1774, n1775, n1776, n1777, n1778, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2156, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2187, n2188, n2189, n2190, n2192, n2193,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2267, n2269, n2270,
    n2271, n2272, n2274, n2275, n2277, n2278, n2279, n2280;
  assign n92 = a & d;
  assign n93 = s & n92;
  assign n94 = t & n93;
  assign n95 = u & n94;
  assign n96 = ~v & n95;
  assign n97 = b0 & n96;
  assign n98 = ~d0 & n97;
  assign n99 = ~e0 & n98;
  assign n100 = ~a & ~e;
  assign n101 = s & n100;
  assign n102 = t & n101;
  assign n103 = u & n102;
  assign n104 = ~v & n103;
  assign n105 = ~b0 & n104;
  assign n106 = c0 & n105;
  assign n107 = d0 & n106;
  assign n108 = ~e0 & n107;
  assign n109 = a & ~f;
  assign n110 = s & n109;
  assign n111 = t & n110;
  assign n112 = u & n111;
  assign n113 = ~v & n112;
  assign n114 = ~b0 & n113;
  assign n115 = ~c0 & n114;
  assign n116 = d0 & n115;
  assign n117 = e0 & n116;
  assign n118 = a & ~l;
  assign n119 = s & n118;
  assign n120 = t & n119;
  assign n121 = ~u & n120;
  assign n122 = ~v & n121;
  assign n123 = a0 & n122;
  assign n124 = c0 & n123;
  assign n125 = ~d0 & n124;
  assign n126 = e0 & n125;
  assign n127 = a & l;
  assign n128 = s & n127;
  assign n129 = t & n128;
  assign n130 = ~u & n129;
  assign n131 = ~v & n130;
  assign n132 = a0 & n131;
  assign n133 = c0 & n132;
  assign n134 = ~d0 & n133;
  assign n135 = e0 & n134;
  assign n136 = a & s;
  assign n137 = t & n136;
  assign n138 = ~u & n137;
  assign n139 = ~v & n138;
  assign n140 = a0 & n139;
  assign n141 = ~c0 & n140;
  assign n142 = d0 & n141;
  assign n143 = ~e0 & n142;
  assign n144 = a & k;
  assign n145 = ~l & n144;
  assign n146 = s & n145;
  assign n147 = t & n146;
  assign n148 = ~u & n147;
  assign n149 = ~v & n148;
  assign n150 = z & n149;
  assign n151 = d0 & n150;
  assign n152 = ~e0 & n151;
  assign n153 = l & n144;
  assign n154 = s & n153;
  assign n155 = t & n154;
  assign n156 = ~u & n155;
  assign n157 = ~v & n156;
  assign n158 = z & n157;
  assign n159 = d0 & n158;
  assign n160 = ~e0 & n159;
  assign n161 = w & n139;
  assign n162 = d0 & n161;
  assign n163 = ~e0 & n162;
  assign n164 = ~t & n128;
  assign n165 = u & n164;
  assign n166 = ~v & n165;
  assign n167 = a0 & n166;
  assign n168 = c0 & n167;
  assign n169 = ~d0 & n168;
  assign n170 = e0 & n169;
  assign n171 = ~t & n119;
  assign n172 = u & n171;
  assign n173 = ~v & n172;
  assign n174 = a0 & n173;
  assign n175 = c0 & n174;
  assign n176 = ~d0 & n175;
  assign n177 = e0 & n176;
  assign n178 = a & ~r;
  assign n179 = s & n178;
  assign n180 = ~t & n179;
  assign n181 = u & n180;
  assign n182 = ~v & n181;
  assign n183 = a0 & n182;
  assign n184 = ~c0 & n183;
  assign n185 = d0 & n184;
  assign n186 = ~e0 & n185;
  assign n187 = a & r;
  assign n188 = s & n187;
  assign n189 = ~t & n188;
  assign n190 = u & n189;
  assign n191 = ~v & n190;
  assign n192 = a0 & n191;
  assign n193 = ~c0 & n192;
  assign n194 = d0 & n193;
  assign n195 = ~e0 & n194;
  assign n196 = a & ~s;
  assign n197 = t & n196;
  assign n198 = u & n197;
  assign n199 = ~v & n198;
  assign n200 = w & n199;
  assign n201 = c0 & n200;
  assign n202 = d0 & n201;
  assign n203 = ~e0 & n202;
  assign n204 = ~s & n109;
  assign n205 = t & n204;
  assign n206 = u & n205;
  assign n207 = ~v & n206;
  assign n208 = w & n207;
  assign n209 = ~c0 & n208;
  assign n210 = d0 & n209;
  assign n211 = ~e0 & n210;
  assign n212 = a & ~c;
  assign n213 = ~d & n212;
  assign n214 = ~s & n213;
  assign n215 = ~t & n214;
  assign n216 = u & n215;
  assign n217 = ~v & n216;
  assign n218 = c0 & n217;
  assign n219 = ~d0 & n218;
  assign n220 = e0 & n219;
  assign n221 = ~t & n196;
  assign n222 = u & n221;
  assign n223 = ~v & n222;
  assign n224 = x & n223;
  assign n225 = ~c0 & n224;
  assign n226 = d0 & n225;
  assign n227 = ~e0 & n226;
  assign n228 = a & c;
  assign n229 = ~d & n228;
  assign n230 = ~s & n229;
  assign n231 = ~t & n230;
  assign n232 = ~u & n231;
  assign n233 = ~v & n232;
  assign n234 = c0 & n233;
  assign n235 = ~d0 & n234;
  assign n236 = e0 & n235;
  assign n237 = a & ~d;
  assign n238 = ~f & n237;
  assign n239 = ~s & n238;
  assign n240 = ~t & n239;
  assign n241 = ~u & n240;
  assign n242 = ~v & n241;
  assign n243 = ~c0 & n242;
  assign n244 = d0 & n243;
  assign n245 = ~e0 & n244;
  assign n246 = l & n109;
  assign n247 = ~p & n246;
  assign n248 = s & n247;
  assign n249 = ~t & n248;
  assign n250 = u & n249;
  assign n251 = v & n250;
  assign n252 = a0 & n251;
  assign n253 = ~c0 & n252;
  assign n254 = ~d0 & n253;
  assign n255 = e0 & n254;
  assign n256 = ~l & n109;
  assign n257 = ~p & n256;
  assign n258 = s & n257;
  assign n259 = ~t & n258;
  assign n260 = u & n259;
  assign n261 = v & n260;
  assign n262 = a0 & n261;
  assign n263 = ~c0 & n262;
  assign n264 = ~d0 & n263;
  assign n265 = e0 & n264;
  assign n266 = k & n109;
  assign n267 = l & n266;
  assign n268 = ~p & n267;
  assign n269 = s & n268;
  assign n270 = ~t & n269;
  assign n271 = u & n270;
  assign n272 = v & n271;
  assign n273 = z & n272;
  assign n274 = ~c0 & n273;
  assign n275 = ~d0 & n274;
  assign n276 = e0 & n275;
  assign n277 = ~l & n266;
  assign n278 = ~p & n277;
  assign n279 = s & n278;
  assign n280 = ~t & n279;
  assign n281 = u & n280;
  assign n282 = v & n281;
  assign n283 = z & n282;
  assign n284 = ~c0 & n283;
  assign n285 = ~d0 & n284;
  assign n286 = e0 & n285;
  assign n287 = ~p & n109;
  assign n288 = s & n287;
  assign n289 = ~t & n288;
  assign n290 = u & n289;
  assign n291 = v & n290;
  assign n292 = w & n291;
  assign n293 = ~c0 & n292;
  assign n294 = ~d0 & n293;
  assign n295 = e0 & n294;
  assign n296 = ~s & n287;
  assign n297 = t & n296;
  assign n298 = u & n297;
  assign n299 = v & n298;
  assign n300 = w & n299;
  assign n301 = ~c0 & n300;
  assign n302 = ~d0 & n301;
  assign i2 = e0 & n302;
  assign n304 = ~s & n127;
  assign n305 = ~t & n304;
  assign n306 = u & n305;
  assign n307 = v & n306;
  assign n308 = a0 & n307;
  assign n309 = ~d0 & n308;
  assign n310 = e0 & n309;
  assign n311 = ~s & n118;
  assign n312 = ~t & n311;
  assign n313 = u & n312;
  assign n314 = v & n313;
  assign n315 = a0 & n314;
  assign n316 = ~d0 & n315;
  assign n317 = e0 & n316;
  assign n318 = ~s & n153;
  assign n319 = ~t & n318;
  assign n320 = u & n319;
  assign n321 = v & n320;
  assign n322 = z & n321;
  assign n323 = ~d0 & n322;
  assign n324 = e0 & n323;
  assign n325 = ~s & n145;
  assign n326 = ~t & n325;
  assign n327 = u & n326;
  assign n328 = v & n327;
  assign n329 = z & n328;
  assign n330 = ~d0 & n329;
  assign n331 = e0 & n330;
  assign n332 = v & n222;
  assign n333 = w & n332;
  assign n334 = ~d0 & n333;
  assign n335 = e0 & n334;
  assign n336 = ~n331 & ~n335;
  assign n337 = ~n324 & n336;
  assign n338 = ~n317 & n337;
  assign n339 = ~n310 & n338;
  assign n340 = ~i2 & n339;
  assign n341 = ~n295 & n340;
  assign n342 = ~n286 & n341;
  assign n343 = ~n276 & n342;
  assign n344 = ~n265 & n343;
  assign n345 = ~n255 & n344;
  assign n346 = ~n245 & n345;
  assign n347 = ~n236 & n346;
  assign n348 = ~n227 & n347;
  assign n349 = ~n220 & n348;
  assign n350 = ~n211 & n349;
  assign n351 = ~n203 & n350;
  assign n352 = ~n195 & n351;
  assign n353 = ~n186 & n352;
  assign n354 = ~n177 & n353;
  assign n355 = ~n170 & n354;
  assign n356 = ~n163 & n355;
  assign n357 = ~n160 & n356;
  assign n358 = ~n152 & n357;
  assign n359 = ~n143 & n358;
  assign n360 = ~n135 & n359;
  assign n361 = ~n126 & n360;
  assign n362 = ~n117 & n361;
  assign n363 = ~n108 & n362;
  assign z0 = n99 | ~n363;
  assign n365 = ~m & ~n;
  assign n366 = ~o & n365;
  assign n367 = v & n366;
  assign n368 = ~b0 & n367;
  assign n369 = ~c0 & n368;
  assign n370 = ~d0 & n369;
  assign z1 = ~e0 & n370;
  assign n372 = ~n324 & ~n331;
  assign n373 = ~n286 & n372;
  assign n374 = ~n276 & n373;
  assign n375 = ~n160 & n374;
  assign a1 = n152 | ~n375;
  assign n377 = s & t;
  assign n378 = u & n377;
  assign n379 = ~v & n378;
  assign n380 = b0 & n379;
  assign n381 = ~d0 & n380;
  assign n382 = e0 & n381;
  assign n383 = ~b0 & n379;
  assign n384 = c0 & n383;
  assign n385 = d0 & n384;
  assign n386 = e0 & n385;
  assign n387 = e & s;
  assign n388 = t & n387;
  assign n389 = u & n388;
  assign n390 = ~v & n389;
  assign n391 = ~b0 & n390;
  assign n392 = c0 & n391;
  assign n393 = d0 & n392;
  assign n394 = ~e0 & n393;
  assign n395 = f & s;
  assign n396 = t & n395;
  assign n397 = u & n396;
  assign n398 = ~v & n397;
  assign n399 = ~b0 & n398;
  assign n400 = ~c0 & n399;
  assign n401 = d0 & n400;
  assign n402 = e0 & n401;
  assign n403 = ~n394 & ~n402;
  assign n404 = ~n386 & n403;
  assign n405 = ~n99 & n404;
  assign a2 = n382 | ~n405;
  assign n407 = ~n317 & n336;
  assign n408 = ~i2 & n407;
  assign n409 = ~n295 & n408;
  assign n410 = ~n286 & n409;
  assign n411 = ~n265 & n410;
  assign n412 = ~n245 & n411;
  assign n413 = ~n220 & n412;
  assign n414 = ~n203 & n413;
  assign n415 = ~n170 & n414;
  assign n416 = ~n163 & n415;
  assign n417 = ~n152 & n416;
  assign n418 = ~n126 & n417;
  assign b1 = n108 | ~n418;
  assign n420 = ~j & ~s;
  assign n421 = ~t & n420;
  assign n422 = ~u & n421;
  assign n423 = v & n422;
  assign n424 = w & n423;
  assign n425 = ~c0 & n424;
  assign n426 = d0 & n425;
  assign n427 = ~e0 & n426;
  assign n428 = ~m0 & n427;
  assign n429 = ~n0 & n428;
  assign n430 = ~o0 & n429;
  assign n431 = ~p0 & n430;
  assign n432 = ~q0 & n431;
  assign n433 = r0 & n432;
  assign n434 = ~s0 & n433;
  assign n435 = ~r0 & n432;
  assign n436 = s0 & n435;
  assign n437 = o0 & n429;
  assign n438 = ~p0 & n437;
  assign n439 = ~q0 & n438;
  assign n440 = ~s & ~t;
  assign n441 = ~u & n440;
  assign n442 = v & n441;
  assign n443 = w & n442;
  assign n444 = ~c0 & n443;
  assign n445 = d0 & n444;
  assign n446 = e0 & n445;
  assign n447 = n0 & n428;
  assign n448 = ~p0 & n447;
  assign n449 = ~q0 & n448;
  assign n450 = ~p0 & n429;
  assign n451 = q0 & n450;
  assign n452 = p0 & n428;
  assign n453 = m0 & n427;
  assign n454 = j & ~s;
  assign n455 = ~t & n454;
  assign n456 = ~u & n455;
  assign n457 = v & n456;
  assign n458 = w & n457;
  assign n459 = ~c0 & n458;
  assign n460 = ~d0 & n459;
  assign n461 = e0 & n460;
  assign n462 = ~f0 & n461;
  assign n463 = ~h0 & n462;
  assign n464 = n0 & n463;
  assign n465 = ~n0 & n463;
  assign n466 = f0 & n461;
  assign n467 = h0 & n461;
  assign n468 = ~d0 & n384;
  assign n469 = e0 & n468;
  assign n470 = ~e0 & n468;
  assign n471 = ~u & n377;
  assign n472 = ~v & n471;
  assign n473 = a0 & n472;
  assign n474 = c0 & n473;
  assign n475 = ~d0 & n474;
  assign n476 = ~e0 & n475;
  assign n477 = ~c0 & n473;
  assign n478 = d0 & n477;
  assign n479 = e0 & n478;
  assign n480 = r & s;
  assign n481 = ~t & n480;
  assign n482 = u & n481;
  assign n483 = ~v & n482;
  assign n484 = a0 & n483;
  assign n485 = c0 & n484;
  assign n486 = ~d0 & n485;
  assign n487 = ~e0 & n486;
  assign n488 = ~c0 & n484;
  assign n489 = d0 & n488;
  assign n490 = ~e0 & n489;
  assign n491 = ~c & ~d;
  assign n492 = ~s & n491;
  assign n493 = t & n492;
  assign n494 = u & n493;
  assign n495 = ~v & n494;
  assign n496 = w & n495;
  assign n497 = c0 & n496;
  assign n498 = ~d0 & n497;
  assign n499 = e0 & n498;
  assign n500 = d & ~s;
  assign n501 = t & n500;
  assign n502 = u & n501;
  assign n503 = ~v & n502;
  assign n504 = w & n503;
  assign n505 = c0 & n504;
  assign n506 = ~d0 & n505;
  assign n507 = e0 & n506;
  assign n508 = ~s & t;
  assign n509 = u & n508;
  assign n510 = ~v & n509;
  assign n511 = w & n510;
  assign n512 = c0 & n511;
  assign n513 = ~d0 & n512;
  assign n514 = ~e0 & n513;
  assign n515 = ~c0 & n511;
  assign n516 = d0 & n515;
  assign n517 = e0 & n516;
  assign n518 = u & n440;
  assign n519 = ~v & n518;
  assign n520 = c0 & n519;
  assign n521 = ~d0 & n520;
  assign n522 = ~e0 & n521;
  assign n523 = ~c0 & n519;
  assign n524 = d0 & n523;
  assign n525 = e0 & n524;
  assign n526 = ~v & n441;
  assign n527 = c0 & n526;
  assign n528 = ~d0 & n527;
  assign n529 = ~e0 & n528;
  assign n530 = ~c0 & n526;
  assign n531 = d0 & n530;
  assign n532 = e0 & n531;
  assign n533 = ~l & s;
  assign n534 = ~t & n533;
  assign n535 = u & n534;
  assign n536 = v & n535;
  assign n537 = a0 & n536;
  assign n538 = ~c0 & n537;
  assign n539 = d0 & n538;
  assign n540 = e0 & n539;
  assign n541 = z & n536;
  assign n542 = ~c0 & n541;
  assign n543 = d0 & n542;
  assign n544 = e0 & n543;
  assign n545 = s & ~t;
  assign n546 = u & n545;
  assign n547 = v & n546;
  assign n548 = w & n547;
  assign n549 = ~c0 & n548;
  assign n550 = d0 & n549;
  assign n551 = e0 & n550;
  assign n552 = ~u & n545;
  assign n553 = v & n552;
  assign n554 = c0 & n553;
  assign n555 = ~d0 & n554;
  assign n556 = ~e0 & n555;
  assign n557 = ~c0 & n553;
  assign n558 = d0 & n557;
  assign n559 = e0 & n558;
  assign n560 = v & n509;
  assign n561 = w & n560;
  assign n562 = ~c0 & n561;
  assign n563 = d0 & n562;
  assign n564 = e0 & n563;
  assign n565 = v & n508;
  assign n566 = c0 & n565;
  assign n567 = d0 & n566;
  assign n568 = ~e0 & n567;
  assign n569 = v & n197;
  assign n570 = c0 & n569;
  assign n571 = ~d0 & n570;
  assign n572 = e0 & n571;
  assign n573 = a0 & n565;
  assign n574 = ~c0 & n573;
  assign n575 = ~d0 & n574;
  assign n576 = e0 & n575;
  assign n577 = k & ~s;
  assign n578 = t & n577;
  assign n579 = v & n578;
  assign n580 = z & n579;
  assign n581 = ~c0 & n580;
  assign n582 = ~d0 & n581;
  assign n583 = e0 & n582;
  assign n584 = y & n565;
  assign n585 = ~c0 & n584;
  assign n586 = ~d0 & n585;
  assign n587 = e0 & n586;
  assign n588 = ~n583 & ~n587;
  assign n589 = ~n576 & n588;
  assign n590 = ~n572 & n589;
  assign n591 = ~n568 & n590;
  assign n592 = ~n564 & n591;
  assign n593 = ~n559 & n592;
  assign n594 = ~n556 & n593;
  assign n595 = ~n551 & n594;
  assign n596 = ~n544 & n595;
  assign n597 = ~n540 & n596;
  assign n598 = ~n532 & n597;
  assign n599 = ~n529 & n598;
  assign n600 = ~n236 & n599;
  assign n601 = ~n525 & n600;
  assign n602 = ~n522 & n601;
  assign n603 = ~n220 & n602;
  assign n604 = ~n517 & n603;
  assign n605 = ~n514 & n604;
  assign n606 = ~n507 & n605;
  assign n607 = ~n203 & n606;
  assign n608 = ~n499 & n607;
  assign n609 = ~n490 & n608;
  assign n610 = ~n487 & n609;
  assign n611 = ~n177 & n610;
  assign n612 = ~n170 & n611;
  assign n613 = ~n479 & n612;
  assign n614 = ~n476 & n613;
  assign n615 = ~n135 & n614;
  assign n616 = ~n126 & n615;
  assign n617 = ~n117 & n616;
  assign n618 = ~n470 & n617;
  assign n619 = ~n469 & n618;
  assign n620 = ~n108 & n619;
  assign n621 = ~n467 & n620;
  assign n622 = ~n466 & n621;
  assign n623 = ~n465 & n622;
  assign n624 = ~n464 & n623;
  assign n625 = ~n453 & n624;
  assign n626 = ~n452 & n625;
  assign n627 = ~n451 & n626;
  assign n628 = ~n449 & n627;
  assign n629 = ~n446 & n628;
  assign n630 = ~n439 & n629;
  assign n631 = ~n436 & n630;
  assign b2 = n434 | ~n631;
  assign n633 = ~n227 & ~n236;
  assign c1 = n99 | ~n633;
  assign n635 = x & n442;
  assign n636 = ~d0 & n635;
  assign n637 = e0 & n636;
  assign n638 = q0 & n448;
  assign n639 = ~d0 & n425;
  assign n640 = e0 & n639;
  assign n641 = ~d & s;
  assign n642 = t & n641;
  assign n643 = u & n642;
  assign n644 = ~v & n643;
  assign n645 = b0 & n644;
  assign n646 = ~d0 & n645;
  assign n647 = ~e0 & n646;
  assign n648 = ~c0 & n383;
  assign n649 = d0 & n648;
  assign n650 = ~e0 & n649;
  assign n651 = ~d0 & n648;
  assign n652 = e0 & n651;
  assign n653 = ~d0 & n477;
  assign n654 = e0 & n653;
  assign n655 = k & s;
  assign n656 = t & n655;
  assign n657 = ~u & n656;
  assign n658 = ~v & n657;
  assign n659 = z & n658;
  assign n660 = ~d0 & n659;
  assign n661 = e0 & n660;
  assign n662 = w & n472;
  assign n663 = ~d0 & n662;
  assign n664 = e0 & n663;
  assign n665 = ~r & s;
  assign n666 = ~t & n665;
  assign n667 = u & n666;
  assign n668 = ~v & n667;
  assign n669 = a0 & n668;
  assign n670 = ~c0 & n669;
  assign n671 = ~d0 & n670;
  assign n672 = e0 & n671;
  assign n673 = ~d0 & n488;
  assign n674 = e0 & n673;
  assign n675 = d0 & n512;
  assign n676 = e0 & n675;
  assign n677 = ~d0 & n515;
  assign n678 = e0 & n677;
  assign n679 = ~u & n508;
  assign n680 = ~v & n679;
  assign n681 = x & n680;
  assign n682 = ~d0 & n681;
  assign n683 = e0 & n682;
  assign n684 = w & n680;
  assign n685 = ~d0 & n684;
  assign n686 = e0 & n685;
  assign n687 = ~g & n491;
  assign n688 = ~s & n687;
  assign n689 = ~t & n688;
  assign n690 = u & n689;
  assign n691 = ~v & n690;
  assign n692 = c0 & n691;
  assign n693 = ~d0 & n692;
  assign n694 = e0 & n693;
  assign n695 = d & ~g;
  assign n696 = ~s & n695;
  assign n697 = ~t & n696;
  assign n698 = u & n697;
  assign n699 = ~v & n698;
  assign n700 = c0 & n699;
  assign n701 = ~d0 & n700;
  assign n702 = e0 & n701;
  assign n703 = x & n519;
  assign n704 = ~c0 & n703;
  assign n705 = ~d0 & n704;
  assign n706 = e0 & n705;
  assign n707 = y & n519;
  assign n708 = ~d0 & n707;
  assign n709 = e0 & n708;
  assign n710 = ~t & n492;
  assign n711 = ~u & n710;
  assign n712 = ~v & n711;
  assign n713 = c0 & n712;
  assign n714 = ~d0 & n713;
  assign n715 = e0 & n714;
  assign n716 = ~d0 & n530;
  assign n717 = e0 & n716;
  assign n718 = v & n378;
  assign n719 = d0 & n718;
  assign n720 = ~e0 & n719;
  assign n721 = u & n137;
  assign n722 = v & n721;
  assign n723 = ~d0 & n722;
  assign n724 = e0 & n723;
  assign n725 = l & s;
  assign n726 = ~t & n725;
  assign n727 = u & n726;
  assign n728 = v & n727;
  assign n729 = a0 & n728;
  assign n730 = ~c0 & n729;
  assign n731 = d0 & n730;
  assign n732 = ~e0 & n731;
  assign n733 = ~e0 & n539;
  assign n734 = z & n728;
  assign n735 = ~c0 & n734;
  assign n736 = d0 & n735;
  assign n737 = ~e0 & n736;
  assign n738 = ~e0 & n543;
  assign n739 = ~e0 & n550;
  assign n740 = ~e0 & n558;
  assign n741 = ~t & n136;
  assign n742 = ~u & n741;
  assign n743 = v & n742;
  assign n744 = ~c0 & n743;
  assign n745 = ~d0 & n744;
  assign n746 = e0 & n745;
  assign n747 = ~e0 & n563;
  assign n748 = b & ~s;
  assign n749 = t & n748;
  assign n750 = ~u & n749;
  assign n751 = v & n750;
  assign n752 = x & n751;
  assign n753 = ~c0 & n752;
  assign n754 = ~d0 & n753;
  assign n755 = e0 & n754;
  assign n756 = w & n751;
  assign n757 = ~c0 & n756;
  assign n758 = ~d0 & n757;
  assign n759 = e0 & n758;
  assign n760 = v & n518;
  assign n761 = y & n760;
  assign n762 = d0 & n761;
  assign n763 = ~e0 & n762;
  assign n764 = y & n332;
  assign n765 = ~d0 & n764;
  assign n766 = e0 & n765;
  assign n767 = a0 & n760;
  assign n768 = d0 & n767;
  assign n769 = ~e0 & n768;
  assign n770 = ~a0 & n760;
  assign n771 = d0 & n770;
  assign n772 = ~e0 & n771;
  assign n773 = ~n335 & ~n772;
  assign n774 = ~n331 & n773;
  assign n775 = ~n324 & n774;
  assign n776 = ~n317 & n775;
  assign n777 = ~n310 & n776;
  assign n778 = ~n769 & n777;
  assign n779 = ~n766 & n778;
  assign n780 = ~n763 & n779;
  assign n781 = ~n759 & n780;
  assign n782 = ~n755 & n781;
  assign n783 = ~n572 & n782;
  assign n784 = ~n568 & n783;
  assign n785 = ~i2 & n784;
  assign n786 = ~n747 & n785;
  assign n787 = ~n746 & n786;
  assign n788 = ~n740 & n787;
  assign n789 = ~n295 & n788;
  assign n790 = ~n739 & n789;
  assign n791 = ~n286 & n790;
  assign n792 = ~n738 & n791;
  assign n793 = ~n276 & n792;
  assign n794 = ~n737 & n793;
  assign n795 = ~n265 & n794;
  assign n796 = ~n733 & n795;
  assign n797 = ~n255 & n796;
  assign n798 = ~n732 & n797;
  assign n799 = ~n724 & n798;
  assign n800 = ~n720 & n799;
  assign n801 = ~n717 & n800;
  assign n802 = ~n245 & n801;
  assign n803 = ~n715 & n802;
  assign n804 = ~n236 & n803;
  assign n805 = ~n709 & n804;
  assign n806 = ~n706 & n805;
  assign n807 = ~n227 & n806;
  assign n808 = ~n702 & n807;
  assign n809 = ~n694 & n808;
  assign n810 = ~n220 & n809;
  assign n811 = ~n686 & n810;
  assign n812 = ~n683 & n811;
  assign n813 = ~n678 & n812;
  assign n814 = ~n211 & n813;
  assign n815 = ~n507 & n814;
  assign n816 = ~n203 & n815;
  assign n817 = ~n676 & n816;
  assign n818 = ~n499 & n817;
  assign n819 = ~n674 & n818;
  assign n820 = ~n672 & n819;
  assign n821 = ~n195 & n820;
  assign n822 = ~n186 & n821;
  assign n823 = ~n177 & n822;
  assign n824 = ~n170 & n823;
  assign n825 = ~n664 & n824;
  assign n826 = ~n163 & n825;
  assign n827 = ~n661 & n826;
  assign n828 = ~n160 & n827;
  assign n829 = ~n152 & n828;
  assign n830 = ~n654 & n829;
  assign n831 = ~n143 & n830;
  assign n832 = ~n135 & n831;
  assign n833 = ~n126 & n832;
  assign n834 = ~n652 & n833;
  assign n835 = ~n650 & n834;
  assign n836 = ~n402 & n835;
  assign n837 = ~n469 & n836;
  assign n838 = ~n394 & n837;
  assign n839 = ~n108 & n838;
  assign n840 = ~n647 & n839;
  assign n841 = ~n382 & n840;
  assign n842 = ~n640 & n841;
  assign n843 = ~n638 & n842;
  assign c2 = n637 | ~n843;
  assign n845 = d0 & n474;
  assign n846 = ~e0 & n845;
  assign n847 = z & n472;
  assign n848 = d0 & n847;
  assign n849 = e0 & n848;
  assign n850 = d0 & n662;
  assign n851 = e0 & n850;
  assign n852 = ~v & n546;
  assign n853 = a0 & n852;
  assign n854 = c0 & n853;
  assign n855 = d0 & n854;
  assign o1 = ~e0 & n855;
  assign n857 = d0 & n670;
  assign n1 = e0 & n857;
  assign n859 = ~v & n750;
  assign n860 = x & n859;
  assign n861 = d0 & n860;
  assign n862 = ~e0 & n861;
  assign n863 = w & n859;
  assign n864 = d0 & n863;
  assign n865 = ~e0 & n864;
  assign n866 = d0 & n520;
  assign n867 = ~e0 & n866;
  assign n868 = d0 & n527;
  assign n869 = ~e0 & n868;
  assign n870 = e0 & n731;
  assign n871 = e0 & n768;
  assign n872 = ~n769 & ~n772;
  assign n873 = ~n871 & n872;
  assign n874 = ~n763 & n873;
  assign n875 = ~n759 & n874;
  assign n876 = ~n755 & n875;
  assign n877 = ~n568 & n876;
  assign n878 = ~n747 & n877;
  assign n879 = ~n740 & n878;
  assign n880 = ~n739 & n879;
  assign n881 = ~n738 & n880;
  assign n882 = ~n737 & n881;
  assign n883 = ~n733 & n882;
  assign n884 = ~n540 & n883;
  assign n885 = ~n732 & n884;
  assign n886 = ~n870 & n885;
  assign n887 = ~n720 & n886;
  assign n888 = ~n532 & n887;
  assign n889 = ~n869 & n888;
  assign n890 = ~n525 & n889;
  assign n891 = ~n867 & n890;
  assign n892 = ~n865 & n891;
  assign n893 = ~n862 & n892;
  assign n894 = ~n517 & n893;
  assign n895 = ~n676 & n894;
  assign n896 = ~n490 & n895;
  assign n897 = ~n1 & n896;
  assign n898 = ~o1 & n897;
  assign n899 = ~n851 & n898;
  assign n900 = ~n849 & n899;
  assign n901 = ~n479 & n900;
  assign n902 = ~n846 & n901;
  assign n903 = ~n470 & n902;
  assign n904 = ~n386 & n903;
  assign n905 = ~n382 & n904;
  assign n906 = ~n640 & n905;
  assign n907 = ~n464 & n906;
  assign n908 = ~n453 & n907;
  assign n909 = ~n452 & n908;
  assign n910 = ~n451 & n909;
  assign n911 = ~n449 & n910;
  assign n912 = ~n638 & n911;
  assign n913 = ~n446 & n912;
  assign d1 = n436 | ~n913;
  assign n915 = ~i & q;
  assign n916 = s & n915;
  assign n917 = ~t & n916;
  assign n918 = u & n917;
  assign n919 = v & n918;
  assign n920 = c0 & n919;
  assign n921 = ~h & ~q;
  assign n922 = s & n921;
  assign n923 = ~t & n922;
  assign n924 = u & n923;
  assign n925 = v & n924;
  assign n926 = c0 & n925;
  assign n927 = ~f & p;
  assign n928 = s & n927;
  assign n929 = ~t & n928;
  assign n930 = u & n929;
  assign n931 = v & n930;
  assign n932 = ~c0 & n931;
  assign n933 = ~d0 & n932;
  assign n934 = e0 & n933;
  assign n935 = ~s & n921;
  assign n936 = t & n935;
  assign n937 = u & n936;
  assign n938 = v & n937;
  assign n939 = w & n938;
  assign n940 = c0 & n939;
  assign n941 = ~d0 & n940;
  assign n942 = ~e0 & n941;
  assign n943 = ~s & n915;
  assign n944 = t & n943;
  assign n945 = u & n944;
  assign n946 = v & n945;
  assign n947 = w & n946;
  assign n948 = c0 & n947;
  assign n949 = ~d0 & n948;
  assign n950 = ~e0 & n949;
  assign n951 = ~s & n927;
  assign n952 = t & n951;
  assign n953 = u & n952;
  assign n954 = v & n953;
  assign n955 = w & n954;
  assign n956 = ~c0 & n955;
  assign n957 = ~d0 & n956;
  assign n958 = e0 & n957;
  assign n959 = n & ~o;
  assign n960 = ~v & n959;
  assign n961 = ~b0 & n960;
  assign n962 = ~c0 & n961;
  assign n963 = ~d0 & n962;
  assign n964 = ~e0 & n963;
  assign n965 = ~o & s;
  assign n966 = ~t & n965;
  assign n967 = ~u & n966;
  assign n968 = ~v & n967;
  assign n969 = ~b0 & n968;
  assign n970 = ~c0 & n969;
  assign n971 = ~d0 & n970;
  assign n972 = ~e0 & n971;
  assign n973 = ~o & ~s;
  assign n974 = ~t & n973;
  assign n975 = u & n974;
  assign n976 = ~v & n975;
  assign n977 = ~x & n976;
  assign n978 = ~b0 & n977;
  assign n979 = ~c0 & n978;
  assign n980 = ~d0 & n979;
  assign n981 = ~e0 & n980;
  assign n982 = ~n972 & ~n981;
  assign n983 = ~n964 & n982;
  assign n984 = ~z1 & n983;
  assign n985 = ~n772 & n984;
  assign n986 = ~n769 & n985;
  assign n987 = ~n763 & n986;
  assign n988 = ~n587 & n987;
  assign n989 = ~n583 & n988;
  assign n990 = ~n576 & n989;
  assign n991 = ~n568 & n990;
  assign n992 = ~n958 & n991;
  assign n993 = ~n747 & n992;
  assign n994 = ~n950 & n993;
  assign n995 = ~n942 & n994;
  assign n996 = ~n740 & n995;
  assign n997 = ~n556 & n996;
  assign n998 = ~n739 & n997;
  assign n999 = ~n934 & n998;
  assign n1000 = ~n926 & n999;
  assign n1001 = ~n920 & n1000;
  assign n1002 = ~n738 & n1001;
  assign n1003 = ~n544 & n1002;
  assign n1004 = ~n737 & n1003;
  assign n1005 = ~n733 & n1004;
  assign n1006 = ~n732 & n1005;
  assign n1007 = ~n720 & n1006;
  assign n1008 = ~n245 & n1007;
  assign n1009 = ~n529 & n1008;
  assign n1010 = ~n227 & n1009;
  assign n1011 = ~n522 & n1010;
  assign n1012 = ~n211 & n1011;
  assign n1013 = ~n514 & n1012;
  assign n1014 = ~n203 & n1013;
  assign n1015 = ~n195 & n1014;
  assign n1016 = ~n186 & n1015;
  assign n1017 = ~n487 & n1016;
  assign n1018 = ~n163 & n1017;
  assign n1019 = ~n160 & n1018;
  assign n1020 = ~n152 & n1019;
  assign n1021 = ~n143 & n1020;
  assign n1022 = ~n476 & n1021;
  assign n1023 = ~n650 & n1022;
  assign n1024 = ~n470 & n1023;
  assign n1025 = ~n108 & n1024;
  assign n1026 = ~n647 & n1025;
  assign n1027 = ~n99 & n1026;
  assign n1028 = ~n467 & n1027;
  assign n1029 = ~n638 & n1028;
  assign d2 = n439 | ~n1029;
  assign n1031 = e0 & n736;
  assign n1032 = e0 & n567;
  assign n1033 = v & n679;
  assign n1034 = x & n1033;
  assign n1035 = ~c0 & n1034;
  assign n1036 = d0 & n1035;
  assign n1037 = ~e0 & n1036;
  assign n1038 = w & n1033;
  assign n1039 = ~c0 & n1038;
  assign n1040 = d0 & n1039;
  assign n1041 = ~e0 & n1040;
  assign n1042 = e0 & n762;
  assign n1043 = e0 & n771;
  assign n1044 = ~n772 & ~n1043;
  assign n1045 = ~n769 & n1044;
  assign n1046 = ~n871 & n1045;
  assign n1047 = ~n763 & n1046;
  assign n1048 = ~n1042 & n1047;
  assign n1049 = ~n759 & n1048;
  assign n1050 = ~n755 & n1049;
  assign n1051 = ~n1041 & n1050;
  assign n1052 = ~n1037 & n1051;
  assign n1053 = ~n568 & n1052;
  assign n1054 = ~n1032 & n1053;
  assign n1055 = ~n747 & n1054;
  assign n1056 = ~n564 & n1055;
  assign n1057 = ~n740 & n1056;
  assign n1058 = ~n559 & n1057;
  assign n1059 = ~n739 & n1058;
  assign n1060 = ~n551 & n1059;
  assign n1061 = ~n738 & n1060;
  assign n1062 = ~n544 & n1061;
  assign n1063 = ~n1031 & n1062;
  assign n1064 = ~n733 & n1063;
  assign n1065 = ~n540 & n1064;
  assign n1066 = ~n732 & n1065;
  assign n1067 = ~n870 & n1066;
  assign n1068 = ~n720 & n1067;
  assign n1069 = ~n532 & n1068;
  assign n1070 = ~n869 & n1069;
  assign n1071 = ~n525 & n1070;
  assign n1072 = ~n867 & n1071;
  assign n1073 = ~n517 & n1072;
  assign n1074 = ~n490 & n1073;
  assign n1075 = ~n487 & n1074;
  assign n1076 = ~n479 & n1075;
  assign n1077 = ~n476 & n1076;
  assign n1078 = ~n470 & n1077;
  assign n1079 = ~n647 & n1078;
  assign n1080 = ~n382 & n1079;
  assign e1 = n434 | ~n1080;
  assign n1082 = d0 & n635;
  assign n1083 = ~e0 & n1082;
  assign n1084 = ~f0 & n1083;
  assign n1085 = ~g0 & n1084;
  assign n1086 = ~h0 & n1085;
  assign n1087 = ~i0 & n1086;
  assign n1088 = ~j0 & n1087;
  assign n1089 = ~k0 & n1088;
  assign n1090 = ~l0 & n1089;
  assign n1091 = l0 & n1089;
  assign n1092 = k0 & n1088;
  assign n1093 = j0 & n1087;
  assign n1094 = i0 & n1086;
  assign n1095 = h0 & n1085;
  assign n1096 = g0 & n1084;
  assign n1097 = f0 & n1083;
  assign n1098 = ~s0 & n435;
  assign n1099 = c0 & n443;
  assign n1100 = e0 & n1099;
  assign n1101 = ~c0 & n380;
  assign n1102 = d0 & n1101;
  assign n1103 = ~e0 & n1102;
  assign n1104 = ~k & s;
  assign n1105 = t & n1104;
  assign n1106 = ~u & n1105;
  assign n1107 = ~v & n1106;
  assign n1108 = z & n1107;
  assign n1109 = ~d0 & n1108;
  assign n1110 = e0 & n1109;
  assign n1111 = x & n852;
  assign n1112 = e0 & n1111;
  assign n1113 = w & n852;
  assign n1114 = e0 & n1113;
  assign n1115 = ~t & n1104;
  assign n1116 = ~u & n1115;
  assign n1117 = ~v & n1116;
  assign n1118 = z & n1117;
  assign n1119 = e0 & n1118;
  assign n1120 = ~t & n655;
  assign n1121 = ~u & n1120;
  assign n1122 = ~v & n1121;
  assign n1123 = z & n1122;
  assign n1124 = e0 & n1123;
  assign n1125 = ~v & n552;
  assign n1126 = w & n1125;
  assign n1127 = e0 & n1126;
  assign n1128 = c & ~d;
  assign n1129 = ~s & n1128;
  assign n1130 = t & n1129;
  assign n1131 = u & n1130;
  assign n1132 = ~v & n1131;
  assign n1133 = w & n1132;
  assign n1134 = c0 & n1133;
  assign n1135 = ~d0 & n1134;
  assign n1136 = e0 & n1135;
  assign n1137 = f & ~s;
  assign n1138 = t & n1137;
  assign n1139 = u & n1138;
  assign n1140 = ~v & n1139;
  assign n1141 = w & n1140;
  assign n1142 = ~c0 & n1141;
  assign n1143 = d0 & n1142;
  assign n1144 = ~e0 & n1143;
  assign n1145 = a0 & n510;
  assign n1146 = ~c0 & n1145;
  assign n1147 = ~d0 & n1146;
  assign n1148 = e0 & n1147;
  assign n1149 = x & n510;
  assign n1150 = ~c0 & n1149;
  assign n1151 = ~d0 & n1150;
  assign n1152 = e0 & n1151;
  assign n1153 = g & n491;
  assign n1154 = ~s & n1153;
  assign n1155 = ~t & n1154;
  assign n1156 = u & n1155;
  assign n1157 = ~v & n1156;
  assign n1158 = c0 & n1157;
  assign n1159 = ~d0 & n1158;
  assign n1160 = e0 & n1159;
  assign n1161 = d & g;
  assign n1162 = ~s & n1161;
  assign n1163 = ~t & n1162;
  assign n1164 = u & n1163;
  assign n1165 = ~v & n1164;
  assign n1166 = c0 & n1165;
  assign n1167 = ~d0 & n1166;
  assign n1168 = e0 & n1167;
  assign n1169 = a0 & n519;
  assign n1170 = ~d0 & n1169;
  assign n1171 = e0 & n1170;
  assign n1172 = d0 & n707;
  assign n1173 = ~e0 & n1172;
  assign n1174 = w & n519;
  assign n1175 = ~d0 & n1174;
  assign l2 = e0 & n1175;
  assign n1177 = ~d & f;
  assign n1178 = ~s & n1177;
  assign n1179 = ~t & n1178;
  assign n1180 = ~u & n1179;
  assign n1181 = ~v & n1180;
  assign n1182 = ~c0 & n1181;
  assign n1183 = d0 & n1182;
  assign n1184 = ~e0 & n1183;
  assign n1185 = ~t & n500;
  assign n1186 = ~u & n1185;
  assign n1187 = ~v & n1186;
  assign n1188 = ~c0 & n1187;
  assign n1189 = d0 & n1188;
  assign n1190 = ~e0 & n1189;
  assign n1191 = e0 & n719;
  assign n1192 = w & n718;
  assign n1193 = e0 & n1192;
  assign n1194 = v & n1106;
  assign n1195 = z & n1194;
  assign n1196 = e0 & n1195;
  assign n1197 = v & n471;
  assign n1198 = a0 & n1197;
  assign n1199 = e0 & n1198;
  assign n1200 = v & n657;
  assign n1201 = z & n1200;
  assign n1202 = e0 & n1201;
  assign n1203 = w & n1197;
  assign n1204 = e0 & n1203;
  assign n1205 = h & ~q;
  assign n1206 = s & n1205;
  assign n1207 = ~t & n1206;
  assign n1208 = u & n1207;
  assign n1209 = v & n1208;
  assign n1210 = c0 & n1209;
  assign n1211 = i & q;
  assign n1212 = s & n1211;
  assign n1213 = ~t & n1212;
  assign n1214 = u & n1213;
  assign n1215 = v & n1214;
  assign n1216 = c0 & n1215;
  assign n1217 = ~k & n109;
  assign n1218 = ~p & n1217;
  assign n1219 = s & n1218;
  assign n1220 = ~t & n1219;
  assign n1221 = u & n1220;
  assign n1222 = v & n1221;
  assign n1223 = z & n1222;
  assign n1224 = ~c0 & n1223;
  assign n1225 = ~d0 & n1224;
  assign n1226 = e0 & n1225;
  assign n1227 = f & ~k;
  assign n1228 = s & n1227;
  assign n1229 = ~t & n1228;
  assign n1230 = u & n1229;
  assign n1231 = v & n1230;
  assign n1232 = z & n1231;
  assign n1233 = ~c0 & n1232;
  assign n1234 = ~d0 & n1233;
  assign n1235 = e0 & n1234;
  assign n1236 = f & k;
  assign n1237 = s & n1236;
  assign n1238 = ~t & n1237;
  assign n1239 = u & n1238;
  assign n1240 = v & n1239;
  assign n1241 = z & n1240;
  assign n1242 = ~c0 & n1241;
  assign n1243 = ~d0 & n1242;
  assign n1244 = e0 & n1243;
  assign n1245 = ~t & n395;
  assign n1246 = u & n1245;
  assign n1247 = v & n1246;
  assign n1248 = ~z & n1247;
  assign n1249 = ~c0 & n1248;
  assign n1250 = ~d0 & n1249;
  assign n1251 = e0 & n1250;
  assign n1252 = e0 & n555;
  assign n1253 = ~s & n1205;
  assign n1254 = t & n1253;
  assign n1255 = u & n1254;
  assign n1256 = v & n1255;
  assign n1257 = w & n1256;
  assign n1258 = c0 & n1257;
  assign n1259 = ~d0 & n1258;
  assign n1260 = ~e0 & n1259;
  assign n1261 = ~s & n1211;
  assign n1262 = t & n1261;
  assign n1263 = u & n1262;
  assign n1264 = v & n1263;
  assign n1265 = w & n1264;
  assign n1266 = c0 & n1265;
  assign n1267 = ~d0 & n1266;
  assign n1268 = ~e0 & n1267;
  assign n1269 = v & n1139;
  assign n1270 = w & n1269;
  assign n1271 = ~c0 & n1270;
  assign n1272 = ~d0 & n1271;
  assign n1273 = e0 & n1272;
  assign n1274 = ~k & ~s;
  assign n1275 = t & n1274;
  assign n1276 = v & n1275;
  assign n1277 = z & n1276;
  assign n1278 = ~c0 & n1277;
  assign n1279 = ~d0 & n1278;
  assign n1280 = e0 & n1279;
  assign n1281 = ~t & n1274;
  assign n1282 = u & n1281;
  assign n1283 = v & n1282;
  assign n1284 = z & n1283;
  assign n1285 = o & ~b0;
  assign n1286 = ~c0 & n1285;
  assign n1287 = ~d0 & n1286;
  assign n1288 = ~e0 & n1287;
  assign n1289 = a0 & n718;
  assign n1290 = e0 & n1289;
  assign n1291 = ~n981 & ~n1288;
  assign n1292 = ~n972 & n1291;
  assign n1293 = ~n964 & n1292;
  assign n1294 = ~z1 & n1293;
  assign n1295 = ~n335 & n1294;
  assign n1296 = ~n772 & n1295;
  assign n1297 = ~n1043 & n1296;
  assign n1298 = ~n1284 & n1297;
  assign n1299 = ~n331 & n1298;
  assign n1300 = ~n324 & n1299;
  assign n1301 = ~n317 & n1300;
  assign n1302 = ~n310 & n1301;
  assign n1303 = ~n769 & n1302;
  assign n1304 = ~n871 & n1303;
  assign n1305 = ~n766 & n1304;
  assign n1306 = ~n763 & n1305;
  assign n1307 = ~n1042 & n1306;
  assign n1308 = ~n587 & n1307;
  assign n1309 = ~n583 & n1308;
  assign n1310 = ~n576 & n1309;
  assign n1311 = ~n759 & n1310;
  assign n1312 = ~n755 & n1311;
  assign n1313 = ~n1280 & n1312;
  assign n1314 = ~n1041 & n1313;
  assign n1315 = ~n1037 & n1314;
  assign n1316 = ~n572 & n1315;
  assign n1317 = ~n568 & n1316;
  assign n1318 = ~n1032 & n1317;
  assign n1319 = ~n1273 & n1318;
  assign n1320 = ~n958 & n1319;
  assign n1321 = ~i2 & n1320;
  assign n1322 = ~n747 & n1321;
  assign n1323 = ~n564 & n1322;
  assign n1324 = ~n950 & n1323;
  assign n1325 = ~n1268 & n1324;
  assign n1326 = ~n942 & n1325;
  assign n1327 = ~n1260 & n1326;
  assign n1328 = ~n746 & n1327;
  assign n1329 = ~n740 & n1328;
  assign n1330 = ~n559 & n1329;
  assign n1331 = ~n556 & n1330;
  assign n1332 = ~n1252 & n1331;
  assign n1333 = ~n295 & n1332;
  assign n1334 = ~n739 & n1333;
  assign n1335 = ~n551 & n1334;
  assign n1336 = ~n934 & n1335;
  assign n1337 = ~n926 & n1336;
  assign n1338 = ~n1251 & n1337;
  assign n1339 = ~n1244 & n1338;
  assign n1340 = ~n1235 & n1339;
  assign n1341 = ~n1226 & n1340;
  assign n1342 = ~n1216 & n1341;
  assign n1343 = ~n1210 & n1342;
  assign n1344 = ~n920 & n1343;
  assign n1345 = ~n286 & n1344;
  assign n1346 = ~n738 & n1345;
  assign n1347 = ~n544 & n1346;
  assign n1348 = ~n276 & n1347;
  assign n1349 = ~n737 & n1348;
  assign n1350 = ~n1031 & n1349;
  assign n1351 = ~n265 & n1350;
  assign n1352 = ~n733 & n1351;
  assign n1353 = ~n540 & n1352;
  assign n1354 = ~n255 & n1353;
  assign n1355 = ~n732 & n1354;
  assign n1356 = ~n870 & n1355;
  assign n1357 = ~n1204 & n1356;
  assign n1358 = ~n1202 & n1357;
  assign n1359 = ~n1199 & n1358;
  assign n1360 = ~n1196 & n1359;
  assign n1361 = ~n1193 & n1360;
  assign n1362 = ~n724 & n1361;
  assign n1363 = ~n720 & n1362;
  assign n1364 = ~n1191 & n1363;
  assign n1365 = ~n717 & n1364;
  assign n1366 = ~n1190 & n1365;
  assign n1367 = ~n1184 & n1366;
  assign n1368 = ~n245 & n1367;
  assign n1369 = ~n532 & n1368;
  assign n1370 = ~n529 & n1369;
  assign n1371 = ~n715 & n1370;
  assign n1372 = ~n236 & n1371;
  assign n1373 = ~n869 & n1372;
  assign n1374 = ~l2 & n1373;
  assign n1375 = ~n709 & n1374;
  assign n1376 = ~n1173 & n1375;
  assign n1377 = ~n1171 & n1376;
  assign n1378 = ~n706 & n1377;
  assign n1379 = ~n227 & n1378;
  assign n1380 = ~n525 & n1379;
  assign n1381 = ~n522 & n1380;
  assign n1382 = ~n702 & n1381;
  assign n1383 = ~n694 & n1382;
  assign n1384 = ~n1168 & n1383;
  assign n1385 = ~n1160 & n1384;
  assign n1386 = ~n220 & n1385;
  assign n1387 = ~n867 & n1386;
  assign n1388 = ~n686 & n1387;
  assign n1389 = ~n865 & n1388;
  assign n1390 = ~n683 & n1389;
  assign n1391 = ~n862 & n1390;
  assign n1392 = ~n678 & n1391;
  assign n1393 = ~n1152 & n1392;
  assign n1394 = ~n1148 & n1393;
  assign n1395 = ~n1144 & n1394;
  assign n1396 = ~n211 & n1395;
  assign n1397 = ~n517 & n1396;
  assign n1398 = ~n514 & n1397;
  assign n1399 = ~n507 & n1398;
  assign n1400 = ~n203 & n1399;
  assign n1401 = ~n676 & n1400;
  assign n1402 = ~n499 & n1401;
  assign n1403 = ~n1136 & n1402;
  assign n1404 = ~n1127 & n1403;
  assign n1405 = ~n1124 & n1404;
  assign n1406 = ~n1119 & n1405;
  assign n1407 = ~n1114 & n1406;
  assign n1408 = ~n1112 & n1407;
  assign n1409 = ~n674 & n1408;
  assign n1410 = ~n672 & n1409;
  assign n1411 = ~n195 & n1410;
  assign n1412 = ~n490 & n1411;
  assign n1413 = ~n186 & n1412;
  assign n1414 = ~n487 & n1413;
  assign n1415 = ~n1 & n1414;
  assign n1416 = ~n177 & n1415;
  assign n1417 = ~n170 & n1416;
  assign n1418 = ~o1 & n1417;
  assign n1419 = ~n664 & n1418;
  assign n1420 = ~n163 & n1419;
  assign n1421 = ~n851 & n1420;
  assign n1422 = ~n1110 & n1421;
  assign n1423 = ~n661 & n1422;
  assign n1424 = ~n160 & n1423;
  assign n1425 = ~n152 & n1424;
  assign n1426 = ~n849 & n1425;
  assign n1427 = ~n654 & n1426;
  assign n1428 = ~n143 & n1427;
  assign n1429 = ~n479 & n1428;
  assign n1430 = ~n476 & n1429;
  assign n1431 = ~n135 & n1430;
  assign n1432 = ~n126 & n1431;
  assign n1433 = ~n846 & n1432;
  assign n1434 = ~n652 & n1433;
  assign n1435 = ~n650 & n1434;
  assign n1436 = ~n402 & n1435;
  assign n1437 = ~n117 & n1436;
  assign n1438 = ~n470 & n1437;
  assign n1439 = ~n469 & n1438;
  assign n1440 = ~n394 & n1439;
  assign n1441 = ~n108 & n1440;
  assign n1442 = ~n386 & n1441;
  assign n1443 = ~n647 & n1442;
  assign n1444 = ~n99 & n1443;
  assign n1445 = ~n382 & n1444;
  assign n1446 = ~n1103 & n1445;
  assign n1447 = ~n640 & n1446;
  assign n1448 = ~n467 & n1447;
  assign n1449 = ~n466 & n1448;
  assign n1450 = ~n465 & n1449;
  assign n1451 = ~n464 & n1450;
  assign n1452 = ~n453 & n1451;
  assign n1453 = ~n452 & n1452;
  assign n1454 = ~n451 & n1453;
  assign n1455 = ~n449 & n1454;
  assign n1456 = ~n638 & n1455;
  assign n1457 = ~n446 & n1456;
  assign n1458 = ~n1100 & n1457;
  assign n1459 = ~n439 & n1458;
  assign n1460 = ~n436 & n1459;
  assign n1461 = ~n1098 & n1460;
  assign n1462 = ~n434 & n1461;
  assign n1463 = ~n637 & n1462;
  assign n1464 = ~n1097 & n1463;
  assign n1465 = ~n1096 & n1464;
  assign n1466 = ~n1095 & n1465;
  assign n1467 = ~n1094 & n1466;
  assign n1468 = ~n1093 & n1467;
  assign n1469 = ~n1092 & n1468;
  assign n1470 = ~n1091 & n1469;
  assign n1471 = ~n1090 & n1470;
  assign e2 = n1290 | ~n1471;
  assign n1473 = ~n1041 & n1048;
  assign n1474 = ~n1037 & n1473;
  assign n1475 = ~n568 & n1474;
  assign n1476 = ~n1032 & n1475;
  assign n1477 = ~n747 & n1476;
  assign n1478 = ~n564 & n1477;
  assign n1479 = ~n740 & n1478;
  assign n1480 = ~n559 & n1479;
  assign n1481 = ~n739 & n1480;
  assign n1482 = ~n551 & n1481;
  assign n1483 = ~n738 & n1482;
  assign n1484 = ~n544 & n1483;
  assign n1485 = ~n737 & n1484;
  assign n1486 = ~n1031 & n1485;
  assign n1487 = ~n733 & n1486;
  assign n1488 = ~n540 & n1487;
  assign n1489 = ~n732 & n1488;
  assign n1490 = ~n870 & n1489;
  assign n1491 = ~n1202 & n1490;
  assign n1492 = ~n1199 & n1491;
  assign n1493 = ~n720 & n1492;
  assign n1494 = ~n1191 & n1493;
  assign n1495 = ~n532 & n1494;
  assign n1496 = ~n869 & n1495;
  assign n1497 = ~n525 & n1496;
  assign n1498 = ~n867 & n1497;
  assign n1499 = ~n865 & n1498;
  assign n1500 = ~n862 & n1499;
  assign n1501 = ~n517 & n1500;
  assign n1502 = ~n676 & n1501;
  assign n1503 = ~n490 & n1502;
  assign n1504 = ~n487 & n1503;
  assign n1505 = ~n1 & n1504;
  assign n1506 = ~o1 & n1505;
  assign n1507 = ~n851 & n1506;
  assign n1508 = ~n849 & n1507;
  assign n1509 = ~n479 & n1508;
  assign n1510 = ~n476 & n1509;
  assign n1511 = ~n846 & n1510;
  assign n1512 = ~n470 & n1511;
  assign n1513 = ~n386 & n1512;
  assign n1514 = ~n647 & n1513;
  assign n1515 = ~n382 & n1514;
  assign n1516 = ~n640 & n1515;
  assign n1517 = ~n436 & n1516;
  assign f1 = n1098 | ~n1517;
  assign n1519 = ~a & s;
  assign n1520 = t & n1519;
  assign n1521 = u & n1520;
  assign n1522 = v & n1521;
  assign n1523 = y & n1522;
  assign n1524 = ~d0 & n1523;
  assign n1525 = e0 & n1524;
  assign n1526 = ~t & n1519;
  assign n1527 = ~u & n1526;
  assign n1528 = v & n1527;
  assign n1529 = ~c0 & n1528;
  assign n1530 = ~d0 & n1529;
  assign n1531 = e0 & n1530;
  assign n1532 = ~a & ~s;
  assign n1533 = ~t & n1532;
  assign n1534 = u & n1533;
  assign n1535 = v & n1534;
  assign n1536 = y & n1535;
  assign n1537 = ~d0 & n1536;
  assign n1538 = e0 & n1537;
  assign n1539 = ~d0 & n562;
  assign n1540 = e0 & n1539;
  assign n1541 = ~a & n1540;
  assign n1542 = ~f & n1541;
  assign n1543 = ~p & n1542;
  assign n1544 = e0 & n528;
  assign n1545 = ~a & n1544;
  assign n1546 = ~d & n1545;
  assign n1547 = ~c & n1546;
  assign n1548 = e0 & n521;
  assign n1549 = ~a & n1548;
  assign n1550 = ~d & n1549;
  assign n1551 = c & n1550;
  assign n1552 = ~c0 & n547;
  assign n1553 = ~d0 & n1552;
  assign n1554 = e0 & n1553;
  assign n1555 = ~a & n1554;
  assign n1556 = ~f & n1555;
  assign n1557 = ~p & n1556;
  assign n1558 = ~c0 & n379;
  assign n1559 = d0 & n1558;
  assign n1560 = e0 & n1559;
  assign n1561 = ~a & n1560;
  assign n1562 = ~b0 & n1561;
  assign n1563 = ~f & n1562;
  assign n1564 = ~e0 & n531;
  assign n1565 = ~a & n1564;
  assign n1566 = ~d & n1565;
  assign n1567 = ~f & n1566;
  assign n1568 = ~e0 & n516;
  assign n1569 = ~a & n1568;
  assign n1570 = ~f & n1569;
  assign n1571 = c0 & n379;
  assign n1572 = d0 & n1571;
  assign n1573 = ~e0 & n1572;
  assign n1574 = ~a & n1573;
  assign n1575 = ~b0 & n1574;
  assign n1576 = ~e & n1575;
  assign n1577 = ~c0 & n852;
  assign n1578 = d0 & n1577;
  assign n1579 = ~e0 & n1578;
  assign n1580 = ~a & n1579;
  assign n1581 = a0 & n1580;
  assign n1582 = ~r & n1581;
  assign n1583 = r & n1581;
  assign n1584 = c0 & n852;
  assign n1585 = ~d0 & n1584;
  assign n1586 = e0 & n1585;
  assign n1587 = ~a & n1586;
  assign n1588 = a0 & n1587;
  assign n1589 = l & n1588;
  assign n1590 = ~e0 & n524;
  assign n1591 = ~a & n1590;
  assign n1592 = x & n1591;
  assign n1593 = ~b & ~s;
  assign n1594 = t & n1593;
  assign n1595 = ~u & n1594;
  assign n1596 = v & n1595;
  assign n1597 = ~c0 & n1596;
  assign n1598 = ~d0 & n1597;
  assign n1599 = e0 & n1598;
  assign n1600 = x & n1599;
  assign n1601 = ~c0 & n472;
  assign n1602 = d0 & n1601;
  assign n1603 = ~e0 & n1602;
  assign n1604 = ~a & n1603;
  assign n1605 = a0 & n1604;
  assign n1606 = c0 & n472;
  assign n1607 = ~d0 & n1606;
  assign n1608 = e0 & n1607;
  assign n1609 = ~a & n1608;
  assign n1610 = a0 & n1609;
  assign n1611 = ~e0 & n675;
  assign n1612 = ~a & n1611;
  assign n1613 = w & n1596;
  assign n1614 = ~c0 & n1613;
  assign n1615 = ~d0 & n1614;
  assign n1616 = e0 & n1615;
  assign n1617 = ~v & n1595;
  assign n1618 = d0 & n1617;
  assign n1619 = ~e0 & n1618;
  assign n1620 = x & n1619;
  assign n1621 = ~d0 & n379;
  assign n1622 = ~a & n1621;
  assign n1623 = d & n1622;
  assign n1624 = b0 & n1623;
  assign n1625 = d0 & n472;
  assign n1626 = ~e0 & n1625;
  assign n1627 = ~a & n1626;
  assign n1628 = z & n1627;
  assign n1629 = ~d0 & n760;
  assign n1630 = e0 & n1629;
  assign n1631 = ~a & n1630;
  assign n1632 = z & n1631;
  assign n1633 = a0 & n1631;
  assign n1634 = ~e0 & n850;
  assign n1635 = ~a & n1634;
  assign n1636 = w & n760;
  assign n1637 = ~d0 & n1636;
  assign n1638 = e0 & n1637;
  assign n1639 = ~a & n1638;
  assign n1640 = w & n1617;
  assign n1641 = d0 & n1640;
  assign n1642 = ~e0 & n1641;
  assign n1643 = ~n1531 & ~n1538;
  assign n1644 = ~n1525 & n1643;
  assign n1645 = ~d0 & n566;
  assign n1646 = e0 & n1645;
  assign n1647 = ~a & n1646;
  assign n1648 = n1644 & ~n1647;
  assign n1649 = ~n1642 & n1648;
  assign n1650 = ~n1639 & n1649;
  assign n1651 = ~n1635 & n1650;
  assign n1652 = ~n1633 & n1651;
  assign n1653 = ~n1632 & n1652;
  assign n1654 = ~n1628 & n1653;
  assign n1655 = ~n1624 & n1654;
  assign n1656 = ~n1620 & n1655;
  assign n1657 = ~n1616 & n1656;
  assign n1658 = ~n1612 & n1657;
  assign n1659 = ~n1610 & n1658;
  assign n1660 = ~n1605 & n1659;
  assign n1661 = ~n1600 & n1660;
  assign n1662 = ~n1592 & n1661;
  assign n1663 = ~n1589 & n1662;
  assign n1664 = ~n1583 & n1663;
  assign n1665 = ~n1582 & n1664;
  assign n1666 = ~n1576 & n1665;
  assign n1667 = ~n1570 & n1666;
  assign n1668 = ~n1567 & n1667;
  assign n1669 = ~n1563 & n1668;
  assign n1670 = ~n1557 & n1669;
  assign n1671 = ~n1551 & n1670;
  assign n1672 = ~n1547 & n1671;
  assign f2 = n1543 | ~n1672;
  assign n1674 = v & n959;
  assign n1675 = ~b0 & n1674;
  assign n1676 = ~c0 & n1675;
  assign n1677 = ~d0 & n1676;
  assign n1678 = ~e0 & n1677;
  assign n1679 = ~n1288 & ~n1678;
  assign n1680 = ~n759 & n1679;
  assign n1681 = ~n755 & n1680;
  assign n1682 = ~n737 & n1681;
  assign n1683 = ~n1202 & n1682;
  assign n1684 = ~n1199 & n1683;
  assign n1685 = ~n1191 & n1684;
  assign n1686 = ~n717 & n1685;
  assign n1687 = ~n706 & n1686;
  assign n1688 = ~n686 & n1687;
  assign n1689 = ~n865 & n1688;
  assign n1690 = ~n683 & n1689;
  assign n1691 = ~n862 & n1690;
  assign n1692 = ~n678 & n1691;
  assign n1693 = ~n1152 & n1692;
  assign n1694 = ~n1148 & n1693;
  assign n1695 = ~n507 & n1694;
  assign n1696 = ~n676 & n1695;
  assign n1697 = ~n499 & n1696;
  assign n1698 = ~n1114 & n1697;
  assign n1699 = ~n1112 & n1698;
  assign n1700 = ~n674 & n1699;
  assign n1701 = ~n672 & n1700;
  assign n1702 = ~n487 & n1701;
  assign n1703 = ~n1 & n1702;
  assign n1704 = ~o1 & n1703;
  assign n1705 = ~n664 & n1704;
  assign n1706 = ~n851 & n1705;
  assign n1707 = ~n661 & n1706;
  assign n1708 = ~n849 & n1707;
  assign n1709 = ~n654 & n1708;
  assign n1710 = ~n476 & n1709;
  assign n1711 = ~n846 & n1710;
  assign n1712 = ~n652 & n1711;
  assign n1713 = ~n386 & n1712;
  assign n1714 = ~n647 & n1713;
  assign n1715 = ~n464 & n1714;
  assign n1716 = ~n451 & n1715;
  assign n1717 = ~n449 & n1716;
  assign n1718 = ~n638 & n1717;
  assign n1719 = ~n446 & n1718;
  assign g1 = n436 | ~n1719;
  assign n1721 = ~n763 & n872;
  assign n1722 = ~n759 & n1721;
  assign n1723 = ~n755 & n1722;
  assign n1724 = ~n568 & n1723;
  assign n1725 = ~n747 & n1724;
  assign n1726 = ~n740 & n1725;
  assign n1727 = ~n739 & n1726;
  assign n1728 = ~n738 & n1727;
  assign n1729 = ~n737 & n1728;
  assign n1730 = ~n733 & n1729;
  assign n1731 = ~n732 & n1730;
  assign n1732 = ~n720 & n1731;
  assign n1733 = ~n869 & n1732;
  assign n1734 = ~n525 & n1733;
  assign n1735 = ~n867 & n1734;
  assign n1736 = ~n865 & n1735;
  assign n1737 = ~n862 & n1736;
  assign n1738 = ~n1144 & n1737;
  assign n1739 = ~n1136 & n1738;
  assign n1740 = ~n1 & n1739;
  assign n1741 = ~o1 & n1740;
  assign n1742 = ~n851 & n1741;
  assign n1743 = ~n849 & n1742;
  assign n1744 = ~n846 & n1743;
  assign n1745 = ~n394 & n1744;
  assign g2 = n382 | ~n1745;
  assign n1747 = ~n755 & ~n871;
  assign n1748 = ~n1032 & n1747;
  assign n1749 = ~n564 & n1748;
  assign n1750 = ~n737 & n1749;
  assign n1751 = ~n540 & n1750;
  assign n1752 = ~n870 & n1751;
  assign n1753 = ~n1199 & n1752;
  assign n1754 = ~n865 & n1753;
  assign n1755 = ~n862 & n1754;
  assign n1756 = ~n507 & n1755;
  assign n1757 = ~n676 & n1756;
  assign n1758 = ~n499 & n1757;
  assign n1759 = ~n487 & n1758;
  assign n1760 = ~n1 & n1759;
  assign n1761 = ~o1 & n1760;
  assign n1762 = ~n851 & n1761;
  assign n1763 = ~n849 & n1762;
  assign n1764 = ~n476 & n1763;
  assign n1765 = ~n846 & n1764;
  assign n1766 = ~n386 & n1765;
  assign n1767 = ~n647 & n1766;
  assign n1768 = ~n467 & n1767;
  assign n1769 = ~n464 & n1768;
  assign n1770 = ~n452 & n1769;
  assign n1771 = ~n449 & n1770;
  assign n1772 = ~n446 & n1771;
  assign h1 = n439 | ~n1772;
  assign n1774 = ~n1251 & ~n1273;
  assign n1775 = ~n1244 & n1774;
  assign n1776 = ~n1190 & n1775;
  assign n1777 = ~n1184 & n1776;
  assign n1778 = ~n1144 & n1777;
  assign h2 = n402 | ~n1778;
  assign n1780 = ~n772 & n1679;
  assign n1781 = ~n769 & n1780;
  assign n1782 = ~n763 & n1781;
  assign n1783 = ~n759 & n1782;
  assign n1784 = ~n755 & n1783;
  assign n1785 = ~n568 & n1784;
  assign n1786 = ~n747 & n1785;
  assign n1787 = ~n746 & n1786;
  assign n1788 = ~n740 & n1787;
  assign n1789 = ~n556 & n1788;
  assign n1790 = ~n739 & n1789;
  assign n1791 = ~n738 & n1790;
  assign n1792 = ~n737 & n1791;
  assign n1793 = ~n733 & n1792;
  assign n1794 = ~n732 & n1793;
  assign n1795 = ~n720 & n1794;
  assign n1796 = ~n1190 & n1795;
  assign n1797 = ~n1184 & n1796;
  assign n1798 = ~n532 & n1797;
  assign n1799 = ~n236 & n1798;
  assign n1800 = ~n869 & n1799;
  assign n1801 = ~n709 & n1800;
  assign n1802 = ~n525 & n1801;
  assign n1803 = ~n1168 & n1802;
  assign n1804 = ~n1160 & n1803;
  assign n1805 = ~n220 & n1804;
  assign n1806 = ~n867 & n1805;
  assign n1807 = ~n686 & n1806;
  assign n1808 = ~n865 & n1807;
  assign n1809 = ~n862 & n1808;
  assign n1810 = ~n1144 & n1809;
  assign n1811 = ~n517 & n1810;
  assign n1812 = ~n676 & n1811;
  assign n1813 = ~n1136 & n1812;
  assign n1814 = ~n674 & n1813;
  assign n1815 = ~n490 & n1814;
  assign n1816 = ~n1 & n1815;
  assign n1817 = ~o1 & n1816;
  assign n1818 = ~n851 & n1817;
  assign n1819 = ~n849 & n1818;
  assign n1820 = ~n654 & n1819;
  assign n1821 = ~n479 & n1820;
  assign n1822 = ~n846 & n1821;
  assign n1823 = ~n402 & n1822;
  assign n1824 = ~n470 & n1823;
  assign n1825 = ~n394 & n1824;
  assign n1826 = ~n386 & n1825;
  assign n1827 = ~n99 & n1826;
  assign n1828 = ~n382 & n1827;
  assign n1829 = ~n1103 & n1828;
  assign n1830 = ~n1100 & n1829;
  assign n1831 = ~n434 & n1830;
  assign n1832 = ~n637 & n1831;
  assign n1833 = ~n1097 & n1832;
  assign n1834 = ~n1096 & n1833;
  assign n1835 = ~n1094 & n1834;
  assign n1836 = ~n1093 & n1835;
  assign i1 = n1091 | ~n1836;
  assign n1838 = ~n769 & n1679;
  assign n1839 = ~n737 & n1838;
  assign n1840 = ~n733 & n1839;
  assign n1841 = ~n732 & n1840;
  assign n1842 = ~n1190 & n1841;
  assign n1843 = ~n1184 & n1842;
  assign n1844 = ~n236 & n1843;
  assign n1845 = ~l2 & n1844;
  assign n1846 = ~n1173 & n1845;
  assign n1847 = ~n1168 & n1846;
  assign n1848 = ~n1160 & n1847;
  assign n1849 = ~n220 & n1848;
  assign n1850 = ~n865 & n1849;
  assign n1851 = ~n862 & n1850;
  assign n1852 = ~n1152 & n1851;
  assign n1853 = ~n1148 & n1852;
  assign n1854 = ~n1144 & n1853;
  assign n1855 = ~n507 & n1854;
  assign n1856 = ~n676 & n1855;
  assign n1857 = ~n499 & n1856;
  assign n1858 = ~n1136 & n1857;
  assign n1859 = ~n1114 & n1858;
  assign n1860 = ~n674 & n1859;
  assign n1861 = ~n672 & n1860;
  assign n1862 = ~n487 & n1861;
  assign n1863 = ~n1 & n1862;
  assign n1864 = ~o1 & n1863;
  assign n1865 = ~n664 & n1864;
  assign n1866 = ~n851 & n1865;
  assign n1867 = ~n661 & n1866;
  assign n1868 = ~n849 & n1867;
  assign n1869 = ~n654 & n1868;
  assign n1870 = ~n476 & n1869;
  assign n1871 = ~n846 & n1870;
  assign n1872 = ~n652 & n1871;
  assign n1873 = ~n650 & n1872;
  assign n1874 = ~n402 & n1873;
  assign n1875 = ~n470 & n1874;
  assign n1876 = ~n394 & n1875;
  assign n1877 = ~n386 & n1876;
  assign n1878 = ~n647 & n1877;
  assign n1879 = ~n99 & n1878;
  assign n1880 = ~n1103 & n1879;
  assign n1881 = ~n640 & n1880;
  assign n1882 = ~n464 & n1881;
  assign n1883 = ~n453 & n1882;
  assign n1884 = ~n452 & n1883;
  assign n1885 = ~n451 & n1884;
  assign n1886 = ~n449 & n1885;
  assign n1887 = ~n638 & n1886;
  assign n1888 = ~n446 & n1887;
  assign j1 = n436 | ~n1888;
  assign n1890 = ~n1043 & n1780;
  assign n1891 = ~n769 & n1890;
  assign n1892 = ~n871 & n1891;
  assign n1893 = ~n763 & n1892;
  assign n1894 = ~n1042 & n1893;
  assign n1895 = ~n759 & n1894;
  assign n1896 = ~n755 & n1895;
  assign n1897 = ~n1041 & n1896;
  assign n1898 = ~n1037 & n1897;
  assign n1899 = ~n568 & n1898;
  assign n1900 = ~n1032 & n1899;
  assign n1901 = ~n747 & n1900;
  assign n1902 = ~n564 & n1901;
  assign n1903 = ~n740 & n1902;
  assign n1904 = ~n559 & n1903;
  assign n1905 = ~n1252 & n1904;
  assign n1906 = ~n739 & n1905;
  assign n1907 = ~n551 & n1906;
  assign n1908 = ~n738 & n1907;
  assign n1909 = ~n544 & n1908;
  assign n1910 = ~n737 & n1909;
  assign n1911 = ~n1031 & n1910;
  assign n1912 = ~n540 & n1911;
  assign n1913 = ~n870 & n1912;
  assign n1914 = ~n1204 & n1913;
  assign n1915 = ~n1202 & n1914;
  assign n1916 = ~n1199 & n1915;
  assign n1917 = ~n720 & n1916;
  assign n1918 = ~n1191 & n1917;
  assign n1919 = ~n532 & n1918;
  assign n1920 = ~n869 & n1919;
  assign n1921 = ~n709 & n1920;
  assign n1922 = ~n525 & n1921;
  assign n1923 = ~n867 & n1922;
  assign n1924 = ~n686 & n1923;
  assign n1925 = ~n1152 & n1924;
  assign n1926 = ~n517 & n1925;
  assign n1927 = ~n507 & n1926;
  assign n1928 = ~n676 & n1927;
  assign n1929 = ~n499 & n1928;
  assign n1930 = ~n1114 & n1929;
  assign n1931 = ~n1112 & n1930;
  assign n1932 = ~n674 & n1931;
  assign n1933 = ~n490 & n1932;
  assign n1934 = ~n487 & n1933;
  assign n1935 = ~n1 & n1934;
  assign n1936 = ~o1 & n1935;
  assign n1937 = ~n851 & n1936;
  assign n1938 = ~n849 & n1937;
  assign n1939 = ~n654 & n1938;
  assign n1940 = ~n479 & n1939;
  assign n1941 = ~n476 & n1940;
  assign n1942 = ~n846 & n1941;
  assign n1943 = ~n650 & n1942;
  assign n1944 = ~n386 & n1943;
  assign n1945 = ~n382 & n1944;
  assign n1946 = ~n1103 & n1945;
  assign n1947 = ~n467 & n1946;
  assign n1948 = ~n1100 & n1947;
  assign n1949 = ~n439 & n1948;
  assign n1950 = ~n1098 & n1949;
  assign n1951 = ~n434 & n1950;
  assign n1952 = ~n637 & n1951;
  assign n1953 = ~n1092 & n1952;
  assign k1 = n1091 | ~n1953;
  assign k2 = n709 | l2;
  assign n1956 = ~n763 & n1780;
  assign n1957 = ~n759 & n1956;
  assign n1958 = ~n755 & n1957;
  assign n1959 = ~n568 & n1958;
  assign n1960 = ~n747 & n1959;
  assign n1961 = ~n746 & n1960;
  assign n1962 = ~n740 & n1961;
  assign n1963 = ~n1252 & n1962;
  assign n1964 = ~n739 & n1963;
  assign n1965 = ~n738 & n1964;
  assign n1966 = ~n720 & n1965;
  assign n1967 = ~n717 & n1966;
  assign n1968 = ~n532 & n1967;
  assign n1969 = ~n869 & n1968;
  assign n1970 = ~n709 & n1969;
  assign n1971 = ~n706 & n1970;
  assign n1972 = ~n525 & n1971;
  assign n1973 = ~n867 & n1972;
  assign n1974 = ~n686 & n1973;
  assign n1975 = ~n865 & n1974;
  assign n1976 = ~n683 & n1975;
  assign n1977 = ~n862 & n1976;
  assign n1978 = ~n678 & n1977;
  assign n1979 = ~n1152 & n1978;
  assign n1980 = ~n1148 & n1979;
  assign n1981 = ~n517 & n1980;
  assign n1982 = ~n1124 & n1981;
  assign n1983 = ~n1114 & n1982;
  assign n1984 = ~n672 & n1983;
  assign n1985 = ~n490 & n1984;
  assign n1986 = ~n664 & n1985;
  assign n1987 = ~n661 & n1986;
  assign n1988 = ~n479 & n1987;
  assign n1989 = ~n652 & n1988;
  assign n1990 = ~n647 & n1989;
  assign n1991 = ~n382 & n1990;
  assign n1992 = ~n1103 & n1991;
  assign n1993 = ~n1094 & n1992;
  assign n1994 = ~n1093 & n1993;
  assign n1995 = ~n1092 & n1994;
  assign l1 = n1091 | ~n1995;
  assign n1997 = ~n746 & n1725;
  assign n1998 = ~n740 & n1997;
  assign n1999 = ~n739 & n1998;
  assign n2000 = ~n738 & n1999;
  assign n2001 = ~n733 & n2000;
  assign n2002 = ~n732 & n2001;
  assign n2003 = ~n720 & n2002;
  assign n2004 = ~n717 & n2003;
  assign n2005 = ~n532 & n2004;
  assign n2006 = ~n869 & n2005;
  assign n2007 = ~l2 & n2006;
  assign n2008 = ~n1173 & n2007;
  assign n2009 = ~n706 & n2008;
  assign n2010 = ~n525 & n2009;
  assign n2011 = ~n867 & n2010;
  assign n2012 = ~n686 & n2011;
  assign n2013 = ~n683 & n2012;
  assign n2014 = ~n862 & n2013;
  assign n2015 = ~n678 & n2014;
  assign n2016 = ~n1152 & n2015;
  assign n2017 = ~n517 & n2016;
  assign n2018 = ~n507 & n2017;
  assign n2019 = ~n499 & n2018;
  assign n2020 = ~n1112 & n2019;
  assign n2021 = ~n674 & n2020;
  assign n2022 = ~n672 & n2021;
  assign n2023 = ~n490 & n2022;
  assign n2024 = ~n487 & n2023;
  assign n2025 = ~n664 & n2024;
  assign n2026 = ~n661 & n2025;
  assign n2027 = ~n654 & n2026;
  assign n2028 = ~n479 & n2027;
  assign n2029 = ~n476 & n2028;
  assign n2030 = ~n652 & n2029;
  assign n2031 = ~n470 & n2030;
  assign n2032 = ~n647 & n2031;
  assign n2033 = ~n382 & n2032;
  assign n2034 = ~n1103 & n2033;
  assign n2035 = ~n1100 & n2034;
  assign n2036 = ~n434 & n2035;
  assign n2037 = ~n1096 & n2036;
  assign n2038 = ~n1095 & n2037;
  assign m1 = n1093 | ~n2038;
  assign n2040 = ~n772 & ~n1288;
  assign n2041 = ~n1043 & n2040;
  assign n2042 = ~n1284 & n2041;
  assign n2043 = ~n769 & n2042;
  assign n2044 = ~n871 & n2043;
  assign n2045 = ~n763 & n2044;
  assign n2046 = ~n1042 & n2045;
  assign n2047 = ~n759 & n2046;
  assign n2048 = ~n755 & n2047;
  assign n2049 = ~n1280 & n2048;
  assign n2050 = ~n1041 & n2049;
  assign n2051 = ~n1037 & n2050;
  assign n2052 = ~n568 & n2051;
  assign n2053 = ~n1032 & n2052;
  assign n2054 = ~n747 & n2053;
  assign n2055 = ~n564 & n2054;
  assign n2056 = ~n746 & n2055;
  assign n2057 = ~n740 & n2056;
  assign n2058 = ~n559 & n2057;
  assign n2059 = ~n556 & n2058;
  assign n2060 = ~n1252 & n2059;
  assign n2061 = ~n739 & n2060;
  assign n2062 = ~n551 & n2061;
  assign n2063 = ~n1235 & n2062;
  assign n2064 = ~n1226 & n2063;
  assign n2065 = ~n738 & n2064;
  assign n2066 = ~n544 & n2065;
  assign n2067 = ~n737 & n2066;
  assign n2068 = ~n1031 & n2067;
  assign n2069 = ~n733 & n2068;
  assign n2070 = ~n540 & n2069;
  assign n2071 = ~n732 & n2070;
  assign n2072 = ~n870 & n2071;
  assign n2073 = ~n1204 & n2072;
  assign n2074 = ~n1202 & n2073;
  assign n2075 = ~n1199 & n2074;
  assign n2076 = ~n1196 & n2075;
  assign n2077 = ~n720 & n2076;
  assign n2078 = ~n1191 & n2077;
  assign n2079 = ~n717 & n2078;
  assign n2080 = ~n1190 & n2079;
  assign n2081 = ~n1184 & n2080;
  assign n2082 = ~n532 & n2081;
  assign n2083 = ~n236 & n2082;
  assign n2084 = ~l2 & n2083;
  assign n2085 = ~n709 & n2084;
  assign n2086 = ~n1173 & n2085;
  assign n2087 = ~n706 & n2086;
  assign n2088 = ~n525 & n2087;
  assign n2089 = ~n1168 & n2088;
  assign n2090 = ~n1160 & n2089;
  assign n2091 = ~n220 & n2090;
  assign n2092 = ~n686 & n2091;
  assign n2093 = ~n865 & n2092;
  assign n2094 = ~n683 & n2093;
  assign n2095 = ~n862 & n2094;
  assign n2096 = ~n678 & n2095;
  assign n2097 = ~n1152 & n2096;
  assign n2098 = ~n1148 & n2097;
  assign n2099 = ~n1144 & n2098;
  assign n2100 = ~n517 & n2099;
  assign n2101 = ~n507 & n2100;
  assign n2102 = ~n676 & n2101;
  assign n2103 = ~n499 & n2102;
  assign n2104 = ~n1136 & n2103;
  assign n2105 = ~n1124 & n2104;
  assign n2106 = ~n1119 & n2105;
  assign n2107 = ~n1114 & n2106;
  assign n2108 = ~n1112 & n2107;
  assign n2109 = ~n674 & n2108;
  assign n2110 = ~n672 & n2109;
  assign n2111 = ~n490 & n2110;
  assign n2112 = ~n487 & n2111;
  assign n2113 = ~n1 & n2112;
  assign n2114 = ~o1 & n2113;
  assign n2115 = ~n664 & n2114;
  assign n2116 = ~n851 & n2115;
  assign n2117 = ~n1110 & n2116;
  assign n2118 = ~n661 & n2117;
  assign n2119 = ~n849 & n2118;
  assign n2120 = ~n654 & n2119;
  assign n2121 = ~n479 & n2120;
  assign n2122 = ~n476 & n2121;
  assign n2123 = ~n846 & n2122;
  assign n2124 = ~n652 & n2123;
  assign n2125 = ~n650 & n2124;
  assign n2126 = ~n402 & n2125;
  assign n2127 = ~n470 & n2126;
  assign n2128 = ~n394 & n2127;
  assign n2129 = ~n386 & n2128;
  assign n2130 = ~n647 & n2129;
  assign n2131 = ~n99 & n2130;
  assign n2132 = ~n382 & n2131;
  assign n2133 = ~n1103 & n2132;
  assign n2134 = ~n640 & n2133;
  assign n2135 = ~n467 & n2134;
  assign n2136 = ~n464 & n2135;
  assign n2137 = ~n453 & n2136;
  assign n2138 = ~n452 & n2137;
  assign n2139 = ~n451 & n2138;
  assign n2140 = ~n449 & n2139;
  assign n2141 = ~n638 & n2140;
  assign n2142 = ~n446 & n2141;
  assign n2143 = ~n1100 & n2142;
  assign n2144 = ~n439 & n2143;
  assign n2145 = ~n436 & n2144;
  assign n2146 = ~n1098 & n2145;
  assign n2147 = ~n434 & n2146;
  assign n2148 = ~n637 & n2147;
  assign n2149 = ~n1097 & n2148;
  assign n2150 = ~n1096 & n2149;
  assign n2151 = ~n1095 & n2150;
  assign n2152 = ~n1094 & n2151;
  assign n2153 = ~n1093 & n2152;
  assign n2154 = ~n1092 & n2153;
  assign p1 = n1091 | ~n2154;
  assign n2156 = ~n733 & ~n769;
  assign q1 = n732 | ~n2156;
  assign n2158 = ~n1284 & ~n1678;
  assign n2159 = ~n1280 & n2158;
  assign n2160 = ~n1235 & n2159;
  assign n2161 = ~n1226 & n2160;
  assign n2162 = ~n1196 & n2161;
  assign n2163 = ~n1193 & n2162;
  assign n2164 = ~n717 & n2163;
  assign n2165 = ~l2 & n2164;
  assign n2166 = ~n709 & n2165;
  assign n2167 = ~n1171 & n2166;
  assign n2168 = ~n706 & n2167;
  assign n2169 = ~n686 & n2168;
  assign n2170 = ~n683 & n2169;
  assign n2171 = ~n678 & n2170;
  assign n2172 = ~n1152 & n2171;
  assign n2173 = ~n1148 & n2172;
  assign n2174 = ~n1127 & n2173;
  assign n2175 = ~n1124 & n2174;
  assign n2176 = ~n1119 & n2175;
  assign n2177 = ~n1114 & n2176;
  assign n2178 = ~n1112 & n2177;
  assign n2179 = ~n674 & n2178;
  assign n2180 = ~n672 & n2179;
  assign n2181 = ~n664 & n2180;
  assign n2182 = ~n1110 & n2181;
  assign n2183 = ~n661 & n2182;
  assign n2184 = ~n654 & n2183;
  assign n2185 = ~n652 & n2184;
  assign s1 = n637 | ~n2185;
  assign n2187 = ~n587 & ~n1538;
  assign n2188 = ~n583 & n2187;
  assign n2189 = ~n576 & n2188;
  assign n2190 = ~n1531 & n2189;
  assign t0 = n1525 | ~n2190;
  assign n2192 = ~n706 & ~n717;
  assign n2193 = ~n678 & n2192;
  assign t1 = n652 | ~n2193;
  assign u0 = n1525 | n1538;
  assign n2196 = ~n1184 & ~n1190;
  assign n2197 = ~n236 & n2196;
  assign n2198 = ~n1168 & n2197;
  assign n2199 = ~n1160 & n2198;
  assign n2200 = ~n220 & n2199;
  assign n2201 = ~n1144 & n2200;
  assign n2202 = ~n1136 & n2201;
  assign n2203 = ~n402 & n2202;
  assign n2204 = ~n394 & n2203;
  assign u1 = n99 | ~n2204;
  assign n2206 = ~n1043 & ~n1284;
  assign n2207 = ~n871 & n2206;
  assign n2208 = ~n1042 & n2207;
  assign n2209 = ~n1280 & n2208;
  assign n2210 = ~n1041 & n2209;
  assign n2211 = ~n1037 & n2210;
  assign n2212 = ~n1032 & n2211;
  assign n2213 = ~n1273 & n2212;
  assign n2214 = ~n1268 & n2213;
  assign n2215 = ~n1260 & n2214;
  assign n2216 = ~n1252 & n2215;
  assign n2217 = ~n1251 & n2216;
  assign n2218 = ~n1244 & n2217;
  assign n2219 = ~n1235 & n2218;
  assign n2220 = ~n1226 & n2219;
  assign n2221 = ~n1216 & n2220;
  assign n2222 = ~n1210 & n2221;
  assign n2223 = ~n1031 & n2222;
  assign n2224 = ~n870 & n2223;
  assign n2225 = ~n1204 & n2224;
  assign n2226 = ~n1202 & n2225;
  assign n2227 = ~n1199 & n2226;
  assign n2228 = ~n1196 & n2227;
  assign n2229 = ~n1193 & n2228;
  assign n2230 = ~n1191 & n2229;
  assign n2231 = ~l2 & n2230;
  assign n2232 = ~n1173 & n2231;
  assign n2233 = ~n1171 & n2232;
  assign n2234 = ~n1127 & n2233;
  assign n2235 = ~n1124 & n2234;
  assign n2236 = ~n1119 & n2235;
  assign n2237 = ~n1100 & n2236;
  assign n2238 = ~n1098 & n2237;
  assign n2239 = ~n1097 & n2238;
  assign n2240 = ~n1096 & n2239;
  assign n2241 = ~n1095 & n2240;
  assign n2242 = ~n1094 & n2241;
  assign n2243 = ~n1093 & n2242;
  assign n2244 = ~n1092 & n2243;
  assign n2245 = ~n1091 & n2244;
  assign v1 = n1090 | ~n2245;
  assign w0 = n576 | n583;
  assign n2248 = n339 & ~n766;
  assign n2249 = ~n572 & n2248;
  assign n2250 = ~i2 & n2249;
  assign n2251 = ~n746 & n2250;
  assign n2252 = ~n295 & n2251;
  assign n2253 = ~n286 & n2252;
  assign n2254 = ~n276 & n2253;
  assign n2255 = ~n265 & n2254;
  assign n2256 = ~n255 & n2255;
  assign n2257 = ~n724 & n2256;
  assign n2258 = ~n245 & n2257;
  assign n2259 = ~n236 & n2258;
  assign n2260 = ~n227 & n2259;
  assign n2261 = ~n220 & n2260;
  assign n2262 = ~n211 & n2261;
  assign n2263 = ~n195 & n2262;
  assign n2264 = ~n143 & n2263;
  assign n2265 = ~n117 & n2264;
  assign w1 = n99 | ~n2265;
  assign n2267 = ~n576 & ~n587;
  assign x0 = n1525 | ~n2267;
  assign n2269 = ~n186 & ~n203;
  assign n2270 = ~n163 & n2269;
  assign n2271 = ~n160 & n2270;
  assign n2272 = ~n152 & n2271;
  assign x1 = n108 | ~n2272;
  assign n2274 = ~n572 & ~n766;
  assign n2275 = ~n746 & n2274;
  assign y0 = n724 | ~n2275;
  assign n2277 = ~n177 & ~n203;
  assign n2278 = ~n170 & n2277;
  assign n2279 = ~n135 & n2278;
  assign n2280 = ~n126 & n2279;
  assign y1 = n108 | ~n2280;
  assign j2 = 1'b0;
  assign v0 = 1'b0;
  assign r1 = l2;
endmodule


