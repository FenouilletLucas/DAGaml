// Benchmark "too_large" written by ABC on Tue May 16 16:07:53 2017

module too_large ( 
    g0, h0, i0, j0, k0, l0, a, b, c, d, e, f, g, h, i, j, k, l, m0, m, n,
    o, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0,
    n0, o0, p0  );
  input  g0, h0, i0, j0, k0, l0, a, b, c, d, e, f, g, h, i, j, k, l, m0,
    m, n, o, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0;
  output n0, o0, p0;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
    n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
    n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
    n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
    n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
    n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
    n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
    n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
    n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
    n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
    n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
    n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
    n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
    n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
    n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
    n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
    n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
    n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
    n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
    n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
    n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
    n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
    n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
    n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
    n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
    n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
    n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
    n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
    n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
    n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
    n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
    n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
    n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
    n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
    n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
    n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
    n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
    n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
    n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
    n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
    n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
    n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
    n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
    n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
    n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
    n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
    n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
    n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
    n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
    n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
    n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
    n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
    n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
    n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
    n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
    n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
    n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
    n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747;
  assign n42 = ~n & ~q;
  assign n43 = ~r & n42;
  assign n44 = w & n43;
  assign n45 = ~x & n44;
  assign n46 = ~y & n45;
  assign n47 = ~a0 & n46;
  assign n48 = ~b0 & n47;
  assign n49 = ~c0 & n48;
  assign n50 = d0 & n49;
  assign n51 = w & ~x;
  assign n52 = ~y & n51;
  assign n53 = ~c0 & n52;
  assign n54 = d0 & n53;
  assign n55 = ~e0 & n54;
  assign n56 = ~f0 & n55;
  assign n57 = ~g0 & n56;
  assign n58 = i0 & n57;
  assign n59 = ~m & ~n;
  assign n60 = ~q & n59;
  assign n61 = w & n60;
  assign n62 = ~x & n61;
  assign n63 = ~y & n62;
  assign n64 = ~a0 & n63;
  assign n65 = ~b0 & n64;
  assign n66 = ~c0 & n65;
  assign n67 = d0 & n66;
  assign n68 = w & ~y;
  assign n69 = ~a0 & n68;
  assign n70 = ~c0 & n69;
  assign n71 = d0 & n70;
  assign n72 = ~e0 & n71;
  assign n73 = ~f0 & n72;
  assign n74 = ~g0 & n73;
  assign n75 = ~i0 & n74;
  assign n76 = ~o & ~q;
  assign n77 = ~r & n76;
  assign n78 = w & n77;
  assign n79 = ~x & n78;
  assign n80 = ~y & n79;
  assign n81 = ~a0 & n80;
  assign n82 = ~b0 & n81;
  assign n83 = ~c0 & n82;
  assign n84 = d0 & n83;
  assign n85 = ~b0 & n46;
  assign n86 = ~c0 & n85;
  assign n87 = d0 & n86;
  assign n88 = i0 & n87;
  assign n89 = ~m & ~o;
  assign n90 = ~q & n89;
  assign n91 = w & n90;
  assign n92 = ~x & n91;
  assign n93 = ~y & n92;
  assign n94 = ~a0 & n93;
  assign n95 = ~b0 & n94;
  assign n96 = ~c0 & n95;
  assign n97 = d0 & n96;
  assign n98 = ~b0 & n63;
  assign n99 = ~c0 & n98;
  assign n100 = d0 & n99;
  assign n101 = i0 & n100;
  assign n102 = w & ~c0;
  assign n103 = d0 & n102;
  assign n104 = ~e0 & n103;
  assign n105 = ~f0 & n104;
  assign n106 = ~g0 & n105;
  assign n107 = ~i0 & n106;
  assign n108 = j0 & n107;
  assign n109 = ~x & n77;
  assign n110 = ~y & n109;
  assign n111 = z & n110;
  assign n112 = ~a0 & n111;
  assign n113 = ~b0 & n112;
  assign n114 = ~c0 & n113;
  assign n115 = h0 & n114;
  assign n116 = o & ~x;
  assign n117 = ~y & n116;
  assign n118 = ~c0 & n117;
  assign n119 = ~d0 & n118;
  assign n120 = ~e0 & n119;
  assign n121 = ~f0 & n120;
  assign n122 = ~g0 & n121;
  assign n123 = h0 & n122;
  assign n124 = i0 & n123;
  assign n125 = ~x & n90;
  assign n126 = ~y & n125;
  assign n127 = z & n126;
  assign n128 = ~a0 & n127;
  assign n129 = ~b0 & n128;
  assign n130 = ~c0 & n129;
  assign n131 = h0 & n130;
  assign n132 = ~b0 & n80;
  assign n133 = ~c0 & n132;
  assign n134 = d0 & n133;
  assign n135 = i0 & n134;
  assign n136 = ~b0 & n93;
  assign n137 = ~c0 & n136;
  assign n138 = d0 & n137;
  assign n139 = i0 & n138;
  assign n140 = ~n & o;
  assign n141 = ~q & n140;
  assign n142 = ~r & n141;
  assign n143 = ~x & n142;
  assign n144 = ~y & n143;
  assign n145 = ~b0 & n144;
  assign n146 = ~c0 & n145;
  assign n147 = ~d0 & n146;
  assign n148 = h0 & n147;
  assign n149 = i0 & n148;
  assign n150 = o & n59;
  assign n151 = ~q & n150;
  assign n152 = ~x & n151;
  assign n153 = ~y & n152;
  assign n154 = ~b0 & n153;
  assign n155 = ~c0 & n154;
  assign n156 = ~d0 & n155;
  assign n157 = h0 & n156;
  assign n158 = i0 & n157;
  assign n159 = o & ~c0;
  assign n160 = ~d0 & n159;
  assign n161 = ~e0 & n160;
  assign n162 = ~f0 & n161;
  assign n163 = ~g0 & n162;
  assign n164 = h0 & n163;
  assign n165 = ~i0 & n164;
  assign n166 = j0 & n165;
  assign n167 = ~x & ~y;
  assign n168 = z & n167;
  assign n169 = ~c0 & n168;
  assign n170 = ~d0 & n169;
  assign n171 = ~e0 & n170;
  assign n172 = ~f0 & n171;
  assign n173 = ~g0 & n172;
  assign n174 = h0 & n173;
  assign n175 = i0 & n174;
  assign n176 = ~y & z;
  assign n177 = ~a0 & n176;
  assign n178 = ~c0 & n177;
  assign n179 = ~d0 & n178;
  assign n180 = ~e0 & n179;
  assign n181 = ~f0 & n180;
  assign n182 = ~g0 & n181;
  assign n183 = h0 & n182;
  assign n184 = ~i0 & n183;
  assign n185 = z & ~c0;
  assign n186 = ~d0 & n185;
  assign n187 = ~e0 & n186;
  assign n188 = ~f0 & n187;
  assign n189 = ~g0 & n188;
  assign n190 = h0 & n189;
  assign n191 = ~i0 & n190;
  assign n192 = j0 & n191;
  assign n193 = ~b0 & n111;
  assign n194 = ~c0 & n193;
  assign n195 = ~d0 & n194;
  assign n196 = h0 & n195;
  assign n197 = i0 & n196;
  assign n198 = ~b0 & n45;
  assign n199 = ~c0 & n198;
  assign n200 = d0 & n199;
  assign n201 = ~i0 & n200;
  assign n202 = j0 & n201;
  assign n203 = ~b0 & n127;
  assign n204 = ~c0 & n203;
  assign n205 = ~d0 & n204;
  assign n206 = h0 & n205;
  assign n207 = i0 & n206;
  assign n208 = ~b0 & n62;
  assign n209 = ~c0 & n208;
  assign n210 = d0 & n209;
  assign n211 = ~i0 & n210;
  assign n212 = j0 & n211;
  assign n213 = ~b0 & n79;
  assign n214 = ~c0 & n213;
  assign n215 = d0 & n214;
  assign n216 = ~i0 & n215;
  assign n217 = j0 & n216;
  assign n218 = ~b0 & n92;
  assign n219 = ~c0 & n218;
  assign n220 = d0 & n219;
  assign n221 = ~i0 & n220;
  assign n222 = j0 & n221;
  assign n223 = ~b0 & n143;
  assign n224 = ~c0 & n223;
  assign n225 = ~d0 & n224;
  assign n226 = h0 & n225;
  assign n227 = ~i0 & n226;
  assign n228 = j0 & n227;
  assign n229 = ~b0 & n152;
  assign n230 = ~c0 & n229;
  assign n231 = ~d0 & n230;
  assign n232 = h0 & n231;
  assign n233 = ~i0 & n232;
  assign n234 = j0 & n233;
  assign n235 = u & n43;
  assign n236 = ~v & n235;
  assign n237 = ~w & n236;
  assign n238 = ~x & n237;
  assign n239 = ~y & n238;
  assign n240 = ~a0 & n239;
  assign n241 = ~b0 & n240;
  assign n242 = ~c0 & n241;
  assign n243 = d0 & n242;
  assign n244 = u & n60;
  assign n245 = ~v & n244;
  assign n246 = ~w & n245;
  assign n247 = ~x & n246;
  assign n248 = ~y & n247;
  assign n249 = ~a0 & n248;
  assign n250 = ~b0 & n249;
  assign n251 = ~c0 & n250;
  assign n252 = d0 & n251;
  assign n253 = u & n77;
  assign n254 = ~v & n253;
  assign n255 = ~w & n254;
  assign n256 = ~x & n255;
  assign n257 = ~y & n256;
  assign n258 = ~a0 & n257;
  assign n259 = ~b0 & n258;
  assign n260 = ~c0 & n259;
  assign n261 = d0 & n260;
  assign n262 = u & n90;
  assign n263 = ~v & n262;
  assign n264 = ~w & n263;
  assign n265 = ~x & n264;
  assign n266 = ~y & n265;
  assign n267 = ~a0 & n266;
  assign n268 = ~b0 & n267;
  assign n269 = ~c0 & n268;
  assign n270 = d0 & n269;
  assign n271 = z & n109;
  assign n272 = ~b0 & n271;
  assign n273 = ~c0 & n272;
  assign n274 = ~d0 & n273;
  assign n275 = h0 & n274;
  assign n276 = ~i0 & n275;
  assign n277 = j0 & n276;
  assign n278 = z & n125;
  assign n279 = ~b0 & n278;
  assign n280 = ~c0 & n279;
  assign n281 = ~d0 & n280;
  assign n282 = h0 & n281;
  assign n283 = ~i0 & n282;
  assign n284 = j0 & n283;
  assign n285 = c & ~m;
  assign n286 = ~n & n285;
  assign n287 = ~q & n286;
  assign n288 = ~u & n287;
  assign n289 = ~v & n288;
  assign n290 = ~x & n289;
  assign n291 = ~y & n290;
  assign n292 = ~a0 & n291;
  assign n293 = ~b0 & n292;
  assign n294 = ~c0 & n293;
  assign n295 = d0 & n294;
  assign n296 = ~o & n285;
  assign n297 = ~q & n296;
  assign n298 = ~u & n297;
  assign n299 = ~v & n298;
  assign n300 = ~x & n299;
  assign n301 = ~y & n300;
  assign n302 = ~a0 & n301;
  assign n303 = ~b0 & n302;
  assign n304 = ~c0 & n303;
  assign n305 = d0 & n304;
  assign n306 = ~e & ~f;
  assign n307 = ~g & n306;
  assign n308 = ~j & n307;
  assign n309 = ~n & n308;
  assign n310 = ~q & n309;
  assign n311 = ~r & n310;
  assign n312 = ~x & n311;
  assign n313 = ~b0 & n312;
  assign n314 = ~c0 & n313;
  assign n315 = d0 & n314;
  assign n316 = ~j0 & n315;
  assign n317 = k0 & n316;
  assign n318 = d & n317;
  assign n319 = ~s & n318;
  assign n320 = ~g0 & n319;
  assign n321 = ~v & n320;
  assign n322 = ~y & n321;
  assign n323 = ~a0 & n322;
  assign n324 = ~h & n307;
  assign n325 = ~j & n324;
  assign n326 = ~n & n325;
  assign n327 = ~q & n326;
  assign n328 = ~r & n327;
  assign n329 = ~x & n328;
  assign n330 = ~b0 & n329;
  assign n331 = ~c0 & n330;
  assign n332 = d0 & n331;
  assign n333 = k0 & n332;
  assign n334 = d & n333;
  assign n335 = ~s & n334;
  assign n336 = ~g0 & n335;
  assign n337 = ~v & n336;
  assign n338 = ~y & n337;
  assign n339 = ~a0 & n338;
  assign n340 = ~l & n308;
  assign n341 = ~n & n340;
  assign n342 = ~q & n341;
  assign n343 = ~r & n342;
  assign n344 = ~t & n343;
  assign n345 = ~x & n344;
  assign n346 = ~b0 & n345;
  assign n347 = ~c0 & n346;
  assign n348 = d0 & n347;
  assign n349 = ~j0 & n348;
  assign n350 = k0 & n349;
  assign n351 = ~g0 & n350;
  assign n352 = ~v & n351;
  assign n353 = ~y & n352;
  assign n354 = ~a0 & n353;
  assign n355 = ~l & n325;
  assign n356 = ~n & n355;
  assign n357 = ~q & n356;
  assign n358 = ~r & n357;
  assign n359 = ~t & n358;
  assign n360 = ~x & n359;
  assign n361 = ~b0 & n360;
  assign n362 = ~c0 & n361;
  assign n363 = d0 & n362;
  assign n364 = k0 & n363;
  assign n365 = ~g0 & n364;
  assign n366 = ~v & n365;
  assign n367 = ~y & n366;
  assign n368 = ~a0 & n367;
  assign n369 = ~i & n307;
  assign n370 = ~j & n369;
  assign n371 = ~n & n370;
  assign n372 = ~q & n371;
  assign n373 = ~r & n372;
  assign n374 = ~x & n373;
  assign n375 = ~b0 & n374;
  assign n376 = ~c0 & n375;
  assign n377 = d0 & n376;
  assign n378 = ~j0 & n377;
  assign n379 = k0 & n378;
  assign n380 = d & n379;
  assign n381 = ~s & n380;
  assign n382 = ~v & n381;
  assign n383 = ~y & n382;
  assign n384 = ~a0 & n383;
  assign n385 = ~i & n324;
  assign n386 = ~j & n385;
  assign n387 = ~n & n386;
  assign n388 = ~q & n387;
  assign n389 = ~r & n388;
  assign n390 = ~x & n389;
  assign n391 = ~b0 & n390;
  assign n392 = ~c0 & n391;
  assign n393 = d0 & n392;
  assign n394 = k0 & n393;
  assign n395 = d & n394;
  assign n396 = ~s & n395;
  assign n397 = ~v & n396;
  assign n398 = ~y & n397;
  assign n399 = ~a0 & n398;
  assign n400 = ~l & n370;
  assign n401 = ~n & n400;
  assign n402 = ~q & n401;
  assign n403 = ~r & n402;
  assign n404 = ~t & n403;
  assign n405 = ~x & n404;
  assign n406 = ~b0 & n405;
  assign n407 = ~c0 & n406;
  assign n408 = d0 & n407;
  assign n409 = ~j0 & n408;
  assign n410 = k0 & n409;
  assign n411 = ~v & n410;
  assign n412 = ~y & n411;
  assign n413 = ~a0 & n412;
  assign n414 = ~l & n386;
  assign n415 = ~n & n414;
  assign n416 = ~q & n415;
  assign n417 = ~r & n416;
  assign n418 = ~t & n417;
  assign n419 = ~x & n418;
  assign n420 = ~b0 & n419;
  assign n421 = ~c0 & n420;
  assign n422 = d0 & n421;
  assign n423 = k0 & n422;
  assign n424 = ~v & n423;
  assign n425 = ~y & n424;
  assign n426 = ~a0 & n425;
  assign n427 = ~c & ~e;
  assign n428 = ~f & n427;
  assign n429 = ~g & n428;
  assign n430 = ~j & n429;
  assign n431 = ~n & n430;
  assign n432 = ~q & n431;
  assign n433 = ~r & n432;
  assign n434 = ~x & n433;
  assign n435 = ~b0 & n434;
  assign n436 = ~c0 & n435;
  assign n437 = ~d0 & n436;
  assign n438 = ~j0 & n437;
  assign n439 = k0 & n438;
  assign n440 = d & n439;
  assign n441 = ~s & n440;
  assign n442 = ~g0 & n441;
  assign n443 = ~y & n442;
  assign n444 = ~a0 & n443;
  assign n445 = ~l & n430;
  assign n446 = ~n & n445;
  assign n447 = ~q & n446;
  assign n448 = ~r & n447;
  assign n449 = ~t & n448;
  assign n450 = ~x & n449;
  assign n451 = ~b0 & n450;
  assign n452 = ~c0 & n451;
  assign n453 = ~d0 & n452;
  assign n454 = ~j0 & n453;
  assign n455 = k0 & n454;
  assign n456 = ~g0 & n455;
  assign n457 = ~y & n456;
  assign n458 = ~a0 & n457;
  assign n459 = ~i & n429;
  assign n460 = ~j & n459;
  assign n461 = ~n & n460;
  assign n462 = ~q & n461;
  assign n463 = ~r & n462;
  assign n464 = ~x & n463;
  assign n465 = ~b0 & n464;
  assign n466 = ~c0 & n465;
  assign n467 = ~d0 & n466;
  assign n468 = ~j0 & n467;
  assign n469 = k0 & n468;
  assign n470 = d & n469;
  assign n471 = ~s & n470;
  assign n472 = ~y & n471;
  assign n473 = ~a0 & n472;
  assign n474 = ~l & n460;
  assign n475 = ~n & n474;
  assign n476 = ~q & n475;
  assign n477 = ~r & n476;
  assign n478 = ~t & n477;
  assign n479 = ~x & n478;
  assign n480 = ~b0 & n479;
  assign n481 = ~c0 & n480;
  assign n482 = ~d0 & n481;
  assign n483 = ~j0 & n482;
  assign n484 = k0 & n483;
  assign n485 = ~y & n484;
  assign n486 = ~a0 & n485;
  assign n487 = i0 & n437;
  assign n488 = ~j0 & n487;
  assign n489 = k0 & n488;
  assign n490 = d & n489;
  assign n491 = ~s & n490;
  assign n492 = ~g0 & n491;
  assign n493 = ~y & n492;
  assign n494 = ~h & n429;
  assign n495 = ~j & n494;
  assign n496 = ~n & n495;
  assign n497 = ~q & n496;
  assign n498 = ~r & n497;
  assign n499 = ~x & n498;
  assign n500 = ~b0 & n499;
  assign n501 = ~c0 & n500;
  assign n502 = ~d0 & n501;
  assign n503 = i0 & n502;
  assign n504 = k0 & n503;
  assign n505 = d & n504;
  assign n506 = ~s & n505;
  assign n507 = ~g0 & n506;
  assign n508 = ~y & n507;
  assign n509 = i0 & n453;
  assign n510 = ~j0 & n509;
  assign n511 = k0 & n510;
  assign n512 = ~g0 & n511;
  assign n513 = ~y & n512;
  assign n514 = ~l & n495;
  assign n515 = ~n & n514;
  assign n516 = ~q & n515;
  assign n517 = ~r & n516;
  assign n518 = ~t & n517;
  assign n519 = ~x & n518;
  assign n520 = ~b0 & n519;
  assign n521 = ~c0 & n520;
  assign n522 = ~d0 & n521;
  assign n523 = i0 & n522;
  assign n524 = k0 & n523;
  assign n525 = ~g0 & n524;
  assign n526 = ~y & n525;
  assign n527 = i0 & n467;
  assign n528 = ~j0 & n527;
  assign n529 = k0 & n528;
  assign n530 = d & n529;
  assign n531 = ~s & n530;
  assign n532 = ~y & n531;
  assign n533 = ~i & n494;
  assign n534 = ~j & n533;
  assign n535 = ~n & n534;
  assign n536 = ~q & n535;
  assign n537 = ~r & n536;
  assign n538 = ~x & n537;
  assign n539 = ~b0 & n538;
  assign n540 = ~c0 & n539;
  assign n541 = ~d0 & n540;
  assign n542 = i0 & n541;
  assign n543 = k0 & n542;
  assign n544 = d & n543;
  assign n545 = ~s & n544;
  assign n546 = ~y & n545;
  assign n547 = i0 & n482;
  assign n548 = ~j0 & n547;
  assign n549 = k0 & n548;
  assign n550 = ~y & n549;
  assign n551 = ~l & n534;
  assign n552 = ~n & n551;
  assign n553 = ~q & n552;
  assign n554 = ~r & n553;
  assign n555 = ~t & n554;
  assign n556 = ~x & n555;
  assign n557 = ~b0 & n556;
  assign n558 = ~c0 & n557;
  assign n559 = ~d0 & n558;
  assign n560 = i0 & n559;
  assign n561 = k0 & n560;
  assign n562 = ~y & n561;
  assign n563 = ~i0 & n502;
  assign n564 = j0 & n563;
  assign n565 = k0 & n564;
  assign n566 = d & n565;
  assign n567 = ~s & n566;
  assign n568 = ~g0 & n567;
  assign n569 = ~i0 & n522;
  assign n570 = j0 & n569;
  assign n571 = k0 & n570;
  assign n572 = ~g0 & n571;
  assign n573 = ~i0 & n541;
  assign n574 = j0 & n573;
  assign n575 = k0 & n574;
  assign n576 = d & n575;
  assign n577 = ~s & n576;
  assign n578 = ~i0 & n559;
  assign n579 = j0 & n578;
  assign n580 = k0 & n579;
  assign n581 = ~q & n429;
  assign n582 = ~r & n581;
  assign n583 = ~x & n582;
  assign n584 = ~b0 & n583;
  assign n585 = ~c0 & n584;
  assign n586 = ~j0 & n585;
  assign n587 = k0 & n586;
  assign n588 = ~g0 & n587;
  assign n589 = ~v & n588;
  assign n590 = ~y & n589;
  assign n591 = ~a0 & n590;
  assign n592 = ~o & n591;
  assign n593 = ~b & n592;
  assign n594 = ~f0 & n593;
  assign n595 = ~q & n459;
  assign n596 = ~r & n595;
  assign n597 = ~x & n596;
  assign n598 = ~b0 & n597;
  assign n599 = ~c0 & n598;
  assign n600 = ~j0 & n599;
  assign n601 = k0 & n600;
  assign n602 = ~v & n601;
  assign n603 = ~y & n602;
  assign n604 = ~a0 & n603;
  assign n605 = ~o & n604;
  assign n606 = ~b & n605;
  assign n607 = ~f0 & n606;
  assign n608 = ~d0 & n585;
  assign n609 = ~j0 & n608;
  assign n610 = k0 & n609;
  assign n611 = ~g0 & n610;
  assign n612 = ~y & n611;
  assign n613 = ~a0 & n612;
  assign n614 = ~o & n613;
  assign n615 = ~b & n614;
  assign n616 = ~f0 & n615;
  assign n617 = ~d0 & n599;
  assign n618 = ~j0 & n617;
  assign n619 = k0 & n618;
  assign n620 = ~y & n619;
  assign n621 = ~a0 & n620;
  assign n622 = ~o & n621;
  assign n623 = ~b & n622;
  assign n624 = ~f0 & n623;
  assign n625 = i0 & n608;
  assign n626 = ~j0 & n625;
  assign n627 = k0 & n626;
  assign n628 = ~g0 & n627;
  assign n629 = ~y & n628;
  assign n630 = ~o & n629;
  assign n631 = ~b & n630;
  assign n632 = ~f0 & n631;
  assign n633 = i0 & n617;
  assign n634 = ~j0 & n633;
  assign n635 = k0 & n634;
  assign n636 = ~y & n635;
  assign n637 = ~o & n636;
  assign n638 = ~b & n637;
  assign n639 = ~f0 & n638;
  assign n640 = ~n & n429;
  assign n641 = ~q & n640;
  assign n642 = ~r & n641;
  assign n643 = ~x & n642;
  assign n644 = ~b0 & n643;
  assign n645 = ~c0 & n644;
  assign n646 = ~j0 & n645;
  assign n647 = k0 & n646;
  assign n648 = ~g0 & n647;
  assign n649 = ~v & n648;
  assign n650 = ~y & n649;
  assign n651 = ~a0 & n650;
  assign n652 = ~b & n651;
  assign n653 = ~f0 & n652;
  assign n654 = ~n & n459;
  assign n655 = ~q & n654;
  assign n656 = ~r & n655;
  assign n657 = ~x & n656;
  assign n658 = ~b0 & n657;
  assign n659 = ~c0 & n658;
  assign n660 = ~j0 & n659;
  assign n661 = k0 & n660;
  assign n662 = ~v & n661;
  assign n663 = ~y & n662;
  assign n664 = ~a0 & n663;
  assign n665 = ~b & n664;
  assign n666 = ~f0 & n665;
  assign n667 = ~d0 & n645;
  assign n668 = ~j0 & n667;
  assign n669 = k0 & n668;
  assign n670 = ~g0 & n669;
  assign n671 = ~y & n670;
  assign n672 = ~a0 & n671;
  assign n673 = ~b & n672;
  assign n674 = ~f0 & n673;
  assign n675 = ~d0 & n659;
  assign n676 = ~j0 & n675;
  assign n677 = k0 & n676;
  assign n678 = ~y & n677;
  assign n679 = ~a0 & n678;
  assign n680 = ~b & n679;
  assign n681 = ~f0 & n680;
  assign n682 = i0 & n667;
  assign n683 = ~j0 & n682;
  assign n684 = k0 & n683;
  assign n685 = ~g0 & n684;
  assign n686 = ~y & n685;
  assign n687 = ~b & n686;
  assign n688 = ~f0 & n687;
  assign n689 = i0 & n675;
  assign n690 = ~j0 & n689;
  assign n691 = k0 & n690;
  assign n692 = ~y & n691;
  assign n693 = ~b & n692;
  assign n694 = ~f0 & n693;
  assign n695 = ~g0 & n317;
  assign n696 = ~v & n695;
  assign n697 = ~y & n696;
  assign n698 = ~a0 & n697;
  assign n699 = ~k & n698;
  assign n700 = ~g0 & n333;
  assign n701 = ~v & n700;
  assign n702 = ~y & n701;
  assign n703 = ~a0 & n702;
  assign n704 = ~k & n703;
  assign n705 = ~v & n379;
  assign n706 = ~y & n705;
  assign n707 = ~a0 & n706;
  assign n708 = ~k & n707;
  assign n709 = ~v & n394;
  assign n710 = ~y & n709;
  assign n711 = ~a0 & n710;
  assign n712 = ~k & n711;
  assign n713 = ~g0 & n439;
  assign n714 = ~y & n713;
  assign n715 = ~a0 & n714;
  assign n716 = ~k & n715;
  assign n717 = ~y & n469;
  assign n718 = ~a0 & n717;
  assign n719 = ~k & n718;
  assign n720 = ~g0 & n489;
  assign n721 = ~y & n720;
  assign n722 = ~k & n721;
  assign n723 = ~g0 & n504;
  assign n724 = ~y & n723;
  assign n725 = ~k & n724;
  assign n726 = ~y & n529;
  assign n727 = ~k & n726;
  assign n728 = ~y & n543;
  assign n729 = ~k & n728;
  assign n730 = ~g0 & n565;
  assign n731 = ~k & n730;
  assign n732 = ~k & n575;
  assign n733 = n & n308;
  assign n734 = ~q & n733;
  assign n735 = ~r & n734;
  assign n736 = ~x & n735;
  assign n737 = ~b0 & n736;
  assign n738 = ~c0 & n737;
  assign n739 = d0 & n738;
  assign n740 = ~j0 & n739;
  assign n741 = k0 & n740;
  assign n742 = ~g0 & n741;
  assign n743 = ~v & n742;
  assign n744 = ~y & n743;
  assign n745 = ~a0 & n744;
  assign n746 = ~o & n745;
  assign n747 = n & n325;
  assign n748 = ~q & n747;
  assign n749 = ~r & n748;
  assign n750 = ~x & n749;
  assign n751 = ~b0 & n750;
  assign n752 = ~c0 & n751;
  assign n753 = d0 & n752;
  assign n754 = k0 & n753;
  assign n755 = ~g0 & n754;
  assign n756 = ~v & n755;
  assign n757 = ~y & n756;
  assign n758 = ~a0 & n757;
  assign n759 = ~o & n758;
  assign n760 = n & n370;
  assign n761 = ~q & n760;
  assign n762 = ~r & n761;
  assign n763 = ~x & n762;
  assign n764 = ~b0 & n763;
  assign n765 = ~c0 & n764;
  assign n766 = d0 & n765;
  assign n767 = ~j0 & n766;
  assign n768 = k0 & n767;
  assign n769 = ~v & n768;
  assign n770 = ~y & n769;
  assign n771 = ~a0 & n770;
  assign n772 = ~o & n771;
  assign n773 = n & n386;
  assign n774 = ~q & n773;
  assign n775 = ~r & n774;
  assign n776 = ~x & n775;
  assign n777 = ~b0 & n776;
  assign n778 = ~c0 & n777;
  assign n779 = d0 & n778;
  assign n780 = k0 & n779;
  assign n781 = ~v & n780;
  assign n782 = ~y & n781;
  assign n783 = ~a0 & n782;
  assign n784 = ~o & n783;
  assign n785 = n & n430;
  assign n786 = ~q & n785;
  assign n787 = ~r & n786;
  assign n788 = ~x & n787;
  assign n789 = ~b0 & n788;
  assign n790 = ~c0 & n789;
  assign n791 = ~d0 & n790;
  assign n792 = ~j0 & n791;
  assign n793 = k0 & n792;
  assign n794 = ~g0 & n793;
  assign n795 = ~y & n794;
  assign n796 = ~a0 & n795;
  assign n797 = ~o & n796;
  assign n798 = n & n460;
  assign n799 = ~q & n798;
  assign n800 = ~r & n799;
  assign n801 = ~x & n800;
  assign n802 = ~b0 & n801;
  assign n803 = ~c0 & n802;
  assign n804 = ~d0 & n803;
  assign n805 = ~j0 & n804;
  assign n806 = k0 & n805;
  assign n807 = ~y & n806;
  assign n808 = ~a0 & n807;
  assign n809 = ~o & n808;
  assign n810 = i0 & n791;
  assign n811 = ~j0 & n810;
  assign n812 = k0 & n811;
  assign n813 = ~g0 & n812;
  assign n814 = ~y & n813;
  assign n815 = ~o & n814;
  assign n816 = n & n495;
  assign n817 = ~q & n816;
  assign n818 = ~r & n817;
  assign n819 = ~x & n818;
  assign n820 = ~b0 & n819;
  assign n821 = ~c0 & n820;
  assign n822 = ~d0 & n821;
  assign n823 = i0 & n822;
  assign n824 = k0 & n823;
  assign n825 = ~g0 & n824;
  assign n826 = ~y & n825;
  assign n827 = ~o & n826;
  assign n828 = i0 & n804;
  assign n829 = ~j0 & n828;
  assign n830 = k0 & n829;
  assign n831 = ~y & n830;
  assign n832 = ~o & n831;
  assign n833 = n & n534;
  assign n834 = ~q & n833;
  assign n835 = ~r & n834;
  assign n836 = ~x & n835;
  assign n837 = ~b0 & n836;
  assign n838 = ~c0 & n837;
  assign n839 = ~d0 & n838;
  assign n840 = i0 & n839;
  assign n841 = k0 & n840;
  assign n842 = ~y & n841;
  assign n843 = ~o & n842;
  assign n844 = ~i0 & n822;
  assign n845 = j0 & n844;
  assign n846 = k0 & n845;
  assign n847 = ~g0 & n846;
  assign n848 = ~o & n847;
  assign n849 = ~i0 & n839;
  assign n850 = j0 & n849;
  assign n851 = k0 & n850;
  assign n852 = ~o & n851;
  assign n853 = ~q & n307;
  assign n854 = ~x & n853;
  assign n855 = ~b0 & n854;
  assign n856 = ~c0 & n855;
  assign n857 = d0 & n856;
  assign n858 = ~j0 & n857;
  assign n859 = k0 & n858;
  assign n860 = ~g0 & n859;
  assign n861 = ~v & n860;
  assign n862 = ~y & n861;
  assign n863 = ~a0 & n862;
  assign n864 = ~o & n863;
  assign n865 = ~f0 & n864;
  assign n866 = ~m & n865;
  assign n867 = ~q & n369;
  assign n868 = ~x & n867;
  assign n869 = ~b0 & n868;
  assign n870 = ~c0 & n869;
  assign n871 = d0 & n870;
  assign n872 = ~j0 & n871;
  assign n873 = k0 & n872;
  assign n874 = ~v & n873;
  assign n875 = ~y & n874;
  assign n876 = ~a0 & n875;
  assign n877 = ~o & n876;
  assign n878 = ~f0 & n877;
  assign n879 = ~m & n878;
  assign n880 = ~x & n581;
  assign n881 = ~b0 & n880;
  assign n882 = ~c0 & n881;
  assign n883 = ~d0 & n882;
  assign n884 = ~j0 & n883;
  assign n885 = k0 & n884;
  assign n886 = ~g0 & n885;
  assign n887 = ~y & n886;
  assign n888 = ~a0 & n887;
  assign n889 = ~o & n888;
  assign n890 = ~f0 & n889;
  assign n891 = ~m & n890;
  assign n892 = ~x & n595;
  assign n893 = ~b0 & n892;
  assign n894 = ~c0 & n893;
  assign n895 = ~d0 & n894;
  assign n896 = ~j0 & n895;
  assign n897 = k0 & n896;
  assign n898 = ~y & n897;
  assign n899 = ~a0 & n898;
  assign n900 = ~o & n899;
  assign n901 = ~f0 & n900;
  assign n902 = ~m & n901;
  assign n903 = i0 & n883;
  assign n904 = ~j0 & n903;
  assign n905 = k0 & n904;
  assign n906 = ~g0 & n905;
  assign n907 = ~y & n906;
  assign n908 = ~o & n907;
  assign n909 = ~f0 & n908;
  assign n910 = ~m & n909;
  assign n911 = i0 & n895;
  assign n912 = ~j0 & n911;
  assign n913 = k0 & n912;
  assign n914 = ~y & n913;
  assign n915 = ~o & n914;
  assign n916 = ~f0 & n915;
  assign n917 = ~m & n916;
  assign n918 = ~n & n307;
  assign n919 = ~q & n918;
  assign n920 = ~x & n919;
  assign n921 = ~b0 & n920;
  assign n922 = ~c0 & n921;
  assign n923 = d0 & n922;
  assign n924 = ~j0 & n923;
  assign n925 = k0 & n924;
  assign n926 = ~g0 & n925;
  assign n927 = ~v & n926;
  assign n928 = ~y & n927;
  assign n929 = ~a0 & n928;
  assign n930 = ~f0 & n929;
  assign n931 = ~m & n930;
  assign n932 = ~n & n369;
  assign n933 = ~q & n932;
  assign n934 = ~x & n933;
  assign n935 = ~b0 & n934;
  assign n936 = ~c0 & n935;
  assign n937 = d0 & n936;
  assign n938 = ~j0 & n937;
  assign n939 = k0 & n938;
  assign n940 = ~v & n939;
  assign n941 = ~y & n940;
  assign n942 = ~a0 & n941;
  assign n943 = ~f0 & n942;
  assign n944 = ~m & n943;
  assign n945 = ~x & n641;
  assign n946 = ~b0 & n945;
  assign n947 = ~c0 & n946;
  assign n948 = ~d0 & n947;
  assign n949 = ~j0 & n948;
  assign n950 = k0 & n949;
  assign n951 = ~g0 & n950;
  assign n952 = ~y & n951;
  assign n953 = ~a0 & n952;
  assign n954 = ~f0 & n953;
  assign n955 = ~m & n954;
  assign n956 = ~x & n655;
  assign n957 = ~b0 & n956;
  assign n958 = ~c0 & n957;
  assign n959 = ~d0 & n958;
  assign n960 = ~j0 & n959;
  assign n961 = k0 & n960;
  assign n962 = ~y & n961;
  assign n963 = ~a0 & n962;
  assign n964 = ~f0 & n963;
  assign n965 = ~m & n964;
  assign n966 = i0 & n948;
  assign n967 = ~j0 & n966;
  assign n968 = k0 & n967;
  assign n969 = ~g0 & n968;
  assign n970 = ~y & n969;
  assign n971 = ~f0 & n970;
  assign n972 = ~m & n971;
  assign n973 = i0 & n959;
  assign n974 = ~j0 & n973;
  assign n975 = k0 & n974;
  assign n976 = ~y & n975;
  assign n977 = ~f0 & n976;
  assign n978 = ~m & n977;
  assign n979 = ~q & n494;
  assign n980 = ~r & n979;
  assign n981 = ~x & n980;
  assign n982 = ~b0 & n981;
  assign n983 = ~c0 & n982;
  assign n984 = k0 & n983;
  assign n985 = ~g0 & n984;
  assign n986 = ~v & n985;
  assign n987 = ~y & n986;
  assign n988 = ~a0 & n987;
  assign n989 = ~o & n988;
  assign n990 = ~b & n989;
  assign n991 = ~q & n533;
  assign n992 = ~r & n991;
  assign n993 = ~x & n992;
  assign n994 = ~b0 & n993;
  assign n995 = ~c0 & n994;
  assign n996 = k0 & n995;
  assign n997 = ~v & n996;
  assign n998 = ~y & n997;
  assign n999 = ~a0 & n998;
  assign n1000 = ~o & n999;
  assign n1001 = ~b & n1000;
  assign n1002 = ~d0 & n983;
  assign n1003 = k0 & n1002;
  assign n1004 = ~g0 & n1003;
  assign n1005 = ~y & n1004;
  assign n1006 = ~a0 & n1005;
  assign n1007 = ~o & n1006;
  assign n1008 = ~b & n1007;
  assign n1009 = ~d0 & n995;
  assign n1010 = k0 & n1009;
  assign n1011 = ~y & n1010;
  assign n1012 = ~a0 & n1011;
  assign n1013 = ~o & n1012;
  assign n1014 = ~b & n1013;
  assign n1015 = i0 & n1002;
  assign n1016 = k0 & n1015;
  assign n1017 = ~g0 & n1016;
  assign n1018 = ~y & n1017;
  assign n1019 = ~o & n1018;
  assign n1020 = ~b & n1019;
  assign n1021 = i0 & n1009;
  assign n1022 = k0 & n1021;
  assign n1023 = ~y & n1022;
  assign n1024 = ~o & n1023;
  assign n1025 = ~b & n1024;
  assign n1026 = ~i0 & n1002;
  assign n1027 = j0 & n1026;
  assign n1028 = k0 & n1027;
  assign n1029 = ~g0 & n1028;
  assign n1030 = ~o & n1029;
  assign n1031 = ~b & n1030;
  assign n1032 = ~i0 & n1009;
  assign n1033 = j0 & n1032;
  assign n1034 = k0 & n1033;
  assign n1035 = ~o & n1034;
  assign n1036 = ~b & n1035;
  assign n1037 = ~n & n494;
  assign n1038 = ~q & n1037;
  assign n1039 = ~r & n1038;
  assign n1040 = ~x & n1039;
  assign n1041 = ~b0 & n1040;
  assign n1042 = ~c0 & n1041;
  assign n1043 = k0 & n1042;
  assign n1044 = ~g0 & n1043;
  assign n1045 = ~v & n1044;
  assign n1046 = ~y & n1045;
  assign n1047 = ~a0 & n1046;
  assign n1048 = ~b & n1047;
  assign n1049 = ~n & n533;
  assign n1050 = ~q & n1049;
  assign n1051 = ~r & n1050;
  assign n1052 = ~x & n1051;
  assign n1053 = ~b0 & n1052;
  assign n1054 = ~c0 & n1053;
  assign n1055 = k0 & n1054;
  assign n1056 = ~v & n1055;
  assign n1057 = ~y & n1056;
  assign n1058 = ~a0 & n1057;
  assign n1059 = ~b & n1058;
  assign n1060 = ~d0 & n1042;
  assign n1061 = k0 & n1060;
  assign n1062 = ~g0 & n1061;
  assign n1063 = ~y & n1062;
  assign n1064 = ~a0 & n1063;
  assign n1065 = ~b & n1064;
  assign n1066 = ~d0 & n1054;
  assign n1067 = k0 & n1066;
  assign n1068 = ~y & n1067;
  assign n1069 = ~a0 & n1068;
  assign n1070 = ~b & n1069;
  assign n1071 = i0 & n1060;
  assign n1072 = k0 & n1071;
  assign n1073 = ~g0 & n1072;
  assign n1074 = ~y & n1073;
  assign n1075 = ~b & n1074;
  assign n1076 = i0 & n1066;
  assign n1077 = k0 & n1076;
  assign n1078 = ~y & n1077;
  assign n1079 = ~b & n1078;
  assign n1080 = ~i0 & n1060;
  assign n1081 = j0 & n1080;
  assign n1082 = k0 & n1081;
  assign n1083 = ~g0 & n1082;
  assign n1084 = ~b & n1083;
  assign n1085 = ~i0 & n1066;
  assign n1086 = j0 & n1085;
  assign n1087 = k0 & n1086;
  assign n1088 = ~b & n1087;
  assign n1089 = ~q & n324;
  assign n1090 = ~x & n1089;
  assign n1091 = ~b0 & n1090;
  assign n1092 = ~c0 & n1091;
  assign n1093 = d0 & n1092;
  assign n1094 = k0 & n1093;
  assign n1095 = ~g0 & n1094;
  assign n1096 = ~v & n1095;
  assign n1097 = ~y & n1096;
  assign n1098 = ~a0 & n1097;
  assign n1099 = ~o & n1098;
  assign n1100 = ~m & n1099;
  assign n1101 = ~q & n385;
  assign n1102 = ~x & n1101;
  assign n1103 = ~b0 & n1102;
  assign n1104 = ~c0 & n1103;
  assign n1105 = d0 & n1104;
  assign n1106 = k0 & n1105;
  assign n1107 = ~v & n1106;
  assign n1108 = ~y & n1107;
  assign n1109 = ~a0 & n1108;
  assign n1110 = ~o & n1109;
  assign n1111 = ~m & n1110;
  assign n1112 = ~x & n979;
  assign n1113 = ~b0 & n1112;
  assign n1114 = ~c0 & n1113;
  assign n1115 = ~d0 & n1114;
  assign n1116 = k0 & n1115;
  assign n1117 = ~g0 & n1116;
  assign n1118 = ~y & n1117;
  assign n1119 = ~a0 & n1118;
  assign n1120 = ~o & n1119;
  assign n1121 = ~m & n1120;
  assign n1122 = ~x & n991;
  assign n1123 = ~b0 & n1122;
  assign n1124 = ~c0 & n1123;
  assign n1125 = ~d0 & n1124;
  assign n1126 = k0 & n1125;
  assign n1127 = ~y & n1126;
  assign n1128 = ~a0 & n1127;
  assign n1129 = ~o & n1128;
  assign n1130 = ~m & n1129;
  assign n1131 = i0 & n1115;
  assign n1132 = k0 & n1131;
  assign n1133 = ~g0 & n1132;
  assign n1134 = ~y & n1133;
  assign n1135 = ~o & n1134;
  assign n1136 = ~m & n1135;
  assign n1137 = i0 & n1125;
  assign n1138 = k0 & n1137;
  assign n1139 = ~y & n1138;
  assign n1140 = ~o & n1139;
  assign n1141 = ~m & n1140;
  assign n1142 = ~i0 & n1115;
  assign n1143 = j0 & n1142;
  assign n1144 = k0 & n1143;
  assign n1145 = ~g0 & n1144;
  assign n1146 = ~o & n1145;
  assign n1147 = ~m & n1146;
  assign n1148 = ~i0 & n1125;
  assign n1149 = j0 & n1148;
  assign n1150 = k0 & n1149;
  assign n1151 = ~o & n1150;
  assign n1152 = ~m & n1151;
  assign n1153 = ~n & n324;
  assign n1154 = ~q & n1153;
  assign n1155 = ~x & n1154;
  assign n1156 = ~b0 & n1155;
  assign n1157 = ~c0 & n1156;
  assign n1158 = d0 & n1157;
  assign n1159 = k0 & n1158;
  assign n1160 = ~g0 & n1159;
  assign n1161 = ~v & n1160;
  assign n1162 = ~y & n1161;
  assign n1163 = ~a0 & n1162;
  assign n1164 = ~m & n1163;
  assign n1165 = ~n & n385;
  assign n1166 = ~q & n1165;
  assign n1167 = ~x & n1166;
  assign n1168 = ~b0 & n1167;
  assign n1169 = ~c0 & n1168;
  assign n1170 = d0 & n1169;
  assign n1171 = k0 & n1170;
  assign n1172 = ~v & n1171;
  assign n1173 = ~y & n1172;
  assign n1174 = ~a0 & n1173;
  assign n1175 = ~m & n1174;
  assign n1176 = ~x & n1038;
  assign n1177 = ~b0 & n1176;
  assign n1178 = ~c0 & n1177;
  assign n1179 = ~d0 & n1178;
  assign n1180 = k0 & n1179;
  assign n1181 = ~g0 & n1180;
  assign n1182 = ~y & n1181;
  assign n1183 = ~a0 & n1182;
  assign n1184 = ~m & n1183;
  assign n1185 = ~x & n1050;
  assign n1186 = ~b0 & n1185;
  assign n1187 = ~c0 & n1186;
  assign n1188 = ~d0 & n1187;
  assign n1189 = k0 & n1188;
  assign n1190 = ~y & n1189;
  assign n1191 = ~a0 & n1190;
  assign n1192 = ~m & n1191;
  assign n1193 = i0 & n1179;
  assign n1194 = k0 & n1193;
  assign n1195 = ~g0 & n1194;
  assign n1196 = ~y & n1195;
  assign n1197 = ~m & n1196;
  assign n1198 = i0 & n1188;
  assign n1199 = k0 & n1198;
  assign n1200 = ~y & n1199;
  assign n1201 = ~m & n1200;
  assign n1202 = ~i0 & n1179;
  assign n1203 = j0 & n1202;
  assign n1204 = k0 & n1203;
  assign n1205 = ~g0 & n1204;
  assign n1206 = ~m & n1205;
  assign n1207 = ~i0 & n1188;
  assign n1208 = j0 & n1207;
  assign n1209 = k0 & n1208;
  assign n1210 = ~m & n1209;
  assign n1211 = ~c & ~q;
  assign n1212 = ~r & n1211;
  assign n1213 = ~x & n1212;
  assign n1214 = ~b0 & n1213;
  assign n1215 = ~c0 & n1214;
  assign n1216 = ~j0 & n1215;
  assign n1217 = k0 & n1216;
  assign n1218 = ~g0 & n1217;
  assign n1219 = ~v & n1218;
  assign n1220 = ~y & n1219;
  assign n1221 = ~a0 & n1220;
  assign n1222 = ~o & n1221;
  assign n1223 = ~f0 & n1222;
  assign n1224 = ~e0 & n1223;
  assign n1225 = ~c & ~i;
  assign n1226 = ~q & n1225;
  assign n1227 = ~r & n1226;
  assign n1228 = ~x & n1227;
  assign n1229 = ~b0 & n1228;
  assign n1230 = ~c0 & n1229;
  assign n1231 = ~j0 & n1230;
  assign n1232 = k0 & n1231;
  assign n1233 = ~v & n1232;
  assign n1234 = ~y & n1233;
  assign n1235 = ~a0 & n1234;
  assign n1236 = ~o & n1235;
  assign n1237 = ~f0 & n1236;
  assign n1238 = ~e0 & n1237;
  assign n1239 = ~c & ~n;
  assign n1240 = ~q & n1239;
  assign n1241 = ~r & n1240;
  assign n1242 = ~x & n1241;
  assign n1243 = ~b0 & n1242;
  assign n1244 = ~c0 & n1243;
  assign n1245 = ~j0 & n1244;
  assign n1246 = k0 & n1245;
  assign n1247 = ~g0 & n1246;
  assign n1248 = ~v & n1247;
  assign n1249 = ~y & n1248;
  assign n1250 = ~a0 & n1249;
  assign n1251 = ~f0 & n1250;
  assign n1252 = ~e0 & n1251;
  assign n1253 = ~n & n1225;
  assign n1254 = ~q & n1253;
  assign n1255 = ~r & n1254;
  assign n1256 = ~x & n1255;
  assign n1257 = ~b0 & n1256;
  assign n1258 = ~c0 & n1257;
  assign n1259 = ~j0 & n1258;
  assign n1260 = k0 & n1259;
  assign n1261 = ~v & n1260;
  assign n1262 = ~y & n1261;
  assign n1263 = ~a0 & n1262;
  assign n1264 = ~f0 & n1263;
  assign n1265 = ~e0 & n1264;
  assign n1266 = ~q & ~x;
  assign n1267 = ~b0 & n1266;
  assign n1268 = ~c0 & n1267;
  assign n1269 = ~j0 & n1268;
  assign n1270 = k0 & n1269;
  assign n1271 = ~g0 & n1270;
  assign n1272 = ~v & n1271;
  assign n1273 = ~y & n1272;
  assign n1274 = ~a0 & n1273;
  assign n1275 = ~o & n1274;
  assign n1276 = ~f0 & n1275;
  assign n1277 = ~m & n1276;
  assign n1278 = ~e0 & n1277;
  assign n1279 = ~i & ~q;
  assign n1280 = ~x & n1279;
  assign n1281 = ~b0 & n1280;
  assign n1282 = ~c0 & n1281;
  assign n1283 = ~j0 & n1282;
  assign n1284 = k0 & n1283;
  assign n1285 = ~v & n1284;
  assign n1286 = ~y & n1285;
  assign n1287 = ~a0 & n1286;
  assign n1288 = ~o & n1287;
  assign n1289 = ~f0 & n1288;
  assign n1290 = ~m & n1289;
  assign n1291 = ~e0 & n1290;
  assign n1292 = ~d0 & n1282;
  assign n1293 = ~j0 & n1292;
  assign n1294 = k0 & n1293;
  assign n1295 = ~y & n1294;
  assign n1296 = ~a0 & n1295;
  assign n1297 = ~o & n1296;
  assign n1298 = ~f0 & n1297;
  assign n1299 = ~m & n1298;
  assign n1300 = ~e0 & n1299;
  assign n1301 = i0 & n1292;
  assign n1302 = ~j0 & n1301;
  assign n1303 = k0 & n1302;
  assign n1304 = ~y & n1303;
  assign n1305 = ~o & n1304;
  assign n1306 = ~f0 & n1305;
  assign n1307 = ~m & n1306;
  assign n1308 = ~e0 & n1307;
  assign n1309 = ~x & n42;
  assign n1310 = ~b0 & n1309;
  assign n1311 = ~c0 & n1310;
  assign n1312 = ~j0 & n1311;
  assign n1313 = k0 & n1312;
  assign n1314 = ~g0 & n1313;
  assign n1315 = ~v & n1314;
  assign n1316 = ~y & n1315;
  assign n1317 = ~a0 & n1316;
  assign n1318 = ~f0 & n1317;
  assign n1319 = ~m & n1318;
  assign n1320 = ~e0 & n1319;
  assign n1321 = ~i & ~n;
  assign n1322 = ~q & n1321;
  assign n1323 = ~x & n1322;
  assign n1324 = ~b0 & n1323;
  assign n1325 = ~c0 & n1324;
  assign n1326 = ~j0 & n1325;
  assign n1327 = k0 & n1326;
  assign n1328 = ~v & n1327;
  assign n1329 = ~y & n1328;
  assign n1330 = ~a0 & n1329;
  assign n1331 = ~f0 & n1330;
  assign n1332 = ~m & n1331;
  assign n1333 = ~e0 & n1332;
  assign n1334 = ~d0 & n1325;
  assign n1335 = ~j0 & n1334;
  assign n1336 = k0 & n1335;
  assign n1337 = ~y & n1336;
  assign n1338 = ~a0 & n1337;
  assign n1339 = ~f0 & n1338;
  assign n1340 = ~m & n1339;
  assign n1341 = ~e0 & n1340;
  assign n1342 = i0 & n1334;
  assign n1343 = ~j0 & n1342;
  assign n1344 = k0 & n1343;
  assign n1345 = ~y & n1344;
  assign n1346 = ~f0 & n1345;
  assign n1347 = ~m & n1346;
  assign n1348 = ~e0 & n1347;
  assign n1349 = ~r & n1279;
  assign n1350 = ~x & n1349;
  assign n1351 = ~b0 & n1350;
  assign n1352 = ~c0 & n1351;
  assign n1353 = ~d0 & n1352;
  assign n1354 = ~j0 & n1353;
  assign n1355 = k0 & n1354;
  assign n1356 = ~y & n1355;
  assign n1357 = ~a0 & n1356;
  assign n1358 = ~o & n1357;
  assign n1359 = ~f0 & n1358;
  assign n1360 = ~e0 & n1359;
  assign n1361 = i0 & n1353;
  assign n1362 = ~j0 & n1361;
  assign n1363 = k0 & n1362;
  assign n1364 = ~y & n1363;
  assign n1365 = ~o & n1364;
  assign n1366 = ~f0 & n1365;
  assign n1367 = ~e0 & n1366;
  assign n1368 = ~r & n1322;
  assign n1369 = ~x & n1368;
  assign n1370 = ~b0 & n1369;
  assign n1371 = ~c0 & n1370;
  assign n1372 = ~d0 & n1371;
  assign n1373 = ~j0 & n1372;
  assign n1374 = k0 & n1373;
  assign n1375 = ~y & n1374;
  assign n1376 = ~a0 & n1375;
  assign n1377 = ~f0 & n1376;
  assign n1378 = ~e0 & n1377;
  assign n1379 = i0 & n1372;
  assign n1380 = ~j0 & n1379;
  assign n1381 = k0 & n1380;
  assign n1382 = ~y & n1381;
  assign n1383 = ~f0 & n1382;
  assign n1384 = ~e0 & n1383;
  assign n1385 = ~c & ~h;
  assign n1386 = ~q & n1385;
  assign n1387 = ~r & n1386;
  assign n1388 = ~x & n1387;
  assign n1389 = ~b0 & n1388;
  assign n1390 = ~c0 & n1389;
  assign n1391 = k0 & n1390;
  assign n1392 = ~g0 & n1391;
  assign n1393 = ~v & n1392;
  assign n1394 = ~y & n1393;
  assign n1395 = ~a0 & n1394;
  assign n1396 = ~o & n1395;
  assign n1397 = ~e0 & n1396;
  assign n1398 = ~i & n1385;
  assign n1399 = ~q & n1398;
  assign n1400 = ~r & n1399;
  assign n1401 = ~x & n1400;
  assign n1402 = ~b0 & n1401;
  assign n1403 = ~c0 & n1402;
  assign n1404 = k0 & n1403;
  assign n1405 = ~v & n1404;
  assign n1406 = ~y & n1405;
  assign n1407 = ~a0 & n1406;
  assign n1408 = ~o & n1407;
  assign n1409 = ~e0 & n1408;
  assign n1410 = ~n & n1385;
  assign n1411 = ~q & n1410;
  assign n1412 = ~r & n1411;
  assign n1413 = ~x & n1412;
  assign n1414 = ~b0 & n1413;
  assign n1415 = ~c0 & n1414;
  assign n1416 = k0 & n1415;
  assign n1417 = ~g0 & n1416;
  assign n1418 = ~v & n1417;
  assign n1419 = ~y & n1418;
  assign n1420 = ~a0 & n1419;
  assign n1421 = ~e0 & n1420;
  assign n1422 = ~n & n1398;
  assign n1423 = ~q & n1422;
  assign n1424 = ~r & n1423;
  assign n1425 = ~x & n1424;
  assign n1426 = ~b0 & n1425;
  assign n1427 = ~c0 & n1426;
  assign n1428 = k0 & n1427;
  assign n1429 = ~v & n1428;
  assign n1430 = ~y & n1429;
  assign n1431 = ~a0 & n1430;
  assign n1432 = ~e0 & n1431;
  assign n1433 = h & ~n;
  assign n1434 = ~q & n1433;
  assign n1435 = ~x & n1434;
  assign n1436 = ~b0 & n1435;
  assign n1437 = ~c0 & n1436;
  assign n1438 = i0 & n1437;
  assign n1439 = d & n1438;
  assign n1440 = ~s & n1439;
  assign n1441 = v & n1440;
  assign n1442 = ~y & n1441;
  assign n1443 = k & n1442;
  assign n1444 = f0 & n1443;
  assign n1445 = ~m & n1444;
  assign n1446 = h & ~l;
  assign n1447 = ~n & n1446;
  assign n1448 = ~q & n1447;
  assign n1449 = ~t & n1448;
  assign n1450 = ~x & n1449;
  assign n1451 = ~b0 & n1450;
  assign n1452 = ~c0 & n1451;
  assign n1453 = i0 & n1452;
  assign n1454 = v & n1453;
  assign n1455 = ~y & n1454;
  assign n1456 = k & n1455;
  assign n1457 = f0 & n1456;
  assign n1458 = ~m & n1457;
  assign n1459 = ~d0 & n1437;
  assign n1460 = i0 & n1459;
  assign n1461 = d & n1460;
  assign n1462 = ~s & n1461;
  assign n1463 = ~y & n1462;
  assign n1464 = k & n1463;
  assign n1465 = f0 & n1464;
  assign n1466 = ~m & n1465;
  assign n1467 = ~d0 & n1452;
  assign n1468 = i0 & n1467;
  assign n1469 = ~y & n1468;
  assign n1470 = k & n1469;
  assign n1471 = f0 & n1470;
  assign n1472 = ~m & n1471;
  assign n1473 = ~i0 & n1437;
  assign n1474 = j0 & n1473;
  assign n1475 = d & n1474;
  assign n1476 = ~s & n1475;
  assign n1477 = v & n1476;
  assign n1478 = k & n1477;
  assign n1479 = f0 & n1478;
  assign n1480 = ~m & n1479;
  assign n1481 = ~i0 & n1452;
  assign n1482 = j0 & n1481;
  assign n1483 = v & n1482;
  assign n1484 = k & n1483;
  assign n1485 = f0 & n1484;
  assign n1486 = ~m & n1485;
  assign n1487 = ~i0 & n1459;
  assign n1488 = j0 & n1487;
  assign n1489 = d & n1488;
  assign n1490 = ~s & n1489;
  assign n1491 = k & n1490;
  assign n1492 = f0 & n1491;
  assign n1493 = ~m & n1492;
  assign n1494 = ~i0 & n1467;
  assign n1495 = j0 & n1494;
  assign n1496 = k & n1495;
  assign n1497 = f0 & n1496;
  assign n1498 = ~m & n1497;
  assign n1499 = ~r & n1434;
  assign n1500 = ~x & n1499;
  assign n1501 = ~b0 & n1500;
  assign n1502 = ~c0 & n1501;
  assign n1503 = i0 & n1502;
  assign n1504 = d & n1503;
  assign n1505 = ~s & n1504;
  assign n1506 = v & n1505;
  assign n1507 = ~y & n1506;
  assign n1508 = k & n1507;
  assign n1509 = f0 & n1508;
  assign n1510 = ~r & n1448;
  assign n1511 = ~t & n1510;
  assign n1512 = ~x & n1511;
  assign n1513 = ~b0 & n1512;
  assign n1514 = ~c0 & n1513;
  assign n1515 = i0 & n1514;
  assign n1516 = v & n1515;
  assign n1517 = ~y & n1516;
  assign n1518 = k & n1517;
  assign n1519 = f0 & n1518;
  assign n1520 = ~d0 & n1502;
  assign n1521 = i0 & n1520;
  assign n1522 = d & n1521;
  assign n1523 = ~s & n1522;
  assign n1524 = ~y & n1523;
  assign n1525 = k & n1524;
  assign n1526 = f0 & n1525;
  assign n1527 = ~d0 & n1514;
  assign n1528 = i0 & n1527;
  assign n1529 = ~y & n1528;
  assign n1530 = k & n1529;
  assign n1531 = f0 & n1530;
  assign n1532 = ~i0 & n1502;
  assign n1533 = j0 & n1532;
  assign n1534 = d & n1533;
  assign n1535 = ~s & n1534;
  assign n1536 = v & n1535;
  assign n1537 = k & n1536;
  assign n1538 = f0 & n1537;
  assign n1539 = ~i0 & n1514;
  assign n1540 = j0 & n1539;
  assign n1541 = v & n1540;
  assign n1542 = k & n1541;
  assign n1543 = f0 & n1542;
  assign n1544 = ~i0 & n1520;
  assign n1545 = j0 & n1544;
  assign n1546 = d & n1545;
  assign n1547 = ~s & n1546;
  assign n1548 = k & n1547;
  assign n1549 = f0 & n1548;
  assign n1550 = ~i0 & n1527;
  assign n1551 = j0 & n1550;
  assign n1552 = k & n1551;
  assign n1553 = f0 & n1552;
  assign n1554 = c & ~j;
  assign n1555 = ~n & n1554;
  assign n1556 = ~q & n1555;
  assign n1557 = ~r & n1556;
  assign n1558 = ~x & n1557;
  assign n1559 = ~b0 & n1558;
  assign n1560 = ~c0 & n1559;
  assign n1561 = d0 & n1560;
  assign n1562 = d & n1561;
  assign n1563 = ~s & n1562;
  assign n1564 = ~v & n1563;
  assign n1565 = ~y & n1564;
  assign n1566 = ~a0 & n1565;
  assign n1567 = ~l & n1554;
  assign n1568 = ~n & n1567;
  assign n1569 = ~q & n1568;
  assign n1570 = ~r & n1569;
  assign n1571 = ~t & n1570;
  assign n1572 = ~x & n1571;
  assign n1573 = ~b0 & n1572;
  assign n1574 = ~c0 & n1573;
  assign n1575 = d0 & n1574;
  assign n1576 = ~v & n1575;
  assign n1577 = ~y & n1576;
  assign n1578 = ~a0 & n1577;
  assign n1579 = ~h & ~q;
  assign n1580 = ~x & n1579;
  assign n1581 = ~b0 & n1580;
  assign n1582 = ~c0 & n1581;
  assign n1583 = k0 & n1582;
  assign n1584 = ~g0 & n1583;
  assign n1585 = ~v & n1584;
  assign n1586 = ~y & n1585;
  assign n1587 = ~a0 & n1586;
  assign n1588 = ~o & n1587;
  assign n1589 = ~m & n1588;
  assign n1590 = ~e0 & n1589;
  assign n1591 = ~h & ~i;
  assign n1592 = ~q & n1591;
  assign n1593 = ~x & n1592;
  assign n1594 = ~b0 & n1593;
  assign n1595 = ~c0 & n1594;
  assign n1596 = k0 & n1595;
  assign n1597 = ~v & n1596;
  assign n1598 = ~y & n1597;
  assign n1599 = ~a0 & n1598;
  assign n1600 = ~o & n1599;
  assign n1601 = ~m & n1600;
  assign n1602 = ~e0 & n1601;
  assign n1603 = ~d0 & n1582;
  assign n1604 = k0 & n1603;
  assign n1605 = ~g0 & n1604;
  assign n1606 = ~y & n1605;
  assign n1607 = ~a0 & n1606;
  assign n1608 = ~o & n1607;
  assign n1609 = ~m & n1608;
  assign n1610 = ~e0 & n1609;
  assign n1611 = ~d0 & n1595;
  assign n1612 = k0 & n1611;
  assign n1613 = ~y & n1612;
  assign n1614 = ~a0 & n1613;
  assign n1615 = ~o & n1614;
  assign n1616 = ~m & n1615;
  assign n1617 = ~e0 & n1616;
  assign n1618 = i0 & n1603;
  assign n1619 = k0 & n1618;
  assign n1620 = ~g0 & n1619;
  assign n1621 = ~y & n1620;
  assign n1622 = ~o & n1621;
  assign n1623 = ~m & n1622;
  assign n1624 = ~e0 & n1623;
  assign n1625 = i0 & n1611;
  assign n1626 = k0 & n1625;
  assign n1627 = ~y & n1626;
  assign n1628 = ~o & n1627;
  assign n1629 = ~m & n1628;
  assign n1630 = ~e0 & n1629;
  assign n1631 = ~i0 & n1603;
  assign n1632 = j0 & n1631;
  assign n1633 = k0 & n1632;
  assign n1634 = ~g0 & n1633;
  assign n1635 = ~o & n1634;
  assign n1636 = ~m & n1635;
  assign n1637 = ~e0 & n1636;
  assign n1638 = ~i0 & n1611;
  assign n1639 = j0 & n1638;
  assign n1640 = k0 & n1639;
  assign n1641 = ~o & n1640;
  assign n1642 = ~m & n1641;
  assign n1643 = ~e0 & n1642;
  assign n1644 = ~h & ~n;
  assign n1645 = ~q & n1644;
  assign n1646 = ~x & n1645;
  assign n1647 = ~b0 & n1646;
  assign n1648 = ~c0 & n1647;
  assign n1649 = k0 & n1648;
  assign n1650 = ~g0 & n1649;
  assign n1651 = ~v & n1650;
  assign n1652 = ~y & n1651;
  assign n1653 = ~a0 & n1652;
  assign n1654 = ~m & n1653;
  assign n1655 = ~e0 & n1654;
  assign n1656 = ~n & n1591;
  assign n1657 = ~q & n1656;
  assign n1658 = ~x & n1657;
  assign n1659 = ~b0 & n1658;
  assign n1660 = ~c0 & n1659;
  assign n1661 = k0 & n1660;
  assign n1662 = ~v & n1661;
  assign n1663 = ~y & n1662;
  assign n1664 = ~a0 & n1663;
  assign n1665 = ~m & n1664;
  assign n1666 = ~e0 & n1665;
  assign n1667 = ~d0 & n1648;
  assign n1668 = k0 & n1667;
  assign n1669 = ~g0 & n1668;
  assign n1670 = ~y & n1669;
  assign n1671 = ~a0 & n1670;
  assign n1672 = ~m & n1671;
  assign n1673 = ~e0 & n1672;
  assign n1674 = ~d0 & n1660;
  assign n1675 = k0 & n1674;
  assign n1676 = ~y & n1675;
  assign n1677 = ~a0 & n1676;
  assign n1678 = ~m & n1677;
  assign n1679 = ~e0 & n1678;
  assign n1680 = i0 & n1667;
  assign n1681 = k0 & n1680;
  assign n1682 = ~g0 & n1681;
  assign n1683 = ~y & n1682;
  assign n1684 = ~m & n1683;
  assign n1685 = ~e0 & n1684;
  assign n1686 = i0 & n1674;
  assign n1687 = k0 & n1686;
  assign n1688 = ~y & n1687;
  assign n1689 = ~m & n1688;
  assign n1690 = ~e0 & n1689;
  assign n1691 = ~i0 & n1667;
  assign n1692 = j0 & n1691;
  assign n1693 = k0 & n1692;
  assign n1694 = ~g0 & n1693;
  assign n1695 = ~m & n1694;
  assign n1696 = ~e0 & n1695;
  assign n1697 = ~i0 & n1674;
  assign n1698 = j0 & n1697;
  assign n1699 = k0 & n1698;
  assign n1700 = ~m & n1699;
  assign n1701 = ~e0 & n1700;
  assign n1702 = ~r & n1579;
  assign n1703 = ~x & n1702;
  assign n1704 = ~b0 & n1703;
  assign n1705 = ~c0 & n1704;
  assign n1706 = ~d0 & n1705;
  assign n1707 = k0 & n1706;
  assign n1708 = ~g0 & n1707;
  assign n1709 = ~y & n1708;
  assign n1710 = ~a0 & n1709;
  assign n1711 = ~o & n1710;
  assign n1712 = ~e0 & n1711;
  assign n1713 = ~r & n1592;
  assign n1714 = ~x & n1713;
  assign n1715 = ~b0 & n1714;
  assign n1716 = ~c0 & n1715;
  assign n1717 = ~d0 & n1716;
  assign n1718 = k0 & n1717;
  assign n1719 = ~y & n1718;
  assign n1720 = ~a0 & n1719;
  assign n1721 = ~o & n1720;
  assign n1722 = ~e0 & n1721;
  assign n1723 = i0 & n1706;
  assign n1724 = k0 & n1723;
  assign n1725 = ~g0 & n1724;
  assign n1726 = ~y & n1725;
  assign n1727 = ~o & n1726;
  assign n1728 = ~e0 & n1727;
  assign n1729 = i0 & n1717;
  assign n1730 = k0 & n1729;
  assign n1731 = ~y & n1730;
  assign n1732 = ~o & n1731;
  assign n1733 = ~e0 & n1732;
  assign n1734 = ~i0 & n1706;
  assign n1735 = j0 & n1734;
  assign n1736 = k0 & n1735;
  assign n1737 = ~g0 & n1736;
  assign n1738 = ~o & n1737;
  assign n1739 = ~e0 & n1738;
  assign n1740 = ~i0 & n1717;
  assign n1741 = j0 & n1740;
  assign n1742 = k0 & n1741;
  assign n1743 = ~o & n1742;
  assign n1744 = ~e0 & n1743;
  assign n1745 = ~r & n1645;
  assign n1746 = ~x & n1745;
  assign n1747 = ~b0 & n1746;
  assign n1748 = ~c0 & n1747;
  assign n1749 = ~d0 & n1748;
  assign n1750 = k0 & n1749;
  assign n1751 = ~g0 & n1750;
  assign n1752 = ~y & n1751;
  assign n1753 = ~a0 & n1752;
  assign n1754 = ~e0 & n1753;
  assign n1755 = ~r & n1657;
  assign n1756 = ~x & n1755;
  assign n1757 = ~b0 & n1756;
  assign n1758 = ~c0 & n1757;
  assign n1759 = ~d0 & n1758;
  assign n1760 = k0 & n1759;
  assign n1761 = ~y & n1760;
  assign n1762 = ~a0 & n1761;
  assign n1763 = ~e0 & n1762;
  assign n1764 = i0 & n1749;
  assign n1765 = k0 & n1764;
  assign n1766 = ~g0 & n1765;
  assign n1767 = ~y & n1766;
  assign n1768 = ~e0 & n1767;
  assign n1769 = i0 & n1759;
  assign n1770 = k0 & n1769;
  assign n1771 = ~y & n1770;
  assign n1772 = ~e0 & n1771;
  assign n1773 = ~i0 & n1749;
  assign n1774 = j0 & n1773;
  assign n1775 = k0 & n1774;
  assign n1776 = ~g0 & n1775;
  assign n1777 = ~e0 & n1776;
  assign n1778 = ~i0 & n1759;
  assign n1779 = j0 & n1778;
  assign n1780 = k0 & n1779;
  assign n1781 = ~e0 & n1780;
  assign n1782 = h & n;
  assign n1783 = ~q & n1782;
  assign n1784 = ~x & n1783;
  assign n1785 = ~b0 & n1784;
  assign n1786 = ~c0 & n1785;
  assign n1787 = i0 & n1786;
  assign n1788 = v & n1787;
  assign n1789 = ~y & n1788;
  assign n1790 = ~o & n1789;
  assign n1791 = k & n1790;
  assign n1792 = f0 & n1791;
  assign n1793 = ~m & n1792;
  assign n1794 = ~d0 & n1786;
  assign n1795 = i0 & n1794;
  assign n1796 = ~y & n1795;
  assign n1797 = ~o & n1796;
  assign n1798 = k & n1797;
  assign n1799 = f0 & n1798;
  assign n1800 = ~m & n1799;
  assign n1801 = ~i0 & n1786;
  assign n1802 = j0 & n1801;
  assign n1803 = v & n1802;
  assign n1804 = ~o & n1803;
  assign n1805 = k & n1804;
  assign n1806 = f0 & n1805;
  assign n1807 = ~m & n1806;
  assign n1808 = ~i0 & n1794;
  assign n1809 = j0 & n1808;
  assign n1810 = ~o & n1809;
  assign n1811 = k & n1810;
  assign n1812 = f0 & n1811;
  assign n1813 = ~m & n1812;
  assign n1814 = d & n1437;
  assign n1815 = ~s & n1814;
  assign n1816 = ~y & n1815;
  assign n1817 = ~a0 & n1816;
  assign n1818 = k & n1817;
  assign n1819 = f0 & n1818;
  assign n1820 = ~m & n1819;
  assign n1821 = ~y & n1452;
  assign n1822 = ~a0 & n1821;
  assign n1823 = k & n1822;
  assign n1824 = f0 & n1823;
  assign n1825 = ~m & n1824;
  assign n1826 = ~r & n1783;
  assign n1827 = ~x & n1826;
  assign n1828 = ~b0 & n1827;
  assign n1829 = ~c0 & n1828;
  assign n1830 = i0 & n1829;
  assign n1831 = v & n1830;
  assign n1832 = ~y & n1831;
  assign n1833 = ~o & n1832;
  assign n1834 = k & n1833;
  assign n1835 = f0 & n1834;
  assign n1836 = ~d0 & n1829;
  assign n1837 = i0 & n1836;
  assign n1838 = ~y & n1837;
  assign n1839 = ~o & n1838;
  assign n1840 = k & n1839;
  assign n1841 = f0 & n1840;
  assign n1842 = ~i0 & n1829;
  assign n1843 = j0 & n1842;
  assign n1844 = v & n1843;
  assign n1845 = ~o & n1844;
  assign n1846 = k & n1845;
  assign n1847 = f0 & n1846;
  assign n1848 = ~i0 & n1836;
  assign n1849 = j0 & n1848;
  assign n1850 = ~o & n1849;
  assign n1851 = k & n1850;
  assign n1852 = f0 & n1851;
  assign n1853 = d & n1502;
  assign n1854 = ~s & n1853;
  assign n1855 = ~y & n1854;
  assign n1856 = ~a0 & n1855;
  assign n1857 = k & n1856;
  assign n1858 = f0 & n1857;
  assign n1859 = ~y & n1514;
  assign n1860 = ~a0 & n1859;
  assign n1861 = k & n1860;
  assign n1862 = f0 & n1861;
  assign n1863 = ~v & n1561;
  assign n1864 = ~y & n1863;
  assign n1865 = ~a0 & n1864;
  assign n1866 = ~k & n1865;
  assign n1867 = n & n1554;
  assign n1868 = ~q & n1867;
  assign n1869 = ~r & n1868;
  assign n1870 = ~x & n1869;
  assign n1871 = ~b0 & n1870;
  assign n1872 = ~c0 & n1871;
  assign n1873 = d0 & n1872;
  assign n1874 = ~v & n1873;
  assign n1875 = ~y & n1874;
  assign n1876 = ~a0 & n1875;
  assign n1877 = ~o & n1876;
  assign n1878 = ~y & n1786;
  assign n1879 = ~a0 & n1878;
  assign n1880 = ~o & n1879;
  assign n1881 = k & n1880;
  assign n1882 = f0 & n1881;
  assign n1883 = ~m & n1882;
  assign n1884 = h & ~j;
  assign n1885 = ~q & n1884;
  assign n1886 = ~x & n1885;
  assign n1887 = ~b0 & n1886;
  assign n1888 = ~c0 & n1887;
  assign n1889 = i0 & n1888;
  assign n1890 = v & n1889;
  assign n1891 = ~y & n1890;
  assign n1892 = ~o & n1891;
  assign n1893 = f0 & n1892;
  assign n1894 = ~m & n1893;
  assign n1895 = ~d0 & n1888;
  assign n1896 = i0 & n1895;
  assign n1897 = ~y & n1896;
  assign n1898 = ~o & n1897;
  assign n1899 = f0 & n1898;
  assign n1900 = ~m & n1899;
  assign n1901 = ~i0 & n1888;
  assign n1902 = j0 & n1901;
  assign n1903 = v & n1902;
  assign n1904 = ~o & n1903;
  assign n1905 = f0 & n1904;
  assign n1906 = ~m & n1905;
  assign n1907 = ~i0 & n1895;
  assign n1908 = j0 & n1907;
  assign n1909 = ~o & n1908;
  assign n1910 = f0 & n1909;
  assign n1911 = ~m & n1910;
  assign n1912 = ~n & n1884;
  assign n1913 = ~q & n1912;
  assign n1914 = ~x & n1913;
  assign n1915 = ~b0 & n1914;
  assign n1916 = ~c0 & n1915;
  assign n1917 = i0 & n1916;
  assign n1918 = v & n1917;
  assign n1919 = ~y & n1918;
  assign n1920 = f0 & n1919;
  assign n1921 = ~m & n1920;
  assign n1922 = ~d0 & n1916;
  assign n1923 = i0 & n1922;
  assign n1924 = ~y & n1923;
  assign n1925 = f0 & n1924;
  assign n1926 = ~m & n1925;
  assign n1927 = ~i0 & n1916;
  assign n1928 = j0 & n1927;
  assign n1929 = v & n1928;
  assign n1930 = f0 & n1929;
  assign n1931 = ~m & n1930;
  assign n1932 = ~i0 & n1922;
  assign n1933 = j0 & n1932;
  assign n1934 = f0 & n1933;
  assign n1935 = ~m & n1934;
  assign n1936 = ~y & n1829;
  assign n1937 = ~a0 & n1936;
  assign n1938 = ~o & n1937;
  assign n1939 = k & n1938;
  assign n1940 = f0 & n1939;
  assign n1941 = ~r & n1885;
  assign n1942 = ~x & n1941;
  assign n1943 = ~b0 & n1942;
  assign n1944 = ~c0 & n1943;
  assign n1945 = i0 & n1944;
  assign n1946 = v & n1945;
  assign n1947 = ~y & n1946;
  assign n1948 = ~o & n1947;
  assign n1949 = f0 & n1948;
  assign n1950 = ~d0 & n1944;
  assign n1951 = i0 & n1950;
  assign n1952 = ~y & n1951;
  assign n1953 = ~o & n1952;
  assign n1954 = f0 & n1953;
  assign n1955 = ~i0 & n1944;
  assign n1956 = j0 & n1955;
  assign n1957 = v & n1956;
  assign n1958 = ~o & n1957;
  assign n1959 = f0 & n1958;
  assign n1960 = ~i0 & n1950;
  assign n1961 = j0 & n1960;
  assign n1962 = ~o & n1961;
  assign n1963 = f0 & n1962;
  assign n1964 = ~r & n1913;
  assign n1965 = ~x & n1964;
  assign n1966 = ~b0 & n1965;
  assign n1967 = ~c0 & n1966;
  assign n1968 = i0 & n1967;
  assign n1969 = v & n1968;
  assign n1970 = ~y & n1969;
  assign n1971 = f0 & n1970;
  assign n1972 = ~d0 & n1967;
  assign n1973 = i0 & n1972;
  assign n1974 = ~y & n1973;
  assign n1975 = f0 & n1974;
  assign n1976 = ~i0 & n1967;
  assign n1977 = j0 & n1976;
  assign n1978 = v & n1977;
  assign n1979 = f0 & n1978;
  assign n1980 = ~i0 & n1972;
  assign n1981 = j0 & n1980;
  assign n1982 = f0 & n1981;
  assign n1983 = d0 & n1268;
  assign n1984 = ~v & n1983;
  assign n1985 = ~y & n1984;
  assign n1986 = ~a0 & n1985;
  assign n1987 = ~o & n1986;
  assign n1988 = ~m & n1987;
  assign n1989 = a & n1988;
  assign n1990 = d0 & n1311;
  assign n1991 = ~v & n1990;
  assign n1992 = ~y & n1991;
  assign n1993 = ~a0 & n1992;
  assign n1994 = ~m & n1993;
  assign n1995 = a & n1994;
  assign n1996 = ~q & ~r;
  assign n1997 = ~x & n1996;
  assign n1998 = ~b0 & n1997;
  assign n1999 = ~c0 & n1998;
  assign n2000 = d0 & n1999;
  assign n2001 = ~v & n2000;
  assign n2002 = ~y & n2001;
  assign n2003 = ~a0 & n2002;
  assign n2004 = ~o & n2003;
  assign n2005 = a & n2004;
  assign n2006 = ~x & n43;
  assign n2007 = ~b0 & n2006;
  assign n2008 = ~c0 & n2007;
  assign n2009 = d0 & n2008;
  assign n2010 = ~v & n2009;
  assign n2011 = ~y & n2010;
  assign n2012 = ~a0 & n2011;
  assign n2013 = a & n2012;
  assign n2014 = i0 & n1268;
  assign n2015 = v & n2014;
  assign n2016 = ~y & n2015;
  assign n2017 = ~o & n2016;
  assign n2018 = ~m & n2017;
  assign n2019 = h0 & n2018;
  assign n2020 = z & n2019;
  assign n2021 = ~i0 & n1268;
  assign n2022 = j0 & n2021;
  assign n2023 = v & n2022;
  assign n2024 = ~o & n2023;
  assign n2025 = ~m & n2024;
  assign n2026 = h0 & n2025;
  assign n2027 = z & n2026;
  assign n2028 = i0 & n1999;
  assign n2029 = v & n2028;
  assign n2030 = ~y & n2029;
  assign n2031 = ~o & n2030;
  assign n2032 = h0 & n2031;
  assign n2033 = z & n2032;
  assign n2034 = ~i0 & n1999;
  assign n2035 = j0 & n2034;
  assign n2036 = v & n2035;
  assign n2037 = ~o & n2036;
  assign n2038 = h0 & n2037;
  assign n2039 = z & n2038;
  assign n2040 = i0 & n1311;
  assign n2041 = v & n2040;
  assign n2042 = ~y & n2041;
  assign n2043 = o & n2042;
  assign n2044 = ~m & n2043;
  assign n2045 = h0 & n2044;
  assign n2046 = ~i0 & n1311;
  assign n2047 = j0 & n2046;
  assign n2048 = v & n2047;
  assign n2049 = o & n2048;
  assign n2050 = ~m & n2049;
  assign n2051 = h0 & n2050;
  assign n2052 = i0 & n2008;
  assign n2053 = v & n2052;
  assign n2054 = ~y & n2053;
  assign n2055 = o & n2054;
  assign n2056 = h0 & n2055;
  assign n2057 = ~i0 & n2008;
  assign n2058 = j0 & n2057;
  assign n2059 = v & n2058;
  assign n2060 = o & n2059;
  assign n2061 = h0 & n2060;
  assign n2062 = i0 & n1983;
  assign n2063 = ~v & n2062;
  assign n2064 = ~y & n2063;
  assign n2065 = ~o & n2064;
  assign n2066 = ~m & n2065;
  assign n2067 = u & n2066;
  assign n2068 = ~i0 & n1983;
  assign n2069 = j0 & n2068;
  assign n2070 = ~v & n2069;
  assign n2071 = ~o & n2070;
  assign n2072 = ~m & n2071;
  assign n2073 = u & n2072;
  assign n2074 = i0 & n1990;
  assign n2075 = ~v & n2074;
  assign n2076 = ~y & n2075;
  assign n2077 = ~m & n2076;
  assign n2078 = u & n2077;
  assign n2079 = ~i0 & n1990;
  assign n2080 = j0 & n2079;
  assign n2081 = ~v & n2080;
  assign n2082 = ~m & n2081;
  assign n2083 = u & n2082;
  assign n2084 = i0 & n2000;
  assign n2085 = ~v & n2084;
  assign n2086 = ~y & n2085;
  assign n2087 = ~o & n2086;
  assign n2088 = u & n2087;
  assign n2089 = ~i0 & n2000;
  assign n2090 = j0 & n2089;
  assign n2091 = ~v & n2090;
  assign n2092 = ~o & n2091;
  assign n2093 = u & n2092;
  assign n2094 = i0 & n2009;
  assign n2095 = ~v & n2094;
  assign n2096 = ~y & n2095;
  assign n2097 = u & n2096;
  assign n2098 = ~i0 & n2009;
  assign n2099 = j0 & n2098;
  assign n2100 = ~v & n2099;
  assign n2101 = u & n2100;
  assign n2102 = ~y & n1888;
  assign n2103 = ~a0 & n2102;
  assign n2104 = ~o & n2103;
  assign n2105 = f0 & n2104;
  assign n2106 = ~m & n2105;
  assign n2107 = ~y & n1916;
  assign n2108 = ~a0 & n2107;
  assign n2109 = f0 & n2108;
  assign n2110 = ~m & n2109;
  assign n2111 = ~y & n1944;
  assign n2112 = ~a0 & n2111;
  assign n2113 = ~o & n2112;
  assign n2114 = f0 & n2113;
  assign n2115 = ~y & n1967;
  assign n2116 = ~a0 & n2115;
  assign n2117 = f0 & n2116;
  assign n2118 = ~i0 & ~c0;
  assign n2119 = ~g0 & n2118;
  assign n2120 = v & n2119;
  assign n2121 = ~y & n2120;
  assign n2122 = ~a0 & n2121;
  assign n2123 = ~f0 & n2122;
  assign n2124 = ~e0 & n2123;
  assign n2125 = h0 & n2124;
  assign n2126 = z & n2125;
  assign n2127 = ~x & ~c0;
  assign n2128 = i0 & n2127;
  assign n2129 = ~g0 & n2128;
  assign n2130 = v & n2129;
  assign n2131 = ~y & n2130;
  assign n2132 = ~f0 & n2131;
  assign n2133 = ~e0 & n2132;
  assign n2134 = h0 & n2133;
  assign n2135 = z & n2134;
  assign n2136 = o & n2122;
  assign n2137 = ~f0 & n2136;
  assign n2138 = ~e0 & n2137;
  assign n2139 = h0 & n2138;
  assign n2140 = ~c0 & ~d0;
  assign n2141 = ~i0 & n2140;
  assign n2142 = ~g0 & n2141;
  assign n2143 = ~y & n2142;
  assign n2144 = ~a0 & n2143;
  assign n2145 = o & n2144;
  assign n2146 = ~f0 & n2145;
  assign n2147 = ~e0 & n2146;
  assign n2148 = h0 & n2147;
  assign n2149 = o & n2131;
  assign n2150 = ~f0 & n2149;
  assign n2151 = ~e0 & n2150;
  assign n2152 = h0 & n2151;
  assign n2153 = ~y & n1311;
  assign n2154 = ~a0 & n2153;
  assign n2155 = o & n2154;
  assign n2156 = ~m & n2155;
  assign n2157 = h0 & n2156;
  assign n2158 = ~y & n2008;
  assign n2159 = ~a0 & n2158;
  assign n2160 = o & n2159;
  assign n2161 = h0 & n2160;
  assign n2162 = ~c0 & d0;
  assign n2163 = ~i0 & n2162;
  assign n2164 = ~g0 & n2163;
  assign n2165 = ~v & n2164;
  assign n2166 = ~y & n2165;
  assign n2167 = ~a0 & n2166;
  assign n2168 = ~f0 & n2167;
  assign n2169 = ~e0 & n2168;
  assign n2170 = u & n2169;
  assign n2171 = d0 & n2127;
  assign n2172 = i0 & n2171;
  assign n2173 = ~g0 & n2172;
  assign n2174 = ~v & n2173;
  assign n2175 = ~y & n2174;
  assign n2176 = ~f0 & n2175;
  assign n2177 = ~e0 & n2176;
  assign n2178 = u & n2177;
  assign n2179 = ~j0 & n2141;
  assign n2180 = k0 & n2179;
  assign n2181 = ~g0 & n2180;
  assign n2182 = ~y & n2181;
  assign n2183 = ~a0 & n2182;
  assign n2184 = ~f0 & n2183;
  assign n2185 = ~e0 & n2184;
  assign n2186 = ~d0 & n2127;
  assign n2187 = i0 & n2186;
  assign n2188 = ~j0 & n2187;
  assign n2189 = k0 & n2188;
  assign n2190 = ~g0 & n2189;
  assign n2191 = ~y & n2190;
  assign n2192 = ~f0 & n2191;
  assign n2193 = ~e0 & n2192;
  assign n2194 = ~h & ~x;
  assign n2195 = ~c0 & n2194;
  assign n2196 = ~d0 & n2195;
  assign n2197 = i0 & n2196;
  assign n2198 = k0 & n2197;
  assign n2199 = ~g0 & n2198;
  assign n2200 = ~y & n2199;
  assign n2201 = ~f0 & n2200;
  assign n2202 = ~e0 & n2201;
  assign n2203 = j0 & n2118;
  assign n2204 = ~g0 & n2203;
  assign n2205 = v & n2204;
  assign n2206 = ~f0 & n2205;
  assign n2207 = ~e0 & n2206;
  assign n2208 = h0 & n2207;
  assign n2209 = z & n2208;
  assign n2210 = o & n2205;
  assign n2211 = ~f0 & n2210;
  assign n2212 = ~e0 & n2211;
  assign n2213 = h0 & n2212;
  assign n2214 = j0 & n2163;
  assign n2215 = ~g0 & n2214;
  assign n2216 = ~v & n2215;
  assign n2217 = ~f0 & n2216;
  assign n2218 = ~e0 & n2217;
  assign n2219 = u & n2218;
  assign n2220 = ~h & ~c0;
  assign n2221 = ~d0 & n2220;
  assign n2222 = ~i0 & n2221;
  assign n2223 = j0 & n2222;
  assign n2224 = k0 & n2223;
  assign n2225 = ~g0 & n2224;
  assign n2226 = ~f0 & n2225;
  assign n2227 = ~e0 & n2226;
  assign n2228 = ~n295 & ~n305;
  assign n2229 = ~n284 & n2228;
  assign n2230 = ~n277 & n2229;
  assign n2231 = ~n270 & n2230;
  assign n2232 = ~n261 & n2231;
  assign n2233 = ~n252 & n2232;
  assign n2234 = ~n243 & n2233;
  assign n2235 = ~n234 & n2234;
  assign n2236 = ~n228 & n2235;
  assign n2237 = ~n222 & n2236;
  assign n2238 = ~n217 & n2237;
  assign n2239 = ~n212 & n2238;
  assign n2240 = ~n207 & n2239;
  assign n2241 = ~n202 & n2240;
  assign n2242 = ~n197 & n2241;
  assign n2243 = ~n192 & n2242;
  assign n2244 = ~n184 & n2243;
  assign n2245 = ~n175 & n2244;
  assign n2246 = ~n166 & n2245;
  assign n2247 = ~n158 & n2246;
  assign n2248 = ~n149 & n2247;
  assign n2249 = ~n139 & n2248;
  assign n2250 = ~n135 & n2249;
  assign n2251 = ~n131 & n2250;
  assign n2252 = ~n124 & n2251;
  assign n2253 = ~n115 & n2252;
  assign n2254 = ~n108 & n2253;
  assign n2255 = ~n101 & n2254;
  assign n2256 = ~n97 & n2255;
  assign n2257 = ~n88 & n2256;
  assign n2258 = ~n84 & n2257;
  assign n2259 = ~n75 & n2258;
  assign n2260 = ~n67 & n2259;
  assign n2261 = ~n58 & n2260;
  assign n2262 = ~n50 & n2261;
  assign n2263 = ~n2227 & n2262;
  assign n2264 = ~n2219 & n2263;
  assign n2265 = ~n2213 & n2264;
  assign n2266 = ~n2209 & n2265;
  assign n2267 = ~n2202 & n2266;
  assign n2268 = ~n2193 & n2267;
  assign n2269 = ~n2185 & n2268;
  assign n2270 = ~n2178 & n2269;
  assign n2271 = ~n2170 & n2270;
  assign n2272 = ~n2161 & n2271;
  assign n2273 = ~n2157 & n2272;
  assign n2274 = ~n2152 & n2273;
  assign n2275 = ~n2148 & n2274;
  assign n2276 = ~n2139 & n2275;
  assign n2277 = ~n2135 & n2276;
  assign n2278 = ~n2126 & n2277;
  assign n2279 = ~n2117 & n2278;
  assign n2280 = ~n2114 & n2279;
  assign n2281 = ~n2110 & n2280;
  assign n2282 = ~n2106 & n2281;
  assign n2283 = ~n2101 & n2282;
  assign n2284 = ~n2097 & n2283;
  assign n2285 = ~n2093 & n2284;
  assign n2286 = ~n2088 & n2285;
  assign n2287 = ~n2083 & n2286;
  assign n2288 = ~n2078 & n2287;
  assign n2289 = ~n2073 & n2288;
  assign n2290 = ~n2067 & n2289;
  assign n2291 = ~n2061 & n2290;
  assign n2292 = ~n2056 & n2291;
  assign n2293 = ~n2051 & n2292;
  assign n2294 = ~n2045 & n2293;
  assign n2295 = ~n2039 & n2294;
  assign n2296 = ~n2033 & n2295;
  assign n2297 = ~n2027 & n2296;
  assign n2298 = ~n2020 & n2297;
  assign n2299 = ~n2013 & n2298;
  assign n2300 = ~n2005 & n2299;
  assign n2301 = ~n1995 & n2300;
  assign n2302 = ~n1989 & n2301;
  assign n2303 = ~n1982 & n2302;
  assign n2304 = ~n1979 & n2303;
  assign n2305 = ~n1975 & n2304;
  assign n2306 = ~n1971 & n2305;
  assign n2307 = ~n1963 & n2306;
  assign n2308 = ~n1959 & n2307;
  assign n2309 = ~n1954 & n2308;
  assign n2310 = ~n1949 & n2309;
  assign n2311 = ~n1940 & n2310;
  assign n2312 = ~n1935 & n2311;
  assign n2313 = ~n1931 & n2312;
  assign n2314 = ~n1926 & n2313;
  assign n2315 = ~n1921 & n2314;
  assign n2316 = ~n1911 & n2315;
  assign n2317 = ~n1906 & n2316;
  assign n2318 = ~n1900 & n2317;
  assign n2319 = ~n1894 & n2318;
  assign n2320 = ~n1883 & n2319;
  assign n2321 = ~n1877 & n2320;
  assign n2322 = ~n1866 & n2321;
  assign n2323 = ~n1862 & n2322;
  assign n2324 = ~n1858 & n2323;
  assign n2325 = ~n1852 & n2324;
  assign n2326 = ~n1847 & n2325;
  assign n2327 = ~n1841 & n2326;
  assign n2328 = ~n1835 & n2327;
  assign n2329 = ~n1825 & n2328;
  assign n2330 = ~n1820 & n2329;
  assign n2331 = ~n1813 & n2330;
  assign n2332 = ~n1807 & n2331;
  assign n2333 = ~n1800 & n2332;
  assign n2334 = ~n1793 & n2333;
  assign n2335 = ~n1781 & n2334;
  assign n2336 = ~n1777 & n2335;
  assign n2337 = ~n1772 & n2336;
  assign n2338 = ~n1768 & n2337;
  assign n2339 = ~n1763 & n2338;
  assign n2340 = ~n1754 & n2339;
  assign n2341 = ~n1744 & n2340;
  assign n2342 = ~n1739 & n2341;
  assign n2343 = ~n1733 & n2342;
  assign n2344 = ~n1728 & n2343;
  assign n2345 = ~n1722 & n2344;
  assign n2346 = ~n1712 & n2345;
  assign n2347 = ~n1701 & n2346;
  assign n2348 = ~n1696 & n2347;
  assign n2349 = ~n1690 & n2348;
  assign n2350 = ~n1685 & n2349;
  assign n2351 = ~n1679 & n2350;
  assign n2352 = ~n1673 & n2351;
  assign n2353 = ~n1666 & n2352;
  assign n2354 = ~n1655 & n2353;
  assign n2355 = ~n1643 & n2354;
  assign n2356 = ~n1637 & n2355;
  assign n2357 = ~n1630 & n2356;
  assign n2358 = ~n1624 & n2357;
  assign n2359 = ~n1617 & n2358;
  assign n2360 = ~n1610 & n2359;
  assign n2361 = ~n1602 & n2360;
  assign n2362 = ~n1590 & n2361;
  assign n2363 = ~n1578 & n2362;
  assign n2364 = ~n1566 & n2363;
  assign n2365 = ~n1553 & n2364;
  assign n2366 = ~n1549 & n2365;
  assign n2367 = ~n1543 & n2366;
  assign n2368 = ~n1538 & n2367;
  assign n2369 = ~n1531 & n2368;
  assign n2370 = ~n1526 & n2369;
  assign n2371 = ~n1519 & n2370;
  assign n2372 = ~n1509 & n2371;
  assign n2373 = ~n1498 & n2372;
  assign n2374 = ~n1493 & n2373;
  assign n2375 = ~n1486 & n2374;
  assign n2376 = ~n1480 & n2375;
  assign n2377 = ~n1472 & n2376;
  assign n2378 = ~n1466 & n2377;
  assign n2379 = ~n1458 & n2378;
  assign n2380 = ~n1445 & n2379;
  assign n2381 = ~n1432 & n2380;
  assign n2382 = ~n1421 & n2381;
  assign n2383 = ~n1409 & n2382;
  assign n2384 = ~n1397 & n2383;
  assign n2385 = ~n1384 & n2384;
  assign n2386 = ~n1378 & n2385;
  assign n2387 = ~n1367 & n2386;
  assign n2388 = ~n1360 & n2387;
  assign n2389 = ~n1348 & n2388;
  assign n2390 = ~n1341 & n2389;
  assign n2391 = ~n1333 & n2390;
  assign n2392 = ~n1320 & n2391;
  assign n2393 = ~n1308 & n2392;
  assign n2394 = ~n1300 & n2393;
  assign n2395 = ~n1291 & n2394;
  assign n2396 = ~n1278 & n2395;
  assign n2397 = ~n1265 & n2396;
  assign n2398 = ~n1252 & n2397;
  assign n2399 = ~n1238 & n2398;
  assign n2400 = ~n1224 & n2399;
  assign n2401 = ~n1210 & n2400;
  assign n2402 = ~n1206 & n2401;
  assign n2403 = ~n1201 & n2402;
  assign n2404 = ~n1197 & n2403;
  assign n2405 = ~n1192 & n2404;
  assign n2406 = ~n1184 & n2405;
  assign n2407 = ~n1175 & n2406;
  assign n2408 = ~n1164 & n2407;
  assign n2409 = ~n1152 & n2408;
  assign n2410 = ~n1147 & n2409;
  assign n2411 = ~n1141 & n2410;
  assign n2412 = ~n1136 & n2411;
  assign n2413 = ~n1130 & n2412;
  assign n2414 = ~n1121 & n2413;
  assign n2415 = ~n1111 & n2414;
  assign n2416 = ~n1100 & n2415;
  assign n2417 = ~n1088 & n2416;
  assign n2418 = ~n1084 & n2417;
  assign n2419 = ~n1079 & n2418;
  assign n2420 = ~n1075 & n2419;
  assign n2421 = ~n1070 & n2420;
  assign n2422 = ~n1065 & n2421;
  assign n2423 = ~n1059 & n2422;
  assign n2424 = ~n1048 & n2423;
  assign n2425 = ~n1036 & n2424;
  assign n2426 = ~n1031 & n2425;
  assign n2427 = ~n1025 & n2426;
  assign n2428 = ~n1020 & n2427;
  assign n2429 = ~n1014 & n2428;
  assign n2430 = ~n1008 & n2429;
  assign n2431 = ~n1001 & n2430;
  assign n2432 = ~n990 & n2431;
  assign n2433 = ~n978 & n2432;
  assign n2434 = ~n972 & n2433;
  assign n2435 = ~n965 & n2434;
  assign n2436 = ~n955 & n2435;
  assign n2437 = ~n944 & n2436;
  assign n2438 = ~n931 & n2437;
  assign n2439 = ~n917 & n2438;
  assign n2440 = ~n910 & n2439;
  assign n2441 = ~n902 & n2440;
  assign n2442 = ~n891 & n2441;
  assign n2443 = ~n879 & n2442;
  assign n2444 = ~n866 & n2443;
  assign n2445 = ~n852 & n2444;
  assign n2446 = ~n848 & n2445;
  assign n2447 = ~n843 & n2446;
  assign n2448 = ~n832 & n2447;
  assign n2449 = ~n827 & n2448;
  assign n2450 = ~n815 & n2449;
  assign n2451 = ~n809 & n2450;
  assign n2452 = ~n797 & n2451;
  assign n2453 = ~n784 & n2452;
  assign n2454 = ~n772 & n2453;
  assign n2455 = ~n759 & n2454;
  assign n2456 = ~n746 & n2455;
  assign n2457 = ~n732 & n2456;
  assign n2458 = ~n731 & n2457;
  assign n2459 = ~n729 & n2458;
  assign n2460 = ~n727 & n2459;
  assign n2461 = ~n725 & n2460;
  assign n2462 = ~n722 & n2461;
  assign n2463 = ~n719 & n2462;
  assign n2464 = ~n716 & n2463;
  assign n2465 = ~n712 & n2464;
  assign n2466 = ~n708 & n2465;
  assign n2467 = ~n704 & n2466;
  assign n2468 = ~n699 & n2467;
  assign n2469 = ~n694 & n2468;
  assign n2470 = ~n688 & n2469;
  assign n2471 = ~n681 & n2470;
  assign n2472 = ~n674 & n2471;
  assign n2473 = ~n666 & n2472;
  assign n2474 = ~n653 & n2473;
  assign n2475 = ~n639 & n2474;
  assign n2476 = ~n632 & n2475;
  assign n2477 = ~n624 & n2476;
  assign n2478 = ~n616 & n2477;
  assign n2479 = ~n607 & n2478;
  assign n2480 = ~n594 & n2479;
  assign n2481 = ~n580 & n2480;
  assign n2482 = ~n577 & n2481;
  assign n2483 = ~n572 & n2482;
  assign n2484 = ~n568 & n2483;
  assign n2485 = ~n562 & n2484;
  assign n2486 = ~n550 & n2485;
  assign n2487 = ~n546 & n2486;
  assign n2488 = ~n532 & n2487;
  assign n2489 = ~n526 & n2488;
  assign n2490 = ~n513 & n2489;
  assign n2491 = ~n508 & n2490;
  assign n2492 = ~n493 & n2491;
  assign n2493 = ~n486 & n2492;
  assign n2494 = ~n473 & n2493;
  assign n2495 = ~n458 & n2494;
  assign n2496 = ~n444 & n2495;
  assign n2497 = ~n426 & n2496;
  assign n2498 = ~n413 & n2497;
  assign n2499 = ~n399 & n2498;
  assign n2500 = ~n384 & n2499;
  assign n2501 = ~n368 & n2500;
  assign n2502 = ~n354 & n2501;
  assign n2503 = ~n339 & n2502;
  assign n0 = n323 | ~n2503;
  assign n2505 = v & n43;
  assign n2506 = ~w & n2505;
  assign n2507 = ~x & n2506;
  assign n2508 = ~y & n2507;
  assign n2509 = ~a0 & n2508;
  assign n2510 = ~b0 & n2509;
  assign n2511 = ~c0 & n2510;
  assign n2512 = d0 & n2511;
  assign n2513 = v & n60;
  assign n2514 = ~w & n2513;
  assign n2515 = ~x & n2514;
  assign n2516 = ~y & n2515;
  assign n2517 = ~a0 & n2516;
  assign n2518 = ~b0 & n2517;
  assign n2519 = ~c0 & n2518;
  assign n2520 = d0 & n2519;
  assign n2521 = v & n77;
  assign n2522 = ~w & n2521;
  assign n2523 = ~x & n2522;
  assign n2524 = ~y & n2523;
  assign n2525 = ~a0 & n2524;
  assign n2526 = ~b0 & n2525;
  assign n2527 = ~c0 & n2526;
  assign n2528 = d0 & n2527;
  assign n2529 = v & n90;
  assign n2530 = ~w & n2529;
  assign n2531 = ~x & n2530;
  assign n2532 = ~y & n2531;
  assign n2533 = ~a0 & n2532;
  assign n2534 = ~b0 & n2533;
  assign n2535 = ~c0 & n2534;
  assign n2536 = d0 & n2535;
  assign n2537 = ~a & ~e;
  assign n2538 = ~f & n2537;
  assign n2539 = ~g & n2538;
  assign n2540 = ~j & n2539;
  assign n2541 = ~n & n2540;
  assign n2542 = ~q & n2541;
  assign n2543 = ~r & n2542;
  assign n2544 = ~u & n2543;
  assign n2545 = ~x & n2544;
  assign n2546 = ~y & n2545;
  assign n2547 = ~a0 & n2546;
  assign n2548 = ~b0 & n2547;
  assign n2549 = ~c0 & n2548;
  assign n2550 = d0 & n2549;
  assign n2551 = ~h0 & n2550;
  assign n2552 = l0 & n2551;
  assign n2553 = d & n2552;
  assign n2554 = ~s & n2553;
  assign n2555 = ~g0 & n2554;
  assign n2556 = ~j0 & n2555;
  assign n2557 = ~l & n2540;
  assign n2558 = ~n & n2557;
  assign n2559 = ~q & n2558;
  assign n2560 = ~r & n2559;
  assign n2561 = ~t & n2560;
  assign n2562 = ~u & n2561;
  assign n2563 = ~x & n2562;
  assign n2564 = ~y & n2563;
  assign n2565 = ~a0 & n2564;
  assign n2566 = ~b0 & n2565;
  assign n2567 = ~c0 & n2566;
  assign n2568 = d0 & n2567;
  assign n2569 = ~h0 & n2568;
  assign n2570 = l0 & n2569;
  assign n2571 = ~g0 & n2570;
  assign n2572 = ~j0 & n2571;
  assign n2573 = ~i & n2539;
  assign n2574 = ~j & n2573;
  assign n2575 = ~n & n2574;
  assign n2576 = ~q & n2575;
  assign n2577 = ~r & n2576;
  assign n2578 = ~u & n2577;
  assign n2579 = ~x & n2578;
  assign n2580 = ~y & n2579;
  assign n2581 = ~a0 & n2580;
  assign n2582 = ~b0 & n2581;
  assign n2583 = ~c0 & n2582;
  assign n2584 = d0 & n2583;
  assign n2585 = ~h0 & n2584;
  assign n2586 = l0 & n2585;
  assign n2587 = d & n2586;
  assign n2588 = ~s & n2587;
  assign n2589 = ~j0 & n2588;
  assign n2590 = ~l & n2574;
  assign n2591 = ~n & n2590;
  assign n2592 = ~q & n2591;
  assign n2593 = ~r & n2592;
  assign n2594 = ~t & n2593;
  assign n2595 = ~u & n2594;
  assign n2596 = ~x & n2595;
  assign n2597 = ~y & n2596;
  assign n2598 = ~a0 & n2597;
  assign n2599 = ~b0 & n2598;
  assign n2600 = ~c0 & n2599;
  assign n2601 = d0 & n2600;
  assign n2602 = ~h0 & n2601;
  assign n2603 = l0 & n2602;
  assign n2604 = ~j0 & n2603;
  assign n2605 = ~h & n2539;
  assign n2606 = ~j & n2605;
  assign n2607 = ~n & n2606;
  assign n2608 = ~q & n2607;
  assign n2609 = ~r & n2608;
  assign n2610 = ~u & n2609;
  assign n2611 = ~x & n2610;
  assign n2612 = ~y & n2611;
  assign n2613 = ~a0 & n2612;
  assign n2614 = ~b0 & n2613;
  assign n2615 = ~c0 & n2614;
  assign n2616 = d0 & n2615;
  assign n2617 = ~h0 & n2616;
  assign n2618 = l0 & n2617;
  assign n2619 = d & n2618;
  assign n2620 = ~s & n2619;
  assign n2621 = ~g0 & n2620;
  assign n2622 = ~l & n2606;
  assign n2623 = ~n & n2622;
  assign n2624 = ~q & n2623;
  assign n2625 = ~r & n2624;
  assign n2626 = ~t & n2625;
  assign n2627 = ~u & n2626;
  assign n2628 = ~x & n2627;
  assign n2629 = ~y & n2628;
  assign n2630 = ~a0 & n2629;
  assign n2631 = ~b0 & n2630;
  assign n2632 = ~c0 & n2631;
  assign n2633 = d0 & n2632;
  assign n2634 = ~h0 & n2633;
  assign n2635 = l0 & n2634;
  assign n2636 = ~g0 & n2635;
  assign n2637 = ~i & n2605;
  assign n2638 = ~j & n2637;
  assign n2639 = ~n & n2638;
  assign n2640 = ~q & n2639;
  assign n2641 = ~r & n2640;
  assign n2642 = ~u & n2641;
  assign n2643 = ~x & n2642;
  assign n2644 = ~y & n2643;
  assign n2645 = ~a0 & n2644;
  assign n2646 = ~b0 & n2645;
  assign n2647 = ~c0 & n2646;
  assign n2648 = d0 & n2647;
  assign n2649 = ~h0 & n2648;
  assign n2650 = l0 & n2649;
  assign n2651 = d & n2650;
  assign n2652 = ~s & n2651;
  assign n2653 = ~l & n2638;
  assign n2654 = ~n & n2653;
  assign n2655 = ~q & n2654;
  assign n2656 = ~r & n2655;
  assign n2657 = ~t & n2656;
  assign n2658 = ~u & n2657;
  assign n2659 = ~x & n2658;
  assign n2660 = ~y & n2659;
  assign n2661 = ~a0 & n2660;
  assign n2662 = ~b0 & n2661;
  assign n2663 = ~c0 & n2662;
  assign n2664 = d0 & n2663;
  assign n2665 = ~h0 & n2664;
  assign n2666 = l0 & n2665;
  assign n2667 = ~g0 & n2552;
  assign n2668 = ~j0 & n2667;
  assign n2669 = ~k & n2668;
  assign n2670 = ~j0 & n2586;
  assign n2671 = ~k & n2670;
  assign n2672 = ~g0 & n2618;
  assign n2673 = ~k & n2672;
  assign n2674 = ~k & n2650;
  assign n2675 = ~d0 & n331;
  assign n2676 = ~h0 & n2675;
  assign n2677 = l0 & n2676;
  assign n2678 = d & n2677;
  assign n2679 = ~s & n2678;
  assign n2680 = ~g0 & n2679;
  assign n2681 = j0 & n2680;
  assign n2682 = ~c & n2681;
  assign n2683 = ~i0 & n2682;
  assign n2684 = ~d0 & n362;
  assign n2685 = ~h0 & n2684;
  assign n2686 = l0 & n2685;
  assign n2687 = ~g0 & n2686;
  assign n2688 = j0 & n2687;
  assign n2689 = ~c & n2688;
  assign n2690 = ~i0 & n2689;
  assign n2691 = ~d0 & n392;
  assign n2692 = ~h0 & n2691;
  assign n2693 = l0 & n2692;
  assign n2694 = d & n2693;
  assign n2695 = ~s & n2694;
  assign n2696 = j0 & n2695;
  assign n2697 = ~c & n2696;
  assign n2698 = ~i0 & n2697;
  assign n2699 = ~d0 & n421;
  assign n2700 = ~h0 & n2699;
  assign n2701 = l0 & n2700;
  assign n2702 = j0 & n2701;
  assign n2703 = ~c & n2702;
  assign n2704 = ~i0 & n2703;
  assign n2705 = ~y & n312;
  assign n2706 = ~b0 & n2705;
  assign n2707 = ~c0 & n2706;
  assign n2708 = ~d0 & n2707;
  assign n2709 = ~h0 & n2708;
  assign n2710 = l0 & n2709;
  assign n2711 = d & n2710;
  assign n2712 = ~s & n2711;
  assign n2713 = ~g0 & n2712;
  assign n2714 = ~j0 & n2713;
  assign n2715 = ~c & n2714;
  assign n2716 = i0 & n2715;
  assign n2717 = ~y & n345;
  assign n2718 = ~b0 & n2717;
  assign n2719 = ~c0 & n2718;
  assign n2720 = ~d0 & n2719;
  assign n2721 = ~h0 & n2720;
  assign n2722 = l0 & n2721;
  assign n2723 = ~g0 & n2722;
  assign n2724 = ~j0 & n2723;
  assign n2725 = ~c & n2724;
  assign n2726 = i0 & n2725;
  assign n2727 = ~y & n374;
  assign n2728 = ~b0 & n2727;
  assign n2729 = ~c0 & n2728;
  assign n2730 = ~d0 & n2729;
  assign n2731 = ~h0 & n2730;
  assign n2732 = l0 & n2731;
  assign n2733 = d & n2732;
  assign n2734 = ~s & n2733;
  assign n2735 = ~j0 & n2734;
  assign n2736 = ~c & n2735;
  assign n2737 = i0 & n2736;
  assign n2738 = ~y & n405;
  assign n2739 = ~b0 & n2738;
  assign n2740 = ~c0 & n2739;
  assign n2741 = ~d0 & n2740;
  assign n2742 = ~h0 & n2741;
  assign n2743 = l0 & n2742;
  assign n2744 = ~j0 & n2743;
  assign n2745 = ~c & n2744;
  assign n2746 = i0 & n2745;
  assign n2747 = ~y & n329;
  assign n2748 = ~b0 & n2747;
  assign n2749 = ~c0 & n2748;
  assign n2750 = ~d0 & n2749;
  assign n2751 = ~h0 & n2750;
  assign n2752 = l0 & n2751;
  assign n2753 = d & n2752;
  assign n2754 = ~s & n2753;
  assign n2755 = ~g0 & n2754;
  assign n2756 = ~c & n2755;
  assign n2757 = i0 & n2756;
  assign n2758 = ~y & n360;
  assign n2759 = ~b0 & n2758;
  assign n2760 = ~c0 & n2759;
  assign n2761 = ~d0 & n2760;
  assign n2762 = ~h0 & n2761;
  assign n2763 = l0 & n2762;
  assign n2764 = ~g0 & n2763;
  assign n2765 = ~c & n2764;
  assign n2766 = i0 & n2765;
  assign n2767 = ~y & n390;
  assign n2768 = ~b0 & n2767;
  assign n2769 = ~c0 & n2768;
  assign n2770 = ~d0 & n2769;
  assign n2771 = ~h0 & n2770;
  assign n2772 = l0 & n2771;
  assign n2773 = d & n2772;
  assign n2774 = ~s & n2773;
  assign n2775 = ~c & n2774;
  assign n2776 = i0 & n2775;
  assign n2777 = ~y & n419;
  assign n2778 = ~b0 & n2777;
  assign n2779 = ~c0 & n2778;
  assign n2780 = ~d0 & n2779;
  assign n2781 = ~h0 & n2780;
  assign n2782 = l0 & n2781;
  assign n2783 = ~c & n2782;
  assign n2784 = i0 & n2783;
  assign n2785 = ~a0 & n2705;
  assign n2786 = ~b0 & n2785;
  assign n2787 = ~c0 & n2786;
  assign n2788 = ~d0 & n2787;
  assign n2789 = ~h0 & n2788;
  assign n2790 = l0 & n2789;
  assign n2791 = d & n2790;
  assign n2792 = ~s & n2791;
  assign n2793 = ~g0 & n2792;
  assign n2794 = ~j0 & n2793;
  assign n2795 = ~c & n2794;
  assign n2796 = ~a0 & n2717;
  assign n2797 = ~b0 & n2796;
  assign n2798 = ~c0 & n2797;
  assign n2799 = ~d0 & n2798;
  assign n2800 = ~h0 & n2799;
  assign n2801 = l0 & n2800;
  assign n2802 = ~g0 & n2801;
  assign n2803 = ~j0 & n2802;
  assign n2804 = ~c & n2803;
  assign n2805 = ~a0 & n2727;
  assign n2806 = ~b0 & n2805;
  assign n2807 = ~c0 & n2806;
  assign n2808 = ~d0 & n2807;
  assign n2809 = ~h0 & n2808;
  assign n2810 = l0 & n2809;
  assign n2811 = d & n2810;
  assign n2812 = ~s & n2811;
  assign n2813 = ~j0 & n2812;
  assign n2814 = ~c & n2813;
  assign n2815 = ~a0 & n2738;
  assign n2816 = ~b0 & n2815;
  assign n2817 = ~c0 & n2816;
  assign n2818 = ~d0 & n2817;
  assign n2819 = ~h0 & n2818;
  assign n2820 = l0 & n2819;
  assign n2821 = ~j0 & n2820;
  assign n2822 = ~c & n2821;
  assign n2823 = ~q & n2540;
  assign n2824 = ~r & n2823;
  assign n2825 = ~u & n2824;
  assign n2826 = ~x & n2825;
  assign n2827 = ~y & n2826;
  assign n2828 = ~a0 & n2827;
  assign n2829 = ~b0 & n2828;
  assign n2830 = ~c0 & n2829;
  assign n2831 = d0 & n2830;
  assign n2832 = l0 & n2831;
  assign n2833 = d & n2832;
  assign n2834 = ~s & n2833;
  assign n2835 = ~g0 & n2834;
  assign n2836 = ~j0 & n2835;
  assign n2837 = ~o & n2836;
  assign n2838 = ~q & n2557;
  assign n2839 = ~r & n2838;
  assign n2840 = ~t & n2839;
  assign n2841 = ~u & n2840;
  assign n2842 = ~x & n2841;
  assign n2843 = ~y & n2842;
  assign n2844 = ~a0 & n2843;
  assign n2845 = ~b0 & n2844;
  assign n2846 = ~c0 & n2845;
  assign n2847 = d0 & n2846;
  assign n2848 = l0 & n2847;
  assign n2849 = ~g0 & n2848;
  assign n2850 = ~j0 & n2849;
  assign n2851 = ~o & n2850;
  assign n2852 = ~q & n2574;
  assign n2853 = ~r & n2852;
  assign n2854 = ~u & n2853;
  assign n2855 = ~x & n2854;
  assign n2856 = ~y & n2855;
  assign n2857 = ~a0 & n2856;
  assign n2858 = ~b0 & n2857;
  assign n2859 = ~c0 & n2858;
  assign n2860 = d0 & n2859;
  assign n2861 = l0 & n2860;
  assign n2862 = d & n2861;
  assign n2863 = ~s & n2862;
  assign n2864 = ~j0 & n2863;
  assign n2865 = ~o & n2864;
  assign n2866 = ~q & n2590;
  assign n2867 = ~r & n2866;
  assign n2868 = ~t & n2867;
  assign n2869 = ~u & n2868;
  assign n2870 = ~x & n2869;
  assign n2871 = ~y & n2870;
  assign n2872 = ~a0 & n2871;
  assign n2873 = ~b0 & n2872;
  assign n2874 = ~c0 & n2873;
  assign n2875 = d0 & n2874;
  assign n2876 = l0 & n2875;
  assign n2877 = ~j0 & n2876;
  assign n2878 = ~o & n2877;
  assign n2879 = ~q & n2606;
  assign n2880 = ~r & n2879;
  assign n2881 = ~u & n2880;
  assign n2882 = ~x & n2881;
  assign n2883 = ~y & n2882;
  assign n2884 = ~a0 & n2883;
  assign n2885 = ~b0 & n2884;
  assign n2886 = ~c0 & n2885;
  assign n2887 = d0 & n2886;
  assign n2888 = l0 & n2887;
  assign n2889 = d & n2888;
  assign n2890 = ~s & n2889;
  assign n2891 = ~g0 & n2890;
  assign n2892 = ~o & n2891;
  assign n2893 = ~q & n2622;
  assign n2894 = ~r & n2893;
  assign n2895 = ~t & n2894;
  assign n2896 = ~u & n2895;
  assign n2897 = ~x & n2896;
  assign n2898 = ~y & n2897;
  assign n2899 = ~a0 & n2898;
  assign n2900 = ~b0 & n2899;
  assign n2901 = ~c0 & n2900;
  assign n2902 = d0 & n2901;
  assign n2903 = l0 & n2902;
  assign n2904 = ~g0 & n2903;
  assign n2905 = ~o & n2904;
  assign n2906 = ~q & n2638;
  assign n2907 = ~r & n2906;
  assign n2908 = ~u & n2907;
  assign n2909 = ~x & n2908;
  assign n2910 = ~y & n2909;
  assign n2911 = ~a0 & n2910;
  assign n2912 = ~b0 & n2911;
  assign n2913 = ~c0 & n2912;
  assign n2914 = d0 & n2913;
  assign n2915 = l0 & n2914;
  assign n2916 = d & n2915;
  assign n2917 = ~s & n2916;
  assign n2918 = ~o & n2917;
  assign n2919 = ~q & n2653;
  assign n2920 = ~r & n2919;
  assign n2921 = ~t & n2920;
  assign n2922 = ~u & n2921;
  assign n2923 = ~x & n2922;
  assign n2924 = ~y & n2923;
  assign n2925 = ~a0 & n2924;
  assign n2926 = ~b0 & n2925;
  assign n2927 = ~c0 & n2926;
  assign n2928 = d0 & n2927;
  assign n2929 = l0 & n2928;
  assign n2930 = ~o & n2929;
  assign n2931 = ~n & n2539;
  assign n2932 = ~q & n2931;
  assign n2933 = ~r & n2932;
  assign n2934 = ~u & n2933;
  assign n2935 = ~x & n2934;
  assign n2936 = ~y & n2935;
  assign n2937 = ~a0 & n2936;
  assign n2938 = ~b0 & n2937;
  assign n2939 = ~c0 & n2938;
  assign n2940 = d0 & n2939;
  assign n2941 = ~h0 & n2940;
  assign n2942 = l0 & n2941;
  assign n2943 = ~g0 & n2942;
  assign n2944 = ~j0 & n2943;
  assign n2945 = ~b & n2944;
  assign n2946 = ~n & n2573;
  assign n2947 = ~q & n2946;
  assign n2948 = ~r & n2947;
  assign n2949 = ~u & n2948;
  assign n2950 = ~x & n2949;
  assign n2951 = ~y & n2950;
  assign n2952 = ~a0 & n2951;
  assign n2953 = ~b0 & n2952;
  assign n2954 = ~c0 & n2953;
  assign n2955 = d0 & n2954;
  assign n2956 = ~h0 & n2955;
  assign n2957 = l0 & n2956;
  assign n2958 = ~j0 & n2957;
  assign n2959 = ~b & n2958;
  assign n2960 = ~n & n2605;
  assign n2961 = ~q & n2960;
  assign n2962 = ~r & n2961;
  assign n2963 = ~u & n2962;
  assign n2964 = ~x & n2963;
  assign n2965 = ~y & n2964;
  assign n2966 = ~a0 & n2965;
  assign n2967 = ~b0 & n2966;
  assign n2968 = ~c0 & n2967;
  assign n2969 = d0 & n2968;
  assign n2970 = ~h0 & n2969;
  assign n2971 = l0 & n2970;
  assign n2972 = ~g0 & n2971;
  assign n2973 = ~b & n2972;
  assign n2974 = ~n & n2637;
  assign n2975 = ~q & n2974;
  assign n2976 = ~r & n2975;
  assign n2977 = ~u & n2976;
  assign n2978 = ~x & n2977;
  assign n2979 = ~y & n2978;
  assign n2980 = ~a0 & n2979;
  assign n2981 = ~b0 & n2980;
  assign n2982 = ~c0 & n2981;
  assign n2983 = d0 & n2982;
  assign n2984 = ~h0 & n2983;
  assign n2985 = l0 & n2984;
  assign n2986 = ~b & n2985;
  assign n2987 = ~g0 & n2677;
  assign n2988 = j0 & n2987;
  assign n2989 = ~c & n2988;
  assign n2990 = ~i0 & n2989;
  assign n2991 = ~k & n2990;
  assign n2992 = j0 & n2693;
  assign n2993 = ~c & n2992;
  assign n2994 = ~i0 & n2993;
  assign n2995 = ~k & n2994;
  assign n2996 = ~g0 & n2710;
  assign n2997 = ~j0 & n2996;
  assign n2998 = ~c & n2997;
  assign n2999 = i0 & n2998;
  assign n3000 = ~k & n2999;
  assign n3001 = ~j0 & n2732;
  assign n3002 = ~c & n3001;
  assign n3003 = i0 & n3002;
  assign n3004 = ~k & n3003;
  assign n3005 = ~g0 & n2752;
  assign n3006 = ~c & n3005;
  assign n3007 = i0 & n3006;
  assign n3008 = ~k & n3007;
  assign n3009 = ~c & n2772;
  assign n3010 = i0 & n3009;
  assign n3011 = ~k & n3010;
  assign n3012 = ~g0 & n2790;
  assign n3013 = ~j0 & n3012;
  assign n3014 = ~c & n3013;
  assign n3015 = ~k & n3014;
  assign n3016 = ~j0 & n2810;
  assign n3017 = ~c & n3016;
  assign n3018 = ~k & n3017;
  assign n3019 = ~g0 & n2832;
  assign n3020 = ~j0 & n3019;
  assign n3021 = ~o & n3020;
  assign n3022 = ~k & n3021;
  assign n3023 = ~j0 & n2861;
  assign n3024 = ~o & n3023;
  assign n3025 = ~k & n3024;
  assign n3026 = ~g0 & n2888;
  assign n3027 = ~o & n3026;
  assign n3028 = ~k & n3027;
  assign n3029 = ~o & n2915;
  assign n3030 = ~k & n3029;
  assign n3031 = ~q & n325;
  assign n3032 = ~r & n3031;
  assign n3033 = ~x & n3032;
  assign n3034 = ~b0 & n3033;
  assign n3035 = ~c0 & n3034;
  assign n3036 = ~d0 & n3035;
  assign n3037 = l0 & n3036;
  assign n3038 = d & n3037;
  assign n3039 = ~s & n3038;
  assign n3040 = ~g0 & n3039;
  assign n3041 = j0 & n3040;
  assign n3042 = ~o & n3041;
  assign n3043 = ~c & n3042;
  assign n3044 = ~i0 & n3043;
  assign n3045 = ~q & n355;
  assign n3046 = ~r & n3045;
  assign n3047 = ~t & n3046;
  assign n3048 = ~x & n3047;
  assign n3049 = ~b0 & n3048;
  assign n3050 = ~c0 & n3049;
  assign n3051 = ~d0 & n3050;
  assign n3052 = l0 & n3051;
  assign n3053 = ~g0 & n3052;
  assign n3054 = j0 & n3053;
  assign n3055 = ~o & n3054;
  assign n3056 = ~c & n3055;
  assign n3057 = ~i0 & n3056;
  assign n3058 = ~q & n386;
  assign n3059 = ~r & n3058;
  assign n3060 = ~x & n3059;
  assign n3061 = ~b0 & n3060;
  assign n3062 = ~c0 & n3061;
  assign n3063 = ~d0 & n3062;
  assign n3064 = l0 & n3063;
  assign n3065 = d & n3064;
  assign n3066 = ~s & n3065;
  assign n3067 = j0 & n3066;
  assign n3068 = ~o & n3067;
  assign n3069 = ~c & n3068;
  assign n3070 = ~i0 & n3069;
  assign n3071 = ~q & n414;
  assign n3072 = ~r & n3071;
  assign n3073 = ~t & n3072;
  assign n3074 = ~x & n3073;
  assign n3075 = ~b0 & n3074;
  assign n3076 = ~c0 & n3075;
  assign n3077 = ~d0 & n3076;
  assign n3078 = l0 & n3077;
  assign n3079 = j0 & n3078;
  assign n3080 = ~o & n3079;
  assign n3081 = ~c & n3080;
  assign n3082 = ~i0 & n3081;
  assign n3083 = ~q & n308;
  assign n3084 = ~r & n3083;
  assign n3085 = ~x & n3084;
  assign n3086 = ~y & n3085;
  assign n3087 = ~b0 & n3086;
  assign n3088 = ~c0 & n3087;
  assign n3089 = ~d0 & n3088;
  assign n3090 = l0 & n3089;
  assign n3091 = d & n3090;
  assign n3092 = ~s & n3091;
  assign n3093 = ~g0 & n3092;
  assign n3094 = ~j0 & n3093;
  assign n3095 = ~o & n3094;
  assign n3096 = ~c & n3095;
  assign n3097 = i0 & n3096;
  assign n3098 = ~q & n340;
  assign n3099 = ~r & n3098;
  assign n3100 = ~t & n3099;
  assign n3101 = ~x & n3100;
  assign n3102 = ~y & n3101;
  assign n3103 = ~b0 & n3102;
  assign n3104 = ~c0 & n3103;
  assign n3105 = ~d0 & n3104;
  assign n3106 = l0 & n3105;
  assign n3107 = ~g0 & n3106;
  assign n3108 = ~j0 & n3107;
  assign n3109 = ~o & n3108;
  assign n3110 = ~c & n3109;
  assign n3111 = i0 & n3110;
  assign n3112 = ~q & n370;
  assign n3113 = ~r & n3112;
  assign n3114 = ~x & n3113;
  assign n3115 = ~y & n3114;
  assign n3116 = ~b0 & n3115;
  assign n3117 = ~c0 & n3116;
  assign n3118 = ~d0 & n3117;
  assign n3119 = l0 & n3118;
  assign n3120 = d & n3119;
  assign n3121 = ~s & n3120;
  assign n3122 = ~j0 & n3121;
  assign n3123 = ~o & n3122;
  assign n3124 = ~c & n3123;
  assign n3125 = i0 & n3124;
  assign n3126 = ~q & n400;
  assign n3127 = ~r & n3126;
  assign n3128 = ~t & n3127;
  assign n3129 = ~x & n3128;
  assign n3130 = ~y & n3129;
  assign n3131 = ~b0 & n3130;
  assign n3132 = ~c0 & n3131;
  assign n3133 = ~d0 & n3132;
  assign n3134 = l0 & n3133;
  assign n3135 = ~j0 & n3134;
  assign n3136 = ~o & n3135;
  assign n3137 = ~c & n3136;
  assign n3138 = i0 & n3137;
  assign n3139 = ~y & n3033;
  assign n3140 = ~b0 & n3139;
  assign n3141 = ~c0 & n3140;
  assign n3142 = ~d0 & n3141;
  assign n3143 = l0 & n3142;
  assign n3144 = d & n3143;
  assign n3145 = ~s & n3144;
  assign n3146 = ~g0 & n3145;
  assign n3147 = ~o & n3146;
  assign n3148 = ~c & n3147;
  assign n3149 = i0 & n3148;
  assign n3150 = ~y & n3048;
  assign n3151 = ~b0 & n3150;
  assign n3152 = ~c0 & n3151;
  assign n3153 = ~d0 & n3152;
  assign n3154 = l0 & n3153;
  assign n3155 = ~g0 & n3154;
  assign n3156 = ~o & n3155;
  assign n3157 = ~c & n3156;
  assign n3158 = i0 & n3157;
  assign n3159 = ~y & n3060;
  assign n3160 = ~b0 & n3159;
  assign n3161 = ~c0 & n3160;
  assign n3162 = ~d0 & n3161;
  assign n3163 = l0 & n3162;
  assign n3164 = d & n3163;
  assign n3165 = ~s & n3164;
  assign n3166 = ~o & n3165;
  assign n3167 = ~c & n3166;
  assign n3168 = i0 & n3167;
  assign n3169 = ~y & n3074;
  assign n3170 = ~b0 & n3169;
  assign n3171 = ~c0 & n3170;
  assign n3172 = ~d0 & n3171;
  assign n3173 = l0 & n3172;
  assign n3174 = ~o & n3173;
  assign n3175 = ~c & n3174;
  assign n3176 = i0 & n3175;
  assign n3177 = ~a0 & n3086;
  assign n3178 = ~b0 & n3177;
  assign n3179 = ~c0 & n3178;
  assign n3180 = ~d0 & n3179;
  assign n3181 = l0 & n3180;
  assign n3182 = d & n3181;
  assign n3183 = ~s & n3182;
  assign n3184 = ~g0 & n3183;
  assign n3185 = ~j0 & n3184;
  assign n3186 = ~o & n3185;
  assign n3187 = ~c & n3186;
  assign n3188 = ~a0 & n3102;
  assign n3189 = ~b0 & n3188;
  assign n3190 = ~c0 & n3189;
  assign n3191 = ~d0 & n3190;
  assign n3192 = l0 & n3191;
  assign n3193 = ~g0 & n3192;
  assign n3194 = ~j0 & n3193;
  assign n3195 = ~o & n3194;
  assign n3196 = ~c & n3195;
  assign n3197 = ~a0 & n3115;
  assign n3198 = ~b0 & n3197;
  assign n3199 = ~c0 & n3198;
  assign n3200 = ~d0 & n3199;
  assign n3201 = l0 & n3200;
  assign n3202 = d & n3201;
  assign n3203 = ~s & n3202;
  assign n3204 = ~j0 & n3203;
  assign n3205 = ~o & n3204;
  assign n3206 = ~c & n3205;
  assign n3207 = ~a0 & n3130;
  assign n3208 = ~b0 & n3207;
  assign n3209 = ~c0 & n3208;
  assign n3210 = ~d0 & n3209;
  assign n3211 = l0 & n3210;
  assign n3212 = ~j0 & n3211;
  assign n3213 = ~o & n3212;
  assign n3214 = ~c & n3213;
  assign n3215 = n & n2540;
  assign n3216 = ~q & n3215;
  assign n3217 = ~r & n3216;
  assign n3218 = ~u & n3217;
  assign n3219 = ~x & n3218;
  assign n3220 = ~y & n3219;
  assign n3221 = ~a0 & n3220;
  assign n3222 = ~b0 & n3221;
  assign n3223 = ~c0 & n3222;
  assign n3224 = d0 & n3223;
  assign n3225 = l0 & n3224;
  assign n3226 = ~g0 & n3225;
  assign n3227 = ~j0 & n3226;
  assign n3228 = ~o & n3227;
  assign n3229 = n & n2574;
  assign n3230 = ~q & n3229;
  assign n3231 = ~r & n3230;
  assign n3232 = ~u & n3231;
  assign n3233 = ~x & n3232;
  assign n3234 = ~y & n3233;
  assign n3235 = ~a0 & n3234;
  assign n3236 = ~b0 & n3235;
  assign n3237 = ~c0 & n3236;
  assign n3238 = d0 & n3237;
  assign n3239 = l0 & n3238;
  assign n3240 = ~j0 & n3239;
  assign n3241 = ~o & n3240;
  assign n3242 = n & n2606;
  assign n3243 = ~q & n3242;
  assign n3244 = ~r & n3243;
  assign n3245 = ~u & n3244;
  assign n3246 = ~x & n3245;
  assign n3247 = ~y & n3246;
  assign n3248 = ~a0 & n3247;
  assign n3249 = ~b0 & n3248;
  assign n3250 = ~c0 & n3249;
  assign n3251 = d0 & n3250;
  assign n3252 = l0 & n3251;
  assign n3253 = ~g0 & n3252;
  assign n3254 = ~o & n3253;
  assign n3255 = n & n2638;
  assign n3256 = ~q & n3255;
  assign n3257 = ~r & n3256;
  assign n3258 = ~u & n3257;
  assign n3259 = ~x & n3258;
  assign n3260 = ~y & n3259;
  assign n3261 = ~a0 & n3260;
  assign n3262 = ~b0 & n3261;
  assign n3263 = ~c0 & n3262;
  assign n3264 = d0 & n3263;
  assign n3265 = l0 & n3264;
  assign n3266 = ~o & n3265;
  assign n3267 = ~u & n2932;
  assign n3268 = ~x & n3267;
  assign n3269 = ~y & n3268;
  assign n3270 = ~a0 & n3269;
  assign n3271 = ~b0 & n3270;
  assign n3272 = ~c0 & n3271;
  assign n3273 = d0 & n3272;
  assign n3274 = ~h0 & n3273;
  assign n3275 = l0 & n3274;
  assign n3276 = ~g0 & n3275;
  assign n3277 = ~j0 & n3276;
  assign n3278 = ~m & n3277;
  assign n3279 = ~u & n2947;
  assign n3280 = ~x & n3279;
  assign n3281 = ~y & n3280;
  assign n3282 = ~a0 & n3281;
  assign n3283 = ~b0 & n3282;
  assign n3284 = ~c0 & n3283;
  assign n3285 = d0 & n3284;
  assign n3286 = ~h0 & n3285;
  assign n3287 = l0 & n3286;
  assign n3288 = ~j0 & n3287;
  assign n3289 = ~m & n3288;
  assign n3290 = ~u & n2961;
  assign n3291 = ~x & n3290;
  assign n3292 = ~y & n3291;
  assign n3293 = ~a0 & n3292;
  assign n3294 = ~b0 & n3293;
  assign n3295 = ~c0 & n3294;
  assign n3296 = d0 & n3295;
  assign n3297 = ~h0 & n3296;
  assign n3298 = l0 & n3297;
  assign n3299 = ~g0 & n3298;
  assign n3300 = ~m & n3299;
  assign n3301 = ~u & n2975;
  assign n3302 = ~x & n3301;
  assign n3303 = ~y & n3302;
  assign n3304 = ~a0 & n3303;
  assign n3305 = ~b0 & n3304;
  assign n3306 = ~c0 & n3305;
  assign n3307 = d0 & n3306;
  assign n3308 = ~h0 & n3307;
  assign n3309 = l0 & n3308;
  assign n3310 = ~m & n3309;
  assign n3311 = ~r & n1154;
  assign n3312 = ~x & n3311;
  assign n3313 = ~b0 & n3312;
  assign n3314 = ~c0 & n3313;
  assign n3315 = ~d0 & n3314;
  assign n3316 = ~h0 & n3315;
  assign n3317 = l0 & n3316;
  assign n3318 = ~g0 & n3317;
  assign n3319 = j0 & n3318;
  assign n3320 = ~c & n3319;
  assign n3321 = ~i0 & n3320;
  assign n3322 = ~b & n3321;
  assign n3323 = ~r & n1166;
  assign n3324 = ~x & n3323;
  assign n3325 = ~b0 & n3324;
  assign n3326 = ~c0 & n3325;
  assign n3327 = ~d0 & n3326;
  assign n3328 = ~h0 & n3327;
  assign n3329 = l0 & n3328;
  assign n3330 = j0 & n3329;
  assign n3331 = ~c & n3330;
  assign n3332 = ~i0 & n3331;
  assign n3333 = ~b & n3332;
  assign n3334 = ~r & n919;
  assign n3335 = ~x & n3334;
  assign n3336 = ~y & n3335;
  assign n3337 = ~b0 & n3336;
  assign n3338 = ~c0 & n3337;
  assign n3339 = ~d0 & n3338;
  assign n3340 = ~h0 & n3339;
  assign n3341 = l0 & n3340;
  assign n3342 = ~g0 & n3341;
  assign n3343 = ~j0 & n3342;
  assign n3344 = ~c & n3343;
  assign n3345 = i0 & n3344;
  assign n3346 = ~b & n3345;
  assign n3347 = ~r & n933;
  assign n3348 = ~x & n3347;
  assign n3349 = ~y & n3348;
  assign n3350 = ~b0 & n3349;
  assign n3351 = ~c0 & n3350;
  assign n3352 = ~d0 & n3351;
  assign n3353 = ~h0 & n3352;
  assign n3354 = l0 & n3353;
  assign n3355 = ~j0 & n3354;
  assign n3356 = ~c & n3355;
  assign n3357 = i0 & n3356;
  assign n3358 = ~b & n3357;
  assign n3359 = ~y & n3312;
  assign n3360 = ~b0 & n3359;
  assign n3361 = ~c0 & n3360;
  assign n3362 = ~d0 & n3361;
  assign n3363 = ~h0 & n3362;
  assign n3364 = l0 & n3363;
  assign n3365 = ~g0 & n3364;
  assign n3366 = ~c & n3365;
  assign n3367 = i0 & n3366;
  assign n3368 = ~b & n3367;
  assign n3369 = ~y & n3324;
  assign n3370 = ~b0 & n3369;
  assign n3371 = ~c0 & n3370;
  assign n3372 = ~d0 & n3371;
  assign n3373 = ~h0 & n3372;
  assign n3374 = l0 & n3373;
  assign n3375 = ~c & n3374;
  assign n3376 = i0 & n3375;
  assign n3377 = ~b & n3376;
  assign n3378 = ~a0 & n3336;
  assign n3379 = ~b0 & n3378;
  assign n3380 = ~c0 & n3379;
  assign n3381 = ~d0 & n3380;
  assign n3382 = ~h0 & n3381;
  assign n3383 = l0 & n3382;
  assign n3384 = ~g0 & n3383;
  assign n3385 = ~j0 & n3384;
  assign n3386 = ~c & n3385;
  assign n3387 = ~b & n3386;
  assign n3388 = ~a0 & n3349;
  assign n3389 = ~b0 & n3388;
  assign n3390 = ~c0 & n3389;
  assign n3391 = ~d0 & n3390;
  assign n3392 = ~h0 & n3391;
  assign n3393 = l0 & n3392;
  assign n3394 = ~j0 & n3393;
  assign n3395 = ~c & n3394;
  assign n3396 = ~b & n3395;
  assign n3397 = ~q & n2539;
  assign n3398 = ~r & n3397;
  assign n3399 = ~u & n3398;
  assign n3400 = ~x & n3399;
  assign n3401 = ~y & n3400;
  assign n3402 = ~a0 & n3401;
  assign n3403 = ~b0 & n3402;
  assign n3404 = ~c0 & n3403;
  assign n3405 = d0 & n3404;
  assign n3406 = l0 & n3405;
  assign n3407 = ~g0 & n3406;
  assign n3408 = ~j0 & n3407;
  assign n3409 = ~o & n3408;
  assign n3410 = ~b & n3409;
  assign n3411 = ~q & n2573;
  assign n3412 = ~r & n3411;
  assign n3413 = ~u & n3412;
  assign n3414 = ~x & n3413;
  assign n3415 = ~y & n3414;
  assign n3416 = ~a0 & n3415;
  assign n3417 = ~b0 & n3416;
  assign n3418 = ~c0 & n3417;
  assign n3419 = d0 & n3418;
  assign n3420 = l0 & n3419;
  assign n3421 = ~j0 & n3420;
  assign n3422 = ~o & n3421;
  assign n3423 = ~b & n3422;
  assign n3424 = ~q & n2605;
  assign n3425 = ~r & n3424;
  assign n3426 = ~u & n3425;
  assign n3427 = ~x & n3426;
  assign n3428 = ~y & n3427;
  assign n3429 = ~a0 & n3428;
  assign n3430 = ~b0 & n3429;
  assign n3431 = ~c0 & n3430;
  assign n3432 = d0 & n3431;
  assign n3433 = l0 & n3432;
  assign n3434 = ~g0 & n3433;
  assign n3435 = ~o & n3434;
  assign n3436 = ~b & n3435;
  assign n3437 = ~q & n2637;
  assign n3438 = ~r & n3437;
  assign n3439 = ~u & n3438;
  assign n3440 = ~x & n3439;
  assign n3441 = ~y & n3440;
  assign n3442 = ~a0 & n3441;
  assign n3443 = ~b0 & n3442;
  assign n3444 = ~c0 & n3443;
  assign n3445 = d0 & n3444;
  assign n3446 = l0 & n3445;
  assign n3447 = ~o & n3446;
  assign n3448 = ~b & n3447;
  assign n3449 = ~g0 & n3037;
  assign n3450 = j0 & n3449;
  assign n3451 = ~o & n3450;
  assign n3452 = ~c & n3451;
  assign n3453 = ~i0 & n3452;
  assign n3454 = ~k & n3453;
  assign n3455 = j0 & n3064;
  assign n3456 = ~o & n3455;
  assign n3457 = ~c & n3456;
  assign n3458 = ~i0 & n3457;
  assign n3459 = ~k & n3458;
  assign n3460 = ~g0 & n3090;
  assign n3461 = ~j0 & n3460;
  assign n3462 = ~o & n3461;
  assign n3463 = ~c & n3462;
  assign n3464 = i0 & n3463;
  assign n3465 = ~k & n3464;
  assign n3466 = ~j0 & n3119;
  assign n3467 = ~o & n3466;
  assign n3468 = ~c & n3467;
  assign n3469 = i0 & n3468;
  assign n3470 = ~k & n3469;
  assign n3471 = ~g0 & n3143;
  assign n3472 = ~o & n3471;
  assign n3473 = ~c & n3472;
  assign n3474 = i0 & n3473;
  assign n3475 = ~k & n3474;
  assign n3476 = ~o & n3163;
  assign n3477 = ~c & n3476;
  assign n3478 = i0 & n3477;
  assign n3479 = ~k & n3478;
  assign n3480 = ~g0 & n3181;
  assign n3481 = ~j0 & n3480;
  assign n3482 = ~o & n3481;
  assign n3483 = ~c & n3482;
  assign n3484 = ~k & n3483;
  assign n3485 = ~j0 & n3201;
  assign n3486 = ~o & n3485;
  assign n3487 = ~c & n3486;
  assign n3488 = ~k & n3487;
  assign n3489 = ~d0 & n752;
  assign n3490 = l0 & n3489;
  assign n3491 = ~g0 & n3490;
  assign n3492 = j0 & n3491;
  assign n3493 = ~o & n3492;
  assign n3494 = ~c & n3493;
  assign n3495 = ~i0 & n3494;
  assign n3496 = ~d0 & n778;
  assign n3497 = l0 & n3496;
  assign n3498 = j0 & n3497;
  assign n3499 = ~o & n3498;
  assign n3500 = ~c & n3499;
  assign n3501 = ~i0 & n3500;
  assign n3502 = ~y & n736;
  assign n3503 = ~b0 & n3502;
  assign n3504 = ~c0 & n3503;
  assign n3505 = ~d0 & n3504;
  assign n3506 = l0 & n3505;
  assign n3507 = ~g0 & n3506;
  assign n3508 = ~j0 & n3507;
  assign n3509 = ~o & n3508;
  assign n3510 = ~c & n3509;
  assign n3511 = i0 & n3510;
  assign n3512 = ~y & n763;
  assign n3513 = ~b0 & n3512;
  assign n3514 = ~c0 & n3513;
  assign n3515 = ~d0 & n3514;
  assign n3516 = l0 & n3515;
  assign n3517 = ~j0 & n3516;
  assign n3518 = ~o & n3517;
  assign n3519 = ~c & n3518;
  assign n3520 = i0 & n3519;
  assign n3521 = ~y & n750;
  assign n3522 = ~b0 & n3521;
  assign n3523 = ~c0 & n3522;
  assign n3524 = ~d0 & n3523;
  assign n3525 = l0 & n3524;
  assign n3526 = ~g0 & n3525;
  assign n3527 = ~o & n3526;
  assign n3528 = ~c & n3527;
  assign n3529 = i0 & n3528;
  assign n3530 = ~y & n776;
  assign n3531 = ~b0 & n3530;
  assign n3532 = ~c0 & n3531;
  assign n3533 = ~d0 & n3532;
  assign n3534 = l0 & n3533;
  assign n3535 = ~o & n3534;
  assign n3536 = ~c & n3535;
  assign n3537 = i0 & n3536;
  assign n3538 = ~a0 & n3502;
  assign n3539 = ~b0 & n3538;
  assign n3540 = ~c0 & n3539;
  assign n3541 = ~d0 & n3540;
  assign n3542 = l0 & n3541;
  assign n3543 = ~g0 & n3542;
  assign n3544 = ~j0 & n3543;
  assign n3545 = ~o & n3544;
  assign n3546 = ~c & n3545;
  assign n3547 = ~a0 & n3512;
  assign n3548 = ~b0 & n3547;
  assign n3549 = ~c0 & n3548;
  assign n3550 = ~d0 & n3549;
  assign n3551 = l0 & n3550;
  assign n3552 = ~j0 & n3551;
  assign n3553 = ~o & n3552;
  assign n3554 = ~c & n3553;
  assign n3555 = ~d0 & n1157;
  assign n3556 = ~h0 & n3555;
  assign n3557 = l0 & n3556;
  assign n3558 = ~g0 & n3557;
  assign n3559 = j0 & n3558;
  assign n3560 = ~c & n3559;
  assign n3561 = ~i0 & n3560;
  assign n3562 = ~m & n3561;
  assign n3563 = ~d0 & n1169;
  assign n3564 = ~h0 & n3563;
  assign n3565 = l0 & n3564;
  assign n3566 = j0 & n3565;
  assign n3567 = ~c & n3566;
  assign n3568 = ~i0 & n3567;
  assign n3569 = ~m & n3568;
  assign n3570 = ~y & n920;
  assign n3571 = ~b0 & n3570;
  assign n3572 = ~c0 & n3571;
  assign n3573 = ~d0 & n3572;
  assign n3574 = ~h0 & n3573;
  assign n3575 = l0 & n3574;
  assign n3576 = ~g0 & n3575;
  assign n3577 = ~j0 & n3576;
  assign n3578 = ~c & n3577;
  assign n3579 = i0 & n3578;
  assign n3580 = ~m & n3579;
  assign n3581 = ~y & n934;
  assign n3582 = ~b0 & n3581;
  assign n3583 = ~c0 & n3582;
  assign n3584 = ~d0 & n3583;
  assign n3585 = ~h0 & n3584;
  assign n3586 = l0 & n3585;
  assign n3587 = ~j0 & n3586;
  assign n3588 = ~c & n3587;
  assign n3589 = i0 & n3588;
  assign n3590 = ~m & n3589;
  assign n3591 = ~y & n1155;
  assign n3592 = ~b0 & n3591;
  assign n3593 = ~c0 & n3592;
  assign n3594 = ~d0 & n3593;
  assign n3595 = ~h0 & n3594;
  assign n3596 = l0 & n3595;
  assign n3597 = ~g0 & n3596;
  assign n3598 = ~c & n3597;
  assign n3599 = i0 & n3598;
  assign n3600 = ~m & n3599;
  assign n3601 = ~y & n1167;
  assign n3602 = ~b0 & n3601;
  assign n3603 = ~c0 & n3602;
  assign n3604 = ~d0 & n3603;
  assign n3605 = ~h0 & n3604;
  assign n3606 = l0 & n3605;
  assign n3607 = ~c & n3606;
  assign n3608 = i0 & n3607;
  assign n3609 = ~m & n3608;
  assign n3610 = ~a0 & n3570;
  assign n3611 = ~b0 & n3610;
  assign n3612 = ~c0 & n3611;
  assign n3613 = ~d0 & n3612;
  assign n3614 = ~h0 & n3613;
  assign n3615 = l0 & n3614;
  assign n3616 = ~g0 & n3615;
  assign n3617 = ~j0 & n3616;
  assign n3618 = ~c & n3617;
  assign n3619 = ~m & n3618;
  assign n3620 = ~a0 & n3581;
  assign n3621 = ~b0 & n3620;
  assign n3622 = ~c0 & n3621;
  assign n3623 = ~d0 & n3622;
  assign n3624 = ~h0 & n3623;
  assign n3625 = l0 & n3624;
  assign n3626 = ~j0 & n3625;
  assign n3627 = ~c & n3626;
  assign n3628 = ~m & n3627;
  assign n3629 = ~u & n3397;
  assign n3630 = ~x & n3629;
  assign n3631 = ~y & n3630;
  assign n3632 = ~a0 & n3631;
  assign n3633 = ~b0 & n3632;
  assign n3634 = ~c0 & n3633;
  assign n3635 = d0 & n3634;
  assign n3636 = l0 & n3635;
  assign n3637 = ~g0 & n3636;
  assign n3638 = ~j0 & n3637;
  assign n3639 = ~o & n3638;
  assign n3640 = ~m & n3639;
  assign n3641 = ~u & n3411;
  assign n3642 = ~x & n3641;
  assign n3643 = ~y & n3642;
  assign n3644 = ~a0 & n3643;
  assign n3645 = ~b0 & n3644;
  assign n3646 = ~c0 & n3645;
  assign n3647 = d0 & n3646;
  assign n3648 = l0 & n3647;
  assign n3649 = ~j0 & n3648;
  assign n3650 = ~o & n3649;
  assign n3651 = ~m & n3650;
  assign n3652 = ~u & n3424;
  assign n3653 = ~x & n3652;
  assign n3654 = ~y & n3653;
  assign n3655 = ~a0 & n3654;
  assign n3656 = ~b0 & n3655;
  assign n3657 = ~c0 & n3656;
  assign n3658 = d0 & n3657;
  assign n3659 = l0 & n3658;
  assign n3660 = ~g0 & n3659;
  assign n3661 = ~o & n3660;
  assign n3662 = ~m & n3661;
  assign n3663 = ~u & n3437;
  assign n3664 = ~x & n3663;
  assign n3665 = ~y & n3664;
  assign n3666 = ~a0 & n3665;
  assign n3667 = ~b0 & n3666;
  assign n3668 = ~c0 & n3667;
  assign n3669 = d0 & n3668;
  assign n3670 = l0 & n3669;
  assign n3671 = ~o & n3670;
  assign n3672 = ~m & n3671;
  assign n3673 = ~r & n1089;
  assign n3674 = ~x & n3673;
  assign n3675 = ~b0 & n3674;
  assign n3676 = ~c0 & n3675;
  assign n3677 = ~d0 & n3676;
  assign n3678 = l0 & n3677;
  assign n3679 = ~g0 & n3678;
  assign n3680 = j0 & n3679;
  assign n3681 = ~o & n3680;
  assign n3682 = ~c & n3681;
  assign n3683 = ~i0 & n3682;
  assign n3684 = ~b & n3683;
  assign n3685 = ~r & n1101;
  assign n3686 = ~x & n3685;
  assign n3687 = ~b0 & n3686;
  assign n3688 = ~c0 & n3687;
  assign n3689 = ~d0 & n3688;
  assign n3690 = l0 & n3689;
  assign n3691 = j0 & n3690;
  assign n3692 = ~o & n3691;
  assign n3693 = ~c & n3692;
  assign n3694 = ~i0 & n3693;
  assign n3695 = ~b & n3694;
  assign n3696 = ~r & n853;
  assign n3697 = ~x & n3696;
  assign n3698 = ~y & n3697;
  assign n3699 = ~b0 & n3698;
  assign n3700 = ~c0 & n3699;
  assign n3701 = ~d0 & n3700;
  assign n3702 = l0 & n3701;
  assign n3703 = ~g0 & n3702;
  assign n3704 = ~j0 & n3703;
  assign n3705 = ~o & n3704;
  assign n3706 = ~c & n3705;
  assign n3707 = i0 & n3706;
  assign n3708 = ~b & n3707;
  assign n3709 = ~r & n867;
  assign n3710 = ~x & n3709;
  assign n3711 = ~y & n3710;
  assign n3712 = ~b0 & n3711;
  assign n3713 = ~c0 & n3712;
  assign n3714 = ~d0 & n3713;
  assign n3715 = l0 & n3714;
  assign n3716 = ~j0 & n3715;
  assign n3717 = ~o & n3716;
  assign n3718 = ~c & n3717;
  assign n3719 = i0 & n3718;
  assign n3720 = ~b & n3719;
  assign n3721 = ~y & n3674;
  assign n3722 = ~b0 & n3721;
  assign n3723 = ~c0 & n3722;
  assign n3724 = ~d0 & n3723;
  assign n3725 = l0 & n3724;
  assign n3726 = ~g0 & n3725;
  assign n3727 = ~o & n3726;
  assign n3728 = ~c & n3727;
  assign n3729 = i0 & n3728;
  assign n3730 = ~b & n3729;
  assign n3731 = ~y & n3686;
  assign n3732 = ~b0 & n3731;
  assign n3733 = ~c0 & n3732;
  assign n3734 = ~d0 & n3733;
  assign n3735 = l0 & n3734;
  assign n3736 = ~o & n3735;
  assign n3737 = ~c & n3736;
  assign n3738 = i0 & n3737;
  assign n3739 = ~b & n3738;
  assign n3740 = ~a0 & n3698;
  assign n3741 = ~b0 & n3740;
  assign n3742 = ~c0 & n3741;
  assign n3743 = ~d0 & n3742;
  assign n3744 = l0 & n3743;
  assign n3745 = ~g0 & n3744;
  assign n3746 = ~j0 & n3745;
  assign n3747 = ~o & n3746;
  assign n3748 = ~c & n3747;
  assign n3749 = ~b & n3748;
  assign n3750 = ~a0 & n3711;
  assign n3751 = ~b0 & n3750;
  assign n3752 = ~c0 & n3751;
  assign n3753 = ~d0 & n3752;
  assign n3754 = l0 & n3753;
  assign n3755 = ~j0 & n3754;
  assign n3756 = ~o & n3755;
  assign n3757 = ~c & n3756;
  assign n3758 = ~b & n3757;
  assign n3759 = ~d0 & n1092;
  assign n3760 = l0 & n3759;
  assign n3761 = ~g0 & n3760;
  assign n3762 = j0 & n3761;
  assign n3763 = ~o & n3762;
  assign n3764 = ~c & n3763;
  assign n3765 = ~i0 & n3764;
  assign n3766 = ~m & n3765;
  assign n3767 = ~d0 & n1104;
  assign n3768 = l0 & n3767;
  assign n3769 = j0 & n3768;
  assign n3770 = ~o & n3769;
  assign n3771 = ~c & n3770;
  assign n3772 = ~i0 & n3771;
  assign n3773 = ~m & n3772;
  assign n3774 = ~y & n854;
  assign n3775 = ~b0 & n3774;
  assign n3776 = ~c0 & n3775;
  assign n3777 = ~d0 & n3776;
  assign n3778 = l0 & n3777;
  assign n3779 = ~g0 & n3778;
  assign n3780 = ~j0 & n3779;
  assign n3781 = ~o & n3780;
  assign n3782 = ~c & n3781;
  assign n3783 = i0 & n3782;
  assign n3784 = ~m & n3783;
  assign n3785 = ~y & n868;
  assign n3786 = ~b0 & n3785;
  assign n3787 = ~c0 & n3786;
  assign n3788 = ~d0 & n3787;
  assign n3789 = l0 & n3788;
  assign n3790 = ~j0 & n3789;
  assign n3791 = ~o & n3790;
  assign n3792 = ~c & n3791;
  assign n3793 = i0 & n3792;
  assign n3794 = ~m & n3793;
  assign n3795 = ~y & n1090;
  assign n3796 = ~b0 & n3795;
  assign n3797 = ~c0 & n3796;
  assign n3798 = ~d0 & n3797;
  assign n3799 = l0 & n3798;
  assign n3800 = ~g0 & n3799;
  assign n3801 = ~o & n3800;
  assign n3802 = ~c & n3801;
  assign n3803 = i0 & n3802;
  assign n3804 = ~m & n3803;
  assign n3805 = ~y & n1102;
  assign n3806 = ~b0 & n3805;
  assign n3807 = ~c0 & n3806;
  assign n3808 = ~d0 & n3807;
  assign n3809 = l0 & n3808;
  assign n3810 = ~o & n3809;
  assign n3811 = ~c & n3810;
  assign n3812 = i0 & n3811;
  assign n3813 = ~m & n3812;
  assign n3814 = ~a0 & n3774;
  assign n3815 = ~b0 & n3814;
  assign n3816 = ~c0 & n3815;
  assign n3817 = ~d0 & n3816;
  assign n3818 = l0 & n3817;
  assign n3819 = ~g0 & n3818;
  assign n3820 = ~j0 & n3819;
  assign n3821 = ~o & n3820;
  assign n3822 = ~c & n3821;
  assign n3823 = ~m & n3822;
  assign n3824 = ~a0 & n3785;
  assign n3825 = ~b0 & n3824;
  assign n3826 = ~c0 & n3825;
  assign n3827 = ~d0 & n3826;
  assign n3828 = l0 & n3827;
  assign n3829 = ~j0 & n3828;
  assign n3830 = ~o & n3829;
  assign n3831 = ~c & n3830;
  assign n3832 = ~m & n3831;
  assign n3833 = ~a & ~n;
  assign n3834 = ~q & n3833;
  assign n3835 = ~u & n3834;
  assign n3836 = ~x & n3835;
  assign n3837 = ~y & n3836;
  assign n3838 = ~a0 & n3837;
  assign n3839 = ~b0 & n3838;
  assign n3840 = ~c0 & n3839;
  assign n3841 = ~h0 & n3840;
  assign n3842 = l0 & n3841;
  assign n3843 = ~g0 & n3842;
  assign n3844 = ~j0 & n3843;
  assign n3845 = ~m & n3844;
  assign n3846 = ~e0 & n3845;
  assign n3847 = ~a & ~i;
  assign n3848 = ~n & n3847;
  assign n3849 = ~q & n3848;
  assign n3850 = ~u & n3849;
  assign n3851 = ~x & n3850;
  assign n3852 = ~y & n3851;
  assign n3853 = ~a0 & n3852;
  assign n3854 = ~b0 & n3853;
  assign n3855 = ~c0 & n3854;
  assign n3856 = ~h0 & n3855;
  assign n3857 = l0 & n3856;
  assign n3858 = ~j0 & n3857;
  assign n3859 = ~m & n3858;
  assign n3860 = ~e0 & n3859;
  assign n3861 = ~a & ~h;
  assign n3862 = ~n & n3861;
  assign n3863 = ~q & n3862;
  assign n3864 = ~u & n3863;
  assign n3865 = ~x & n3864;
  assign n3866 = ~y & n3865;
  assign n3867 = ~a0 & n3866;
  assign n3868 = ~b0 & n3867;
  assign n3869 = ~c0 & n3868;
  assign n3870 = ~h0 & n3869;
  assign n3871 = l0 & n3870;
  assign n3872 = ~g0 & n3871;
  assign n3873 = ~m & n3872;
  assign n3874 = ~e0 & n3873;
  assign n3875 = ~i & n3861;
  assign n3876 = ~n & n3875;
  assign n3877 = ~q & n3876;
  assign n3878 = ~u & n3877;
  assign n3879 = ~x & n3878;
  assign n3880 = ~y & n3879;
  assign n3881 = ~a0 & n3880;
  assign n3882 = ~b0 & n3881;
  assign n3883 = ~c0 & n3882;
  assign n3884 = ~h0 & n3883;
  assign n3885 = l0 & n3884;
  assign n3886 = ~m & n3885;
  assign n3887 = ~e0 & n3886;
  assign n3888 = ~r & n3834;
  assign n3889 = ~u & n3888;
  assign n3890 = ~x & n3889;
  assign n3891 = ~y & n3890;
  assign n3892 = ~a0 & n3891;
  assign n3893 = ~b0 & n3892;
  assign n3894 = ~c0 & n3893;
  assign n3895 = ~h0 & n3894;
  assign n3896 = l0 & n3895;
  assign n3897 = ~g0 & n3896;
  assign n3898 = ~j0 & n3897;
  assign n3899 = ~e0 & n3898;
  assign n3900 = ~r & n3849;
  assign n3901 = ~u & n3900;
  assign n3902 = ~x & n3901;
  assign n3903 = ~y & n3902;
  assign n3904 = ~a0 & n3903;
  assign n3905 = ~b0 & n3904;
  assign n3906 = ~c0 & n3905;
  assign n3907 = ~h0 & n3906;
  assign n3908 = l0 & n3907;
  assign n3909 = ~j0 & n3908;
  assign n3910 = ~e0 & n3909;
  assign n3911 = ~r & n3863;
  assign n3912 = ~u & n3911;
  assign n3913 = ~x & n3912;
  assign n3914 = ~y & n3913;
  assign n3915 = ~a0 & n3914;
  assign n3916 = ~b0 & n3915;
  assign n3917 = ~c0 & n3916;
  assign n3918 = ~h0 & n3917;
  assign n3919 = l0 & n3918;
  assign n3920 = ~g0 & n3919;
  assign n3921 = ~e0 & n3920;
  assign n3922 = ~r & n3877;
  assign n3923 = ~u & n3922;
  assign n3924 = ~x & n3923;
  assign n3925 = ~y & n3924;
  assign n3926 = ~a0 & n3925;
  assign n3927 = ~b0 & n3926;
  assign n3928 = ~c0 & n3927;
  assign n3929 = ~h0 & n3928;
  assign n3930 = l0 & n3929;
  assign n3931 = ~e0 & n3930;
  assign n3932 = ~d0 & n1311;
  assign n3933 = ~h0 & n3932;
  assign n3934 = l0 & n3933;
  assign n3935 = ~g0 & n3934;
  assign n3936 = j0 & n3935;
  assign n3937 = ~i0 & n3936;
  assign n3938 = ~m & n3937;
  assign n3939 = ~e0 & n3938;
  assign n3940 = f0 & n3939;
  assign n3941 = ~y & n1309;
  assign n3942 = ~b0 & n3941;
  assign n3943 = ~c0 & n3942;
  assign n3944 = ~d0 & n3943;
  assign n3945 = ~h0 & n3944;
  assign n3946 = l0 & n3945;
  assign n3947 = ~g0 & n3946;
  assign n3948 = i0 & n3947;
  assign n3949 = ~m & n3948;
  assign n3950 = ~e0 & n3949;
  assign n3951 = f0 & n3950;
  assign n3952 = ~a0 & n3941;
  assign n3953 = ~b0 & n3952;
  assign n3954 = ~c0 & n3953;
  assign n3955 = ~d0 & n3954;
  assign n3956 = ~h0 & n3955;
  assign n3957 = l0 & n3956;
  assign n3958 = ~g0 & n3957;
  assign n3959 = ~m & n3958;
  assign n3960 = ~e0 & n3959;
  assign n3961 = f0 & n3960;
  assign n3962 = ~d0 & n2008;
  assign n3963 = ~h0 & n3962;
  assign n3964 = l0 & n3963;
  assign n3965 = ~g0 & n3964;
  assign n3966 = j0 & n3965;
  assign n3967 = ~i0 & n3966;
  assign n3968 = ~e0 & n3967;
  assign n3969 = f0 & n3968;
  assign n3970 = ~y & n2006;
  assign n3971 = ~b0 & n3970;
  assign n3972 = ~c0 & n3971;
  assign n3973 = ~d0 & n3972;
  assign n3974 = ~h0 & n3973;
  assign n3975 = l0 & n3974;
  assign n3976 = ~g0 & n3975;
  assign n3977 = i0 & n3976;
  assign n3978 = ~e0 & n3977;
  assign n3979 = f0 & n3978;
  assign n3980 = ~a0 & n3970;
  assign n3981 = ~b0 & n3980;
  assign n3982 = ~c0 & n3981;
  assign n3983 = ~d0 & n3982;
  assign n3984 = ~h0 & n3983;
  assign n3985 = l0 & n3984;
  assign n3986 = ~g0 & n3985;
  assign n3987 = ~e0 & n3986;
  assign n3988 = f0 & n3987;
  assign n3989 = ~h0 & n1674;
  assign n3990 = l0 & n3989;
  assign n3991 = j0 & n3990;
  assign n3992 = ~i0 & n3991;
  assign n3993 = ~m & n3992;
  assign n3994 = ~e0 & n3993;
  assign n3995 = ~y & n1323;
  assign n3996 = ~b0 & n3995;
  assign n3997 = ~c0 & n3996;
  assign n3998 = ~d0 & n3997;
  assign n3999 = ~h0 & n3998;
  assign n4000 = l0 & n3999;
  assign n4001 = ~j0 & n4000;
  assign n4002 = i0 & n4001;
  assign n4003 = ~m & n4002;
  assign n4004 = ~e0 & n4003;
  assign n4005 = ~y & n1658;
  assign n4006 = ~b0 & n4005;
  assign n4007 = ~c0 & n4006;
  assign n4008 = ~d0 & n4007;
  assign n4009 = ~h0 & n4008;
  assign n4010 = l0 & n4009;
  assign n4011 = i0 & n4010;
  assign n4012 = ~m & n4011;
  assign n4013 = ~e0 & n4012;
  assign n4014 = ~a & ~q;
  assign n4015 = ~u & n4014;
  assign n4016 = ~x & n4015;
  assign n4017 = ~y & n4016;
  assign n4018 = ~a0 & n4017;
  assign n4019 = ~b0 & n4018;
  assign n4020 = ~c0 & n4019;
  assign n4021 = l0 & n4020;
  assign n4022 = ~g0 & n4021;
  assign n4023 = ~j0 & n4022;
  assign n4024 = ~o & n4023;
  assign n4025 = ~m & n4024;
  assign n4026 = ~e0 & n4025;
  assign n4027 = ~q & n3847;
  assign n4028 = ~u & n4027;
  assign n4029 = ~x & n4028;
  assign n4030 = ~y & n4029;
  assign n4031 = ~a0 & n4030;
  assign n4032 = ~b0 & n4031;
  assign n4033 = ~c0 & n4032;
  assign n4034 = l0 & n4033;
  assign n4035 = ~j0 & n4034;
  assign n4036 = ~o & n4035;
  assign n4037 = ~m & n4036;
  assign n4038 = ~e0 & n4037;
  assign n4039 = ~q & n3861;
  assign n4040 = ~u & n4039;
  assign n4041 = ~x & n4040;
  assign n4042 = ~y & n4041;
  assign n4043 = ~a0 & n4042;
  assign n4044 = ~b0 & n4043;
  assign n4045 = ~c0 & n4044;
  assign n4046 = l0 & n4045;
  assign n4047 = ~g0 & n4046;
  assign n4048 = ~o & n4047;
  assign n4049 = ~m & n4048;
  assign n4050 = ~e0 & n4049;
  assign n4051 = ~q & n3875;
  assign n4052 = ~u & n4051;
  assign n4053 = ~x & n4052;
  assign n4054 = ~y & n4053;
  assign n4055 = ~a0 & n4054;
  assign n4056 = ~b0 & n4055;
  assign n4057 = ~c0 & n4056;
  assign n4058 = l0 & n4057;
  assign n4059 = ~o & n4058;
  assign n4060 = ~m & n4059;
  assign n4061 = ~e0 & n4060;
  assign n4062 = ~a0 & n3995;
  assign n4063 = ~b0 & n4062;
  assign n4064 = ~c0 & n4063;
  assign n4065 = ~d0 & n4064;
  assign n4066 = ~h0 & n4065;
  assign n4067 = l0 & n4066;
  assign n4068 = ~j0 & n4067;
  assign n4069 = ~m & n4068;
  assign n4070 = ~e0 & n4069;
  assign n4071 = ~h0 & n1759;
  assign n4072 = l0 & n4071;
  assign n4073 = j0 & n4072;
  assign n4074 = ~i0 & n4073;
  assign n4075 = ~e0 & n4074;
  assign n4076 = ~y & n1369;
  assign n4077 = ~b0 & n4076;
  assign n4078 = ~c0 & n4077;
  assign n4079 = ~d0 & n4078;
  assign n4080 = ~h0 & n4079;
  assign n4081 = l0 & n4080;
  assign n4082 = ~j0 & n4081;
  assign n4083 = i0 & n4082;
  assign n4084 = ~e0 & n4083;
  assign n4085 = ~y & n1756;
  assign n4086 = ~b0 & n4085;
  assign n4087 = ~c0 & n4086;
  assign n4088 = ~d0 & n4087;
  assign n4089 = ~h0 & n4088;
  assign n4090 = l0 & n4089;
  assign n4091 = i0 & n4090;
  assign n4092 = ~e0 & n4091;
  assign n4093 = ~r & n4014;
  assign n4094 = ~u & n4093;
  assign n4095 = ~x & n4094;
  assign n4096 = ~y & n4095;
  assign n4097 = ~a0 & n4096;
  assign n4098 = ~b0 & n4097;
  assign n4099 = ~c0 & n4098;
  assign n4100 = l0 & n4099;
  assign n4101 = ~g0 & n4100;
  assign n4102 = ~j0 & n4101;
  assign n4103 = ~o & n4102;
  assign n4104 = ~e0 & n4103;
  assign n4105 = ~r & n4027;
  assign n4106 = ~u & n4105;
  assign n4107 = ~x & n4106;
  assign n4108 = ~y & n4107;
  assign n4109 = ~a0 & n4108;
  assign n4110 = ~b0 & n4109;
  assign n4111 = ~c0 & n4110;
  assign n4112 = l0 & n4111;
  assign n4113 = ~j0 & n4112;
  assign n4114 = ~o & n4113;
  assign n4115 = ~e0 & n4114;
  assign n4116 = ~r & n4039;
  assign n4117 = ~u & n4116;
  assign n4118 = ~x & n4117;
  assign n4119 = ~y & n4118;
  assign n4120 = ~a0 & n4119;
  assign n4121 = ~b0 & n4120;
  assign n4122 = ~c0 & n4121;
  assign n4123 = l0 & n4122;
  assign n4124 = ~g0 & n4123;
  assign n4125 = ~o & n4124;
  assign n4126 = ~e0 & n4125;
  assign n4127 = ~r & n4051;
  assign n4128 = ~u & n4127;
  assign n4129 = ~x & n4128;
  assign n4130 = ~y & n4129;
  assign n4131 = ~a0 & n4130;
  assign n4132 = ~b0 & n4131;
  assign n4133 = ~c0 & n4132;
  assign n4134 = l0 & n4133;
  assign n4135 = ~o & n4134;
  assign n4136 = ~e0 & n4135;
  assign n4137 = ~a0 & n4076;
  assign n4138 = ~b0 & n4137;
  assign n4139 = ~c0 & n4138;
  assign n4140 = ~d0 & n4139;
  assign n4141 = ~h0 & n4140;
  assign n4142 = l0 & n4141;
  assign n4143 = ~j0 & n4142;
  assign n4144 = ~e0 & n4143;
  assign n4145 = ~d0 & n1268;
  assign n4146 = l0 & n4145;
  assign n4147 = ~g0 & n4146;
  assign n4148 = j0 & n4147;
  assign n4149 = ~o & n4148;
  assign n4150 = ~i0 & n4149;
  assign n4151 = ~m & n4150;
  assign n4152 = ~e0 & n4151;
  assign n4153 = f0 & n4152;
  assign n4154 = ~y & n1266;
  assign n4155 = ~b0 & n4154;
  assign n4156 = ~c0 & n4155;
  assign n4157 = ~d0 & n4156;
  assign n4158 = l0 & n4157;
  assign n4159 = ~g0 & n4158;
  assign n4160 = ~o & n4159;
  assign n4161 = i0 & n4160;
  assign n4162 = ~m & n4161;
  assign n4163 = ~e0 & n4162;
  assign n4164 = f0 & n4163;
  assign n4165 = ~a0 & n4154;
  assign n4166 = ~b0 & n4165;
  assign n4167 = ~c0 & n4166;
  assign n4168 = ~d0 & n4167;
  assign n4169 = l0 & n4168;
  assign n4170 = ~g0 & n4169;
  assign n4171 = ~o & n4170;
  assign n4172 = ~m & n4171;
  assign n4173 = ~e0 & n4172;
  assign n4174 = f0 & n4173;
  assign n4175 = ~d0 & n1999;
  assign n4176 = l0 & n4175;
  assign n4177 = ~g0 & n4176;
  assign n4178 = j0 & n4177;
  assign n4179 = ~o & n4178;
  assign n4180 = ~i0 & n4179;
  assign n4181 = ~e0 & n4180;
  assign n4182 = f0 & n4181;
  assign n4183 = ~y & n1997;
  assign n4184 = ~b0 & n4183;
  assign n4185 = ~c0 & n4184;
  assign n4186 = ~d0 & n4185;
  assign n4187 = l0 & n4186;
  assign n4188 = ~g0 & n4187;
  assign n4189 = ~o & n4188;
  assign n4190 = i0 & n4189;
  assign n4191 = ~e0 & n4190;
  assign n4192 = f0 & n4191;
  assign n4193 = ~a0 & n4183;
  assign n4194 = ~b0 & n4193;
  assign n4195 = ~c0 & n4194;
  assign n4196 = ~d0 & n4195;
  assign n4197 = l0 & n4196;
  assign n4198 = ~g0 & n4197;
  assign n4199 = ~o & n4198;
  assign n4200 = ~e0 & n4199;
  assign n4201 = f0 & n4200;
  assign n4202 = l0 & n1611;
  assign n4203 = j0 & n4202;
  assign n4204 = ~o & n4203;
  assign n4205 = ~i0 & n4204;
  assign n4206 = ~m & n4205;
  assign n4207 = ~e0 & n4206;
  assign n4208 = ~y & n1280;
  assign n4209 = ~b0 & n4208;
  assign n4210 = ~c0 & n4209;
  assign n4211 = ~d0 & n4210;
  assign n4212 = l0 & n4211;
  assign n4213 = ~j0 & n4212;
  assign n4214 = ~o & n4213;
  assign n4215 = i0 & n4214;
  assign n4216 = ~m & n4215;
  assign n4217 = ~e0 & n4216;
  assign n4218 = ~y & n1593;
  assign n4219 = ~b0 & n4218;
  assign n4220 = ~c0 & n4219;
  assign n4221 = ~d0 & n4220;
  assign n4222 = l0 & n4221;
  assign n4223 = ~o & n4222;
  assign n4224 = i0 & n4223;
  assign n4225 = ~m & n4224;
  assign n4226 = ~e0 & n4225;
  assign n4227 = ~a0 & n4208;
  assign n4228 = ~b0 & n4227;
  assign n4229 = ~c0 & n4228;
  assign n4230 = ~d0 & n4229;
  assign n4231 = l0 & n4230;
  assign n4232 = ~j0 & n4231;
  assign n4233 = ~o & n4232;
  assign n4234 = ~m & n4233;
  assign n4235 = ~e0 & n4234;
  assign n4236 = l0 & n1717;
  assign n4237 = j0 & n4236;
  assign n4238 = ~o & n4237;
  assign n4239 = ~i0 & n4238;
  assign n4240 = ~e0 & n4239;
  assign n4241 = ~y & n1350;
  assign n4242 = ~b0 & n4241;
  assign n4243 = ~c0 & n4242;
  assign n4244 = ~d0 & n4243;
  assign n4245 = l0 & n4244;
  assign n4246 = ~j0 & n4245;
  assign n4247 = ~o & n4246;
  assign n4248 = i0 & n4247;
  assign n4249 = ~e0 & n4248;
  assign n4250 = ~y & n1714;
  assign n4251 = ~b0 & n4250;
  assign n4252 = ~c0 & n4251;
  assign n4253 = ~d0 & n4252;
  assign n4254 = l0 & n4253;
  assign n4255 = ~o & n4254;
  assign n4256 = i0 & n4255;
  assign n4257 = ~e0 & n4256;
  assign n4258 = ~a0 & n4241;
  assign n4259 = ~b0 & n4258;
  assign n4260 = ~c0 & n4259;
  assign n4261 = ~d0 & n4260;
  assign n4262 = l0 & n4261;
  assign n4263 = ~j0 & n4262;
  assign n4264 = ~o & n4263;
  assign n4265 = ~e0 & n4264;
  assign n4266 = ~q & u;
  assign n4267 = ~x & n4266;
  assign n4268 = ~b0 & n4267;
  assign n4269 = ~c0 & n4268;
  assign n4270 = h0 & n4269;
  assign n4271 = j0 & n4270;
  assign n4272 = ~o & n4271;
  assign n4273 = ~i0 & n4272;
  assign n4274 = ~m & n4273;
  assign n4275 = z & n4274;
  assign n4276 = h0 & n3932;
  assign n4277 = j0 & n4276;
  assign n4278 = ~i0 & n4277;
  assign n4279 = ~m & n4278;
  assign n4280 = z & n4279;
  assign n4281 = u & n42;
  assign n4282 = ~x & n4281;
  assign n4283 = ~b0 & n4282;
  assign n4284 = ~c0 & n4283;
  assign n4285 = h0 & n4284;
  assign n4286 = j0 & n4285;
  assign n4287 = ~i0 & n4286;
  assign n4288 = ~m & n4287;
  assign n4289 = z & n4288;
  assign n4290 = ~y & n4267;
  assign n4291 = ~b0 & n4290;
  assign n4292 = ~c0 & n4291;
  assign n4293 = h0 & n4292;
  assign n4294 = ~o & n4293;
  assign n4295 = i0 & n4294;
  assign n4296 = ~m & n4295;
  assign n4297 = z & n4296;
  assign n4298 = h0 & n3944;
  assign n4299 = i0 & n4298;
  assign n4300 = ~m & n4299;
  assign n4301 = z & n4300;
  assign n4302 = ~y & n4282;
  assign n4303 = ~b0 & n4302;
  assign n4304 = ~c0 & n4303;
  assign n4305 = h0 & n4304;
  assign n4306 = i0 & n4305;
  assign n4307 = ~m & n4306;
  assign n4308 = z & n4307;
  assign n4309 = u & n1996;
  assign n4310 = ~x & n4309;
  assign n4311 = ~b0 & n4310;
  assign n4312 = ~c0 & n4311;
  assign n4313 = h0 & n4312;
  assign n4314 = j0 & n4313;
  assign n4315 = ~o & n4314;
  assign n4316 = ~i0 & n4315;
  assign n4317 = z & n4316;
  assign n4318 = h0 & n3962;
  assign n4319 = j0 & n4318;
  assign n4320 = ~i0 & n4319;
  assign n4321 = z & n4320;
  assign n4322 = ~x & n235;
  assign n4323 = ~b0 & n4322;
  assign n4324 = ~c0 & n4323;
  assign n4325 = h0 & n4324;
  assign n4326 = j0 & n4325;
  assign n4327 = ~i0 & n4326;
  assign n4328 = z & n4327;
  assign n4329 = ~y & n4310;
  assign n4330 = ~b0 & n4329;
  assign n4331 = ~c0 & n4330;
  assign n4332 = h0 & n4331;
  assign n4333 = ~o & n4332;
  assign n4334 = i0 & n4333;
  assign n4335 = z & n4334;
  assign n4336 = h0 & n3973;
  assign n4337 = i0 & n4336;
  assign n4338 = z & n4337;
  assign n4339 = ~y & n4322;
  assign n4340 = ~b0 & n4339;
  assign n4341 = ~c0 & n4340;
  assign n4342 = h0 & n4341;
  assign n4343 = i0 & n4342;
  assign n4344 = z & n4343;
  assign n4345 = ~y & ~a0;
  assign n4346 = ~c0 & n4345;
  assign n4347 = ~d0 & n4346;
  assign n4348 = l0 & n4347;
  assign n4349 = ~g0 & n4348;
  assign n4350 = ~j0 & n4349;
  assign n4351 = ~o & n4350;
  assign n4352 = ~i0 & n4351;
  assign n4353 = ~e0 & n4352;
  assign n4354 = ~f0 & n4353;
  assign n4355 = ~h0 & n4347;
  assign n4356 = l0 & n4355;
  assign n4357 = ~g0 & n4356;
  assign n4358 = ~j0 & n4357;
  assign n4359 = ~i0 & n4358;
  assign n4360 = ~e0 & n4359;
  assign n4361 = ~f0 & n4360;
  assign n4362 = ~c0 & n167;
  assign n4363 = ~d0 & n4362;
  assign n4364 = l0 & n4363;
  assign n4365 = ~g0 & n4364;
  assign n4366 = ~j0 & n4365;
  assign n4367 = ~o & n4366;
  assign n4368 = i0 & n4367;
  assign n4369 = ~e0 & n4368;
  assign n4370 = ~f0 & n4369;
  assign n4371 = ~y & n2194;
  assign n4372 = ~c0 & n4371;
  assign n4373 = ~d0 & n4372;
  assign n4374 = l0 & n4373;
  assign n4375 = ~g0 & n4374;
  assign n4376 = ~o & n4375;
  assign n4377 = i0 & n4376;
  assign n4378 = ~e0 & n4377;
  assign n4379 = ~f0 & n4378;
  assign n4380 = ~h0 & n4363;
  assign n4381 = l0 & n4380;
  assign n4382 = ~g0 & n4381;
  assign n4383 = ~j0 & n4382;
  assign n4384 = i0 & n4383;
  assign n4385 = ~e0 & n4384;
  assign n4386 = ~f0 & n4385;
  assign n4387 = ~h0 & n4373;
  assign n4388 = l0 & n4387;
  assign n4389 = ~g0 & n4388;
  assign n4390 = i0 & n4389;
  assign n4391 = ~e0 & n4390;
  assign n4392 = ~f0 & n4391;
  assign n4393 = h & ~q;
  assign n4394 = ~x & n4393;
  assign n4395 = ~b0 & n4394;
  assign n4396 = ~c0 & n4395;
  assign n4397 = ~d0 & n4396;
  assign n4398 = j0 & n4397;
  assign n4399 = ~o & n4398;
  assign n4400 = ~i0 & n4399;
  assign n4401 = ~m & n4400;
  assign n4402 = f0 & n4401;
  assign n4403 = u & n4393;
  assign n4404 = ~x & n4403;
  assign n4405 = ~b0 & n4404;
  assign n4406 = ~c0 & n4405;
  assign n4407 = j0 & n4406;
  assign n4408 = ~o & n4407;
  assign n4409 = ~i0 & n4408;
  assign n4410 = ~m & n4409;
  assign n4411 = f0 & n4410;
  assign n4412 = j0 & n1459;
  assign n4413 = ~i0 & n4412;
  assign n4414 = ~m & n4413;
  assign n4415 = f0 & n4414;
  assign n4416 = u & n1434;
  assign n4417 = ~x & n4416;
  assign n4418 = ~b0 & n4417;
  assign n4419 = ~c0 & n4418;
  assign n4420 = j0 & n4419;
  assign n4421 = ~i0 & n4420;
  assign n4422 = ~m & n4421;
  assign n4423 = f0 & n4422;
  assign n4424 = ~y & n4394;
  assign n4425 = ~b0 & n4424;
  assign n4426 = ~c0 & n4425;
  assign n4427 = ~d0 & n4426;
  assign n4428 = ~o & n4427;
  assign n4429 = i0 & n4428;
  assign n4430 = ~m & n4429;
  assign n4431 = f0 & n4430;
  assign n4432 = ~y & n4404;
  assign n4433 = ~b0 & n4432;
  assign n4434 = ~c0 & n4433;
  assign n4435 = ~o & n4434;
  assign n4436 = i0 & n4435;
  assign n4437 = ~m & n4436;
  assign n4438 = f0 & n4437;
  assign n4439 = ~y & n1435;
  assign n4440 = ~b0 & n4439;
  assign n4441 = ~c0 & n4440;
  assign n4442 = ~d0 & n4441;
  assign n4443 = i0 & n4442;
  assign n4444 = ~m & n4443;
  assign n4445 = f0 & n4444;
  assign n4446 = ~y & n4417;
  assign n4447 = ~b0 & n4446;
  assign n4448 = ~c0 & n4447;
  assign n4449 = i0 & n4448;
  assign n4450 = ~m & n4449;
  assign n4451 = f0 & n4450;
  assign n4452 = ~r & n4393;
  assign n4453 = ~x & n4452;
  assign n4454 = ~b0 & n4453;
  assign n4455 = ~c0 & n4454;
  assign n4456 = ~d0 & n4455;
  assign n4457 = j0 & n4456;
  assign n4458 = ~o & n4457;
  assign n4459 = ~i0 & n4458;
  assign n4460 = f0 & n4459;
  assign n4461 = u & n4452;
  assign n4462 = ~x & n4461;
  assign n4463 = ~b0 & n4462;
  assign n4464 = ~c0 & n4463;
  assign n4465 = j0 & n4464;
  assign n4466 = ~o & n4465;
  assign n4467 = ~i0 & n4466;
  assign n4468 = f0 & n4467;
  assign n4469 = j0 & n1520;
  assign n4470 = ~i0 & n4469;
  assign n4471 = f0 & n4470;
  assign n4472 = u & n1499;
  assign n4473 = ~x & n4472;
  assign n4474 = ~b0 & n4473;
  assign n4475 = ~c0 & n4474;
  assign n4476 = j0 & n4475;
  assign n4477 = ~i0 & n4476;
  assign n4478 = f0 & n4477;
  assign n4479 = ~y & n4453;
  assign n4480 = ~b0 & n4479;
  assign n4481 = ~c0 & n4480;
  assign n4482 = ~d0 & n4481;
  assign n4483 = ~o & n4482;
  assign n4484 = i0 & n4483;
  assign n4485 = f0 & n4484;
  assign n4486 = ~y & n4462;
  assign n4487 = ~b0 & n4486;
  assign n4488 = ~c0 & n4487;
  assign n4489 = ~o & n4488;
  assign n4490 = i0 & n4489;
  assign n4491 = f0 & n4490;
  assign n4492 = ~y & n1500;
  assign n4493 = ~b0 & n4492;
  assign n4494 = ~c0 & n4493;
  assign n4495 = ~d0 & n4494;
  assign n4496 = i0 & n4495;
  assign n4497 = f0 & n4496;
  assign n4498 = ~y & n4473;
  assign n4499 = ~b0 & n4498;
  assign n4500 = ~c0 & n4499;
  assign n4501 = i0 & n4500;
  assign n4502 = f0 & n4501;
  assign n4503 = ~u & n1996;
  assign n4504 = ~x & n4503;
  assign n4505 = ~y & n4504;
  assign n4506 = ~a0 & n4505;
  assign n4507 = ~b0 & n4506;
  assign n4508 = ~c0 & n4507;
  assign n4509 = d0 & n4508;
  assign n4510 = ~o & n4509;
  assign n4511 = c & n4510;
  assign n4512 = ~u & n43;
  assign n4513 = ~x & n4512;
  assign n4514 = ~y & n4513;
  assign n4515 = ~a0 & n4514;
  assign n4516 = ~b0 & n4515;
  assign n4517 = ~c0 & n4516;
  assign n4518 = d0 & n4517;
  assign n4519 = c & n4518;
  assign n4520 = j0 & n1983;
  assign n4521 = ~o & n4520;
  assign n4522 = ~i0 & n4521;
  assign n4523 = ~m & n4522;
  assign n4524 = v & n4523;
  assign n4525 = j0 & n1990;
  assign n4526 = ~i0 & n4525;
  assign n4527 = ~m & n4526;
  assign n4528 = v & n4527;
  assign n4529 = d0 & n4156;
  assign n4530 = ~o & n4529;
  assign n4531 = i0 & n4530;
  assign n4532 = ~m & n4531;
  assign n4533 = v & n4532;
  assign n4534 = d0 & n3943;
  assign n4535 = i0 & n4534;
  assign n4536 = ~m & n4535;
  assign n4537 = v & n4536;
  assign n4538 = j0 & n2000;
  assign n4539 = ~o & n4538;
  assign n4540 = ~i0 & n4539;
  assign n4541 = v & n4540;
  assign n4542 = j0 & n2009;
  assign n4543 = ~i0 & n4542;
  assign n4544 = v & n4543;
  assign n4545 = d0 & n4185;
  assign n4546 = ~o & n4545;
  assign n4547 = i0 & n4546;
  assign n4548 = v & n4547;
  assign n4549 = d0 & n3972;
  assign n4550 = i0 & n4549;
  assign n4551 = v & n4550;
  assign n4552 = u & ~y;
  assign n4553 = ~a0 & n4552;
  assign n4554 = ~c0 & n4553;
  assign n4555 = h0 & n4554;
  assign n4556 = ~g0 & n4555;
  assign n4557 = ~i0 & n4556;
  assign n4558 = ~e0 & n4557;
  assign n4559 = ~f0 & n4558;
  assign n4560 = z & n4559;
  assign n4561 = u & ~x;
  assign n4562 = ~y & n4561;
  assign n4563 = ~c0 & n4562;
  assign n4564 = h0 & n4563;
  assign n4565 = ~g0 & n4564;
  assign n4566 = i0 & n4565;
  assign n4567 = ~e0 & n4566;
  assign n4568 = ~f0 & n4567;
  assign n4569 = z & n4568;
  assign n4570 = h0 & n3954;
  assign n4571 = ~m & n4570;
  assign n4572 = z & n4571;
  assign n4573 = h0 & n3982;
  assign n4574 = z & n4573;
  assign n4575 = l0 & n2221;
  assign n4576 = ~g0 & n4575;
  assign n4577 = j0 & n4576;
  assign n4578 = ~o & n4577;
  assign n4579 = ~i0 & n4578;
  assign n4580 = ~e0 & n4579;
  assign n4581 = ~f0 & n4580;
  assign n4582 = ~h0 & n2221;
  assign n4583 = l0 & n4582;
  assign n4584 = ~g0 & n4583;
  assign n4585 = j0 & n4584;
  assign n4586 = ~i0 & n4585;
  assign n4587 = ~e0 & n4586;
  assign n4588 = ~f0 & n4587;
  assign n4589 = ~a0 & n4424;
  assign n4590 = ~b0 & n4589;
  assign n4591 = ~c0 & n4590;
  assign n4592 = ~o & n4591;
  assign n4593 = ~m & n4592;
  assign n4594 = f0 & n4593;
  assign n4595 = ~a0 & n4439;
  assign n4596 = ~b0 & n4595;
  assign n4597 = ~c0 & n4596;
  assign n4598 = ~m & n4597;
  assign n4599 = f0 & n4598;
  assign n4600 = ~a0 & n4479;
  assign n4601 = ~b0 & n4600;
  assign n4602 = ~c0 & n4601;
  assign n4603 = ~o & n4602;
  assign n4604 = f0 & n4603;
  assign n4605 = ~a0 & n4492;
  assign n4606 = ~b0 & n4605;
  assign n4607 = ~c0 & n4606;
  assign n4608 = f0 & n4607;
  assign n4609 = d0 & n4346;
  assign n4610 = ~g0 & n4609;
  assign n4611 = ~i0 & n4610;
  assign n4612 = ~e0 & n4611;
  assign n4613 = ~f0 & n4612;
  assign n4614 = v & n4613;
  assign n4615 = d0 & n4362;
  assign n4616 = ~g0 & n4615;
  assign n4617 = i0 & n4616;
  assign n4618 = ~e0 & n4617;
  assign n4619 = ~f0 & n4618;
  assign n4620 = v & n4619;
  assign n4621 = u & ~c0;
  assign n4622 = h0 & n4621;
  assign n4623 = ~g0 & n4622;
  assign n4624 = j0 & n4623;
  assign n4625 = ~i0 & n4624;
  assign n4626 = ~e0 & n4625;
  assign n4627 = ~f0 & n4626;
  assign n4628 = z & n4627;
  assign n4629 = ~g0 & n2162;
  assign n4630 = j0 & n4629;
  assign n4631 = ~i0 & n4630;
  assign n4632 = ~e0 & n4631;
  assign n4633 = ~f0 & n4632;
  assign n4634 = v & n4633;
  assign n4635 = ~n222 & n2230;
  assign n4636 = ~n217 & n4635;
  assign n4637 = ~n212 & n4636;
  assign n4638 = ~n207 & n4637;
  assign n4639 = ~n202 & n4638;
  assign n4640 = ~n197 & n4639;
  assign n4641 = ~n192 & n4640;
  assign n4642 = ~n2536 & n4641;
  assign n4643 = ~n2528 & n4642;
  assign n4644 = ~n184 & n4643;
  assign n4645 = ~n175 & n4644;
  assign n4646 = ~n2520 & n4645;
  assign n4647 = ~n2512 & n4646;
  assign n4648 = ~n139 & n4647;
  assign n4649 = ~n135 & n4648;
  assign n4650 = ~n131 & n4649;
  assign n4651 = ~n115 & n4650;
  assign n4652 = ~n108 & n4651;
  assign n4653 = ~n101 & n4652;
  assign n4654 = ~n97 & n4653;
  assign n4655 = ~n88 & n4654;
  assign n4656 = ~n84 & n4655;
  assign n4657 = ~n75 & n4656;
  assign n4658 = ~n67 & n4657;
  assign n4659 = ~n58 & n4658;
  assign n4660 = ~n50 & n4659;
  assign n4661 = ~n4634 & n4660;
  assign n4662 = ~n4628 & n4661;
  assign n4663 = ~n4620 & n4662;
  assign n4664 = ~n4614 & n4663;
  assign n4665 = ~n4608 & n4664;
  assign n4666 = ~n4604 & n4665;
  assign n4667 = ~n4599 & n4666;
  assign n4668 = ~n4594 & n4667;
  assign n4669 = ~n4588 & n4668;
  assign n4670 = ~n4581 & n4669;
  assign n4671 = ~n4574 & n4670;
  assign n4672 = ~n4572 & n4671;
  assign n4673 = ~n4569 & n4672;
  assign n4674 = ~n4560 & n4673;
  assign n4675 = ~n4551 & n4674;
  assign n4676 = ~n4548 & n4675;
  assign n4677 = ~n4544 & n4676;
  assign n4678 = ~n4541 & n4677;
  assign n4679 = ~n4537 & n4678;
  assign n4680 = ~n4533 & n4679;
  assign n4681 = ~n4528 & n4680;
  assign n4682 = ~n4524 & n4681;
  assign n4683 = ~n4519 & n4682;
  assign n4684 = ~n4511 & n4683;
  assign n4685 = ~n4502 & n4684;
  assign n4686 = ~n4497 & n4685;
  assign n4687 = ~n4491 & n4686;
  assign n4688 = ~n4485 & n4687;
  assign n4689 = ~n4478 & n4688;
  assign n4690 = ~n4471 & n4689;
  assign n4691 = ~n4468 & n4690;
  assign n4692 = ~n4460 & n4691;
  assign n4693 = ~n4451 & n4692;
  assign n4694 = ~n4445 & n4693;
  assign n4695 = ~n4438 & n4694;
  assign n4696 = ~n4431 & n4695;
  assign n4697 = ~n4423 & n4696;
  assign n4698 = ~n4415 & n4697;
  assign n4699 = ~n4411 & n4698;
  assign n4700 = ~n4402 & n4699;
  assign n4701 = ~n4392 & n4700;
  assign n4702 = ~n4386 & n4701;
  assign n4703 = ~n4379 & n4702;
  assign n4704 = ~n4370 & n4703;
  assign n4705 = ~n4361 & n4704;
  assign n4706 = ~n4354 & n4705;
  assign n4707 = ~n4344 & n4706;
  assign n4708 = ~n4338 & n4707;
  assign n4709 = ~n4335 & n4708;
  assign n4710 = ~n4328 & n4709;
  assign n4711 = ~n4321 & n4710;
  assign n4712 = ~n4317 & n4711;
  assign n4713 = ~n4308 & n4712;
  assign n4714 = ~n4301 & n4713;
  assign n4715 = ~n4297 & n4714;
  assign n4716 = ~n4289 & n4715;
  assign n4717 = ~n4280 & n4716;
  assign n4718 = ~n4275 & n4717;
  assign n4719 = ~n4265 & n4718;
  assign n4720 = ~n4257 & n4719;
  assign n4721 = ~n4249 & n4720;
  assign n4722 = ~n4240 & n4721;
  assign n4723 = ~n4235 & n4722;
  assign n4724 = ~n4226 & n4723;
  assign n4725 = ~n4217 & n4724;
  assign n4726 = ~n4207 & n4725;
  assign n4727 = ~n4201 & n4726;
  assign n4728 = ~n4192 & n4727;
  assign n4729 = ~n4182 & n4728;
  assign n4730 = ~n4174 & n4729;
  assign n4731 = ~n4164 & n4730;
  assign n4732 = ~n4153 & n4731;
  assign n4733 = ~n4144 & n4732;
  assign n4734 = ~n4136 & n4733;
  assign n4735 = ~n4126 & n4734;
  assign n4736 = ~n4115 & n4735;
  assign n4737 = ~n4104 & n4736;
  assign n4738 = ~n4092 & n4737;
  assign n4739 = ~n4084 & n4738;
  assign n4740 = ~n4075 & n4739;
  assign n4741 = ~n4070 & n4740;
  assign n4742 = ~n4061 & n4741;
  assign n4743 = ~n4050 & n4742;
  assign n4744 = ~n4038 & n4743;
  assign n4745 = ~n4026 & n4744;
  assign n4746 = ~n4013 & n4745;
  assign n4747 = ~n4004 & n4746;
  assign n4748 = ~n3994 & n4747;
  assign n4749 = ~n3988 & n4748;
  assign n4750 = ~n3979 & n4749;
  assign n4751 = ~n3969 & n4750;
  assign n4752 = ~n3961 & n4751;
  assign n4753 = ~n3951 & n4752;
  assign n4754 = ~n3940 & n4753;
  assign n4755 = ~n3931 & n4754;
  assign n4756 = ~n3921 & n4755;
  assign n4757 = ~n3910 & n4756;
  assign n4758 = ~n3899 & n4757;
  assign n4759 = ~n3887 & n4758;
  assign n4760 = ~n3874 & n4759;
  assign n4761 = ~n3860 & n4760;
  assign n4762 = ~n3846 & n4761;
  assign n4763 = ~n3832 & n4762;
  assign n4764 = ~n3823 & n4763;
  assign n4765 = ~n3813 & n4764;
  assign n4766 = ~n3804 & n4765;
  assign n4767 = ~n3794 & n4766;
  assign n4768 = ~n3784 & n4767;
  assign n4769 = ~n3773 & n4768;
  assign n4770 = ~n3766 & n4769;
  assign n4771 = ~n3758 & n4770;
  assign n4772 = ~n3749 & n4771;
  assign n4773 = ~n3739 & n4772;
  assign n4774 = ~n3730 & n4773;
  assign n4775 = ~n3720 & n4774;
  assign n4776 = ~n3708 & n4775;
  assign n4777 = ~n3695 & n4776;
  assign n4778 = ~n3684 & n4777;
  assign n4779 = ~n3672 & n4778;
  assign n4780 = ~n3662 & n4779;
  assign n4781 = ~n3651 & n4780;
  assign n4782 = ~n3640 & n4781;
  assign n4783 = ~n3628 & n4782;
  assign n4784 = ~n3619 & n4783;
  assign n4785 = ~n3609 & n4784;
  assign n4786 = ~n3600 & n4785;
  assign n4787 = ~n3590 & n4786;
  assign n4788 = ~n3580 & n4787;
  assign n4789 = ~n3569 & n4788;
  assign n4790 = ~n3562 & n4789;
  assign n4791 = ~n3554 & n4790;
  assign n4792 = ~n3546 & n4791;
  assign n4793 = ~n3537 & n4792;
  assign n4794 = ~n3529 & n4793;
  assign n4795 = ~n3520 & n4794;
  assign n4796 = ~n3511 & n4795;
  assign n4797 = ~n3501 & n4796;
  assign n4798 = ~n3495 & n4797;
  assign n4799 = ~n3488 & n4798;
  assign n4800 = ~n3484 & n4799;
  assign n4801 = ~n3479 & n4800;
  assign n4802 = ~n3475 & n4801;
  assign n4803 = ~n3470 & n4802;
  assign n4804 = ~n3465 & n4803;
  assign n4805 = ~n3459 & n4804;
  assign n4806 = ~n3454 & n4805;
  assign n4807 = ~n3448 & n4806;
  assign n4808 = ~n3436 & n4807;
  assign n4809 = ~n3423 & n4808;
  assign n4810 = ~n3410 & n4809;
  assign n4811 = ~n3396 & n4810;
  assign n4812 = ~n3387 & n4811;
  assign n4813 = ~n3377 & n4812;
  assign n4814 = ~n3368 & n4813;
  assign n4815 = ~n3358 & n4814;
  assign n4816 = ~n3346 & n4815;
  assign n4817 = ~n3333 & n4816;
  assign n4818 = ~n3322 & n4817;
  assign n4819 = ~n3310 & n4818;
  assign n4820 = ~n3300 & n4819;
  assign n4821 = ~n3289 & n4820;
  assign n4822 = ~n3278 & n4821;
  assign n4823 = ~n3266 & n4822;
  assign n4824 = ~n3254 & n4823;
  assign n4825 = ~n3241 & n4824;
  assign n4826 = ~n3228 & n4825;
  assign n4827 = ~n3214 & n4826;
  assign n4828 = ~n3206 & n4827;
  assign n4829 = ~n3196 & n4828;
  assign n4830 = ~n3187 & n4829;
  assign n4831 = ~n3176 & n4830;
  assign n4832 = ~n3168 & n4831;
  assign n4833 = ~n3158 & n4832;
  assign n4834 = ~n3149 & n4833;
  assign n4835 = ~n3138 & n4834;
  assign n4836 = ~n3125 & n4835;
  assign n4837 = ~n3111 & n4836;
  assign n4838 = ~n3097 & n4837;
  assign n4839 = ~n3082 & n4838;
  assign n4840 = ~n3070 & n4839;
  assign n4841 = ~n3057 & n4840;
  assign n4842 = ~n3044 & n4841;
  assign n4843 = ~n3030 & n4842;
  assign n4844 = ~n3028 & n4843;
  assign n4845 = ~n3025 & n4844;
  assign n4846 = ~n3022 & n4845;
  assign n4847 = ~n3018 & n4846;
  assign n4848 = ~n3015 & n4847;
  assign n4849 = ~n3011 & n4848;
  assign n4850 = ~n3008 & n4849;
  assign n4851 = ~n3004 & n4850;
  assign n4852 = ~n3000 & n4851;
  assign n4853 = ~n2995 & n4852;
  assign n4854 = ~n2991 & n4853;
  assign n4855 = ~n2986 & n4854;
  assign n4856 = ~n2973 & n4855;
  assign n4857 = ~n2959 & n4856;
  assign n4858 = ~n2945 & n4857;
  assign n4859 = ~n2930 & n4858;
  assign n4860 = ~n2918 & n4859;
  assign n4861 = ~n2905 & n4860;
  assign n4862 = ~n2892 & n4861;
  assign n4863 = ~n2878 & n4862;
  assign n4864 = ~n2865 & n4863;
  assign n4865 = ~n2851 & n4864;
  assign n4866 = ~n2837 & n4865;
  assign n4867 = ~n2822 & n4866;
  assign n4868 = ~n2814 & n4867;
  assign n4869 = ~n2804 & n4868;
  assign n4870 = ~n2795 & n4869;
  assign n4871 = ~n2784 & n4870;
  assign n4872 = ~n2776 & n4871;
  assign n4873 = ~n2766 & n4872;
  assign n4874 = ~n2757 & n4873;
  assign n4875 = ~n2746 & n4874;
  assign n4876 = ~n2737 & n4875;
  assign n4877 = ~n2726 & n4876;
  assign n4878 = ~n2716 & n4877;
  assign n4879 = ~n2704 & n4878;
  assign n4880 = ~n2698 & n4879;
  assign n4881 = ~n2690 & n4880;
  assign n4882 = ~n2683 & n4881;
  assign n4883 = ~n2674 & n4882;
  assign n4884 = ~n2673 & n4883;
  assign n4885 = ~n2671 & n4884;
  assign n4886 = ~n2669 & n4885;
  assign n4887 = ~n2666 & n4886;
  assign n4888 = ~n2652 & n4887;
  assign n4889 = ~n2636 & n4888;
  assign n4890 = ~n2621 & n4889;
  assign n4891 = ~n2604 & n4890;
  assign n4892 = ~n2589 & n4891;
  assign n4893 = ~n2572 & n4892;
  assign o0 = n2556 | ~n4893;
  assign n4895 = ~c & j;
  assign n4896 = ~n & n4895;
  assign n4897 = ~y & n4896;
  assign n4898 = ~c0 & n4897;
  assign n4899 = ~j0 & n4898;
  assign n4900 = m0 & n4899;
  assign n4901 = ~h0 & n4900;
  assign n4902 = ~e & n4901;
  assign n4903 = ~f & n4902;
  assign n4904 = ~g & n4903;
  assign n4905 = ~i & n4904;
  assign n4906 = t & n4905;
  assign n4907 = ~d0 & n4906;
  assign n4908 = i0 & n4907;
  assign n4909 = ~d & n4908;
  assign n4910 = ~m & n4909;
  assign n4911 = ~z & n4897;
  assign n4912 = ~c0 & n4911;
  assign n4913 = ~j0 & n4912;
  assign n4914 = m0 & n4913;
  assign n4915 = ~e & n4914;
  assign n4916 = ~f & n4915;
  assign n4917 = ~g & n4916;
  assign n4918 = ~i & n4917;
  assign n4919 = t & n4918;
  assign n4920 = ~d0 & n4919;
  assign n4921 = i0 & n4920;
  assign n4922 = ~d & n4921;
  assign n4923 = ~m & n4922;
  assign n4924 = ~g0 & n4898;
  assign n4925 = ~j0 & n4924;
  assign n4926 = m0 & n4925;
  assign n4927 = ~h0 & n4926;
  assign n4928 = ~e & n4927;
  assign n4929 = ~f & n4928;
  assign n4930 = ~g & n4929;
  assign n4931 = t & n4930;
  assign n4932 = ~d0 & n4931;
  assign n4933 = i0 & n4932;
  assign n4934 = ~d & n4933;
  assign n4935 = ~m & n4934;
  assign n4936 = ~g0 & n4912;
  assign n4937 = ~j0 & n4936;
  assign n4938 = m0 & n4937;
  assign n4939 = ~e & n4938;
  assign n4940 = ~f & n4939;
  assign n4941 = ~g & n4940;
  assign n4942 = t & n4941;
  assign n4943 = ~d0 & n4942;
  assign n4944 = i0 & n4943;
  assign n4945 = ~d & n4944;
  assign n4946 = ~m & n4945;
  assign n4947 = l & n4895;
  assign n4948 = ~n & n4947;
  assign n4949 = ~y & n4948;
  assign n4950 = ~c0 & n4949;
  assign n4951 = ~j0 & n4950;
  assign n4952 = m0 & n4951;
  assign n4953 = ~h0 & n4952;
  assign n4954 = ~e & n4953;
  assign n4955 = ~f & n4954;
  assign n4956 = ~g & n4955;
  assign n4957 = ~i & n4956;
  assign n4958 = ~d0 & n4957;
  assign n4959 = i0 & n4958;
  assign n4960 = ~d & n4959;
  assign n4961 = ~m & n4960;
  assign n4962 = ~z & n4949;
  assign n4963 = ~c0 & n4962;
  assign n4964 = ~j0 & n4963;
  assign n4965 = m0 & n4964;
  assign n4966 = ~e & n4965;
  assign n4967 = ~f & n4966;
  assign n4968 = ~g & n4967;
  assign n4969 = ~i & n4968;
  assign n4970 = ~d0 & n4969;
  assign n4971 = i0 & n4970;
  assign n4972 = ~d & n4971;
  assign n4973 = ~m & n4972;
  assign n4974 = ~g0 & n4950;
  assign n4975 = ~j0 & n4974;
  assign n4976 = m0 & n4975;
  assign n4977 = ~h0 & n4976;
  assign n4978 = ~e & n4977;
  assign n4979 = ~f & n4978;
  assign n4980 = ~g & n4979;
  assign n4981 = ~d0 & n4980;
  assign n4982 = i0 & n4981;
  assign n4983 = ~d & n4982;
  assign n4984 = ~m & n4983;
  assign n4985 = ~g0 & n4963;
  assign n4986 = ~j0 & n4985;
  assign n4987 = m0 & n4986;
  assign n4988 = ~e & n4987;
  assign n4989 = ~f & n4988;
  assign n4990 = ~g & n4989;
  assign n4991 = ~d0 & n4990;
  assign n4992 = i0 & n4991;
  assign n4993 = ~d & n4992;
  assign n4994 = ~m & n4993;
  assign n4995 = ~a0 & n4897;
  assign n4996 = ~c0 & n4995;
  assign n4997 = ~j0 & n4996;
  assign n4998 = m0 & n4997;
  assign n4999 = ~h0 & n4998;
  assign n5000 = ~e & n4999;
  assign n5001 = ~f & n5000;
  assign n5002 = ~g & n5001;
  assign n5003 = ~i & n5002;
  assign n5004 = t & n5003;
  assign n5005 = ~d0 & n5004;
  assign n5006 = ~d & n5005;
  assign n5007 = ~m & n5006;
  assign n5008 = ~a0 & n4911;
  assign n5009 = ~c0 & n5008;
  assign n5010 = ~j0 & n5009;
  assign n5011 = m0 & n5010;
  assign n5012 = ~e & n5011;
  assign n5013 = ~f & n5012;
  assign n5014 = ~g & n5013;
  assign n5015 = ~i & n5014;
  assign n5016 = t & n5015;
  assign n5017 = ~d0 & n5016;
  assign n5018 = ~d & n5017;
  assign n5019 = ~m & n5018;
  assign n5020 = ~g0 & n4996;
  assign n5021 = ~j0 & n5020;
  assign n5022 = m0 & n5021;
  assign n5023 = ~h0 & n5022;
  assign n5024 = ~e & n5023;
  assign n5025 = ~f & n5024;
  assign n5026 = ~g & n5025;
  assign n5027 = t & n5026;
  assign n5028 = ~d0 & n5027;
  assign n5029 = ~d & n5028;
  assign n5030 = ~m & n5029;
  assign n5031 = ~g0 & n5009;
  assign n5032 = ~j0 & n5031;
  assign n5033 = m0 & n5032;
  assign n5034 = ~e & n5033;
  assign n5035 = ~f & n5034;
  assign n5036 = ~g & n5035;
  assign n5037 = t & n5036;
  assign n5038 = ~d0 & n5037;
  assign n5039 = ~d & n5038;
  assign n5040 = ~m & n5039;
  assign n5041 = ~a0 & n4949;
  assign n5042 = ~c0 & n5041;
  assign n5043 = ~j0 & n5042;
  assign n5044 = m0 & n5043;
  assign n5045 = ~h0 & n5044;
  assign n5046 = ~e & n5045;
  assign n5047 = ~f & n5046;
  assign n5048 = ~g & n5047;
  assign n5049 = ~i & n5048;
  assign n5050 = ~d0 & n5049;
  assign n5051 = ~d & n5050;
  assign n5052 = ~m & n5051;
  assign n5053 = ~a0 & n4962;
  assign n5054 = ~c0 & n5053;
  assign n5055 = ~j0 & n5054;
  assign n5056 = m0 & n5055;
  assign n5057 = ~e & n5056;
  assign n5058 = ~f & n5057;
  assign n5059 = ~g & n5058;
  assign n5060 = ~i & n5059;
  assign n5061 = ~d0 & n5060;
  assign n5062 = ~d & n5061;
  assign n5063 = ~m & n5062;
  assign n5064 = ~g0 & n5042;
  assign n5065 = ~j0 & n5064;
  assign n5066 = m0 & n5065;
  assign n5067 = ~h0 & n5066;
  assign n5068 = ~e & n5067;
  assign n5069 = ~f & n5068;
  assign n5070 = ~g & n5069;
  assign n5071 = ~d0 & n5070;
  assign n5072 = ~d & n5071;
  assign n5073 = ~m & n5072;
  assign n5074 = ~g0 & n5054;
  assign n5075 = ~j0 & n5074;
  assign n5076 = m0 & n5075;
  assign n5077 = ~e & n5076;
  assign n5078 = ~f & n5077;
  assign n5079 = ~g & n5078;
  assign n5080 = ~d0 & n5079;
  assign n5081 = ~d & n5080;
  assign n5082 = ~m & n5081;
  assign n5083 = ~w & n4896;
  assign n5084 = ~y & n5083;
  assign n5085 = ~a0 & n5084;
  assign n5086 = ~c0 & n5085;
  assign n5087 = ~j0 & n5086;
  assign n5088 = m0 & n5087;
  assign n5089 = ~h0 & n5088;
  assign n5090 = ~e & n5089;
  assign n5091 = ~f & n5090;
  assign n5092 = ~g & n5091;
  assign n5093 = ~i & n5092;
  assign n5094 = t & n5093;
  assign n5095 = ~d & n5094;
  assign n5096 = ~m & n5095;
  assign n5097 = ~z & n5084;
  assign n5098 = ~a0 & n5097;
  assign n5099 = ~c0 & n5098;
  assign n5100 = ~j0 & n5099;
  assign n5101 = m0 & n5100;
  assign n5102 = ~e & n5101;
  assign n5103 = ~f & n5102;
  assign n5104 = ~g & n5103;
  assign n5105 = ~i & n5104;
  assign n5106 = t & n5105;
  assign n5107 = ~d & n5106;
  assign n5108 = ~m & n5107;
  assign n5109 = ~g0 & n5086;
  assign n5110 = ~j0 & n5109;
  assign n5111 = m0 & n5110;
  assign n5112 = ~h0 & n5111;
  assign n5113 = ~e & n5112;
  assign n5114 = ~f & n5113;
  assign n5115 = ~g & n5114;
  assign n5116 = t & n5115;
  assign n5117 = ~d & n5116;
  assign n5118 = ~m & n5117;
  assign n5119 = ~g0 & n5099;
  assign n5120 = ~j0 & n5119;
  assign n5121 = m0 & n5120;
  assign n5122 = ~e & n5121;
  assign n5123 = ~f & n5122;
  assign n5124 = ~g & n5123;
  assign n5125 = t & n5124;
  assign n5126 = ~d & n5125;
  assign n5127 = ~m & n5126;
  assign n5128 = ~w & n4948;
  assign n5129 = ~y & n5128;
  assign n5130 = ~a0 & n5129;
  assign n5131 = ~c0 & n5130;
  assign n5132 = ~j0 & n5131;
  assign n5133 = m0 & n5132;
  assign n5134 = ~h0 & n5133;
  assign n5135 = ~e & n5134;
  assign n5136 = ~f & n5135;
  assign n5137 = ~g & n5136;
  assign n5138 = ~i & n5137;
  assign n5139 = ~d & n5138;
  assign n5140 = ~m & n5139;
  assign n5141 = ~z & n5129;
  assign n5142 = ~a0 & n5141;
  assign n5143 = ~c0 & n5142;
  assign n5144 = ~j0 & n5143;
  assign n5145 = m0 & n5144;
  assign n5146 = ~e & n5145;
  assign n5147 = ~f & n5146;
  assign n5148 = ~g & n5147;
  assign n5149 = ~i & n5148;
  assign n5150 = ~d & n5149;
  assign n5151 = ~m & n5150;
  assign n5152 = ~g0 & n5131;
  assign n5153 = ~j0 & n5152;
  assign n5154 = m0 & n5153;
  assign n5155 = ~h0 & n5154;
  assign n5156 = ~e & n5155;
  assign n5157 = ~f & n5156;
  assign n5158 = ~g & n5157;
  assign n5159 = ~d & n5158;
  assign n5160 = ~m & n5159;
  assign n5161 = ~g0 & n5143;
  assign n5162 = ~j0 & n5161;
  assign n5163 = m0 & n5162;
  assign n5164 = ~e & n5163;
  assign n5165 = ~f & n5164;
  assign n5166 = ~g & n5165;
  assign n5167 = ~d & n5166;
  assign n5168 = ~m & n5167;
  assign n5169 = s & n4896;
  assign n5170 = ~y & n5169;
  assign n5171 = ~c0 & n5170;
  assign n5172 = ~j0 & n5171;
  assign n5173 = m0 & n5172;
  assign n5174 = ~h0 & n5173;
  assign n5175 = ~e & n5174;
  assign n5176 = ~f & n5175;
  assign n5177 = ~g & n5176;
  assign n5178 = ~i & n5177;
  assign n5179 = t & n5178;
  assign n5180 = ~d0 & n5179;
  assign n5181 = i0 & n5180;
  assign n5182 = ~m & n5181;
  assign n5183 = ~z & n5170;
  assign n5184 = ~c0 & n5183;
  assign n5185 = ~j0 & n5184;
  assign n5186 = m0 & n5185;
  assign n5187 = ~e & n5186;
  assign n5188 = ~f & n5187;
  assign n5189 = ~g & n5188;
  assign n5190 = ~i & n5189;
  assign n5191 = t & n5190;
  assign n5192 = ~d0 & n5191;
  assign n5193 = i0 & n5192;
  assign n5194 = ~m & n5193;
  assign n5195 = ~g0 & n5171;
  assign n5196 = ~j0 & n5195;
  assign n5197 = m0 & n5196;
  assign n5198 = ~h0 & n5197;
  assign n5199 = ~e & n5198;
  assign n5200 = ~f & n5199;
  assign n5201 = ~g & n5200;
  assign n5202 = t & n5201;
  assign n5203 = ~d0 & n5202;
  assign n5204 = i0 & n5203;
  assign n5205 = ~m & n5204;
  assign n5206 = ~g0 & n5184;
  assign n5207 = ~j0 & n5206;
  assign n5208 = m0 & n5207;
  assign n5209 = ~e & n5208;
  assign n5210 = ~f & n5209;
  assign n5211 = ~g & n5210;
  assign n5212 = t & n5211;
  assign n5213 = ~d0 & n5212;
  assign n5214 = i0 & n5213;
  assign n5215 = ~m & n5214;
  assign n5216 = s & n4948;
  assign n5217 = ~y & n5216;
  assign n5218 = ~c0 & n5217;
  assign n5219 = ~j0 & n5218;
  assign n5220 = m0 & n5219;
  assign n5221 = ~h0 & n5220;
  assign n5222 = ~e & n5221;
  assign n5223 = ~f & n5222;
  assign n5224 = ~g & n5223;
  assign n5225 = ~i & n5224;
  assign n5226 = ~d0 & n5225;
  assign n5227 = i0 & n5226;
  assign n5228 = ~m & n5227;
  assign n5229 = ~z & n5217;
  assign n5230 = ~c0 & n5229;
  assign n5231 = ~j0 & n5230;
  assign n5232 = m0 & n5231;
  assign n5233 = ~e & n5232;
  assign n5234 = ~f & n5233;
  assign n5235 = ~g & n5234;
  assign n5236 = ~i & n5235;
  assign n5237 = ~d0 & n5236;
  assign n5238 = i0 & n5237;
  assign n5239 = ~m & n5238;
  assign n5240 = ~g0 & n5218;
  assign n5241 = ~j0 & n5240;
  assign n5242 = m0 & n5241;
  assign n5243 = ~h0 & n5242;
  assign n5244 = ~e & n5243;
  assign n5245 = ~f & n5244;
  assign n5246 = ~g & n5245;
  assign n5247 = ~d0 & n5246;
  assign n5248 = i0 & n5247;
  assign n5249 = ~m & n5248;
  assign n5250 = ~g0 & n5230;
  assign n5251 = ~j0 & n5250;
  assign n5252 = m0 & n5251;
  assign n5253 = ~e & n5252;
  assign n5254 = ~f & n5253;
  assign n5255 = ~g & n5254;
  assign n5256 = ~d0 & n5255;
  assign n5257 = i0 & n5256;
  assign n5258 = ~m & n5257;
  assign n5259 = ~a0 & n5170;
  assign n5260 = ~c0 & n5259;
  assign n5261 = ~j0 & n5260;
  assign n5262 = m0 & n5261;
  assign n5263 = ~h0 & n5262;
  assign n5264 = ~e & n5263;
  assign n5265 = ~f & n5264;
  assign n5266 = ~g & n5265;
  assign n5267 = ~i & n5266;
  assign n5268 = t & n5267;
  assign n5269 = ~d0 & n5268;
  assign n5270 = ~m & n5269;
  assign n5271 = ~a0 & n5183;
  assign n5272 = ~c0 & n5271;
  assign n5273 = ~j0 & n5272;
  assign n5274 = m0 & n5273;
  assign n5275 = ~e & n5274;
  assign n5276 = ~f & n5275;
  assign n5277 = ~g & n5276;
  assign n5278 = ~i & n5277;
  assign n5279 = t & n5278;
  assign n5280 = ~d0 & n5279;
  assign n5281 = ~m & n5280;
  assign n5282 = ~g0 & n5260;
  assign n5283 = ~j0 & n5282;
  assign n5284 = m0 & n5283;
  assign n5285 = ~h0 & n5284;
  assign n5286 = ~e & n5285;
  assign n5287 = ~f & n5286;
  assign n5288 = ~g & n5287;
  assign n5289 = t & n5288;
  assign n5290 = ~d0 & n5289;
  assign n5291 = ~m & n5290;
  assign n5292 = ~g0 & n5272;
  assign n5293 = ~j0 & n5292;
  assign n5294 = m0 & n5293;
  assign n5295 = ~e & n5294;
  assign n5296 = ~f & n5295;
  assign n5297 = ~g & n5296;
  assign n5298 = t & n5297;
  assign n5299 = ~d0 & n5298;
  assign n5300 = ~m & n5299;
  assign n5301 = ~a0 & n5217;
  assign n5302 = ~c0 & n5301;
  assign n5303 = ~j0 & n5302;
  assign n5304 = m0 & n5303;
  assign n5305 = ~h0 & n5304;
  assign n5306 = ~e & n5305;
  assign n5307 = ~f & n5306;
  assign n5308 = ~g & n5307;
  assign n5309 = ~i & n5308;
  assign n5310 = ~d0 & n5309;
  assign n5311 = ~m & n5310;
  assign n5312 = ~a0 & n5229;
  assign n5313 = ~c0 & n5312;
  assign n5314 = ~j0 & n5313;
  assign n5315 = m0 & n5314;
  assign n5316 = ~e & n5315;
  assign n5317 = ~f & n5316;
  assign n5318 = ~g & n5317;
  assign n5319 = ~i & n5318;
  assign n5320 = ~d0 & n5319;
  assign n5321 = ~m & n5320;
  assign n5322 = ~g0 & n5302;
  assign n5323 = ~j0 & n5322;
  assign n5324 = m0 & n5323;
  assign n5325 = ~h0 & n5324;
  assign n5326 = ~e & n5325;
  assign n5327 = ~f & n5326;
  assign n5328 = ~g & n5327;
  assign n5329 = ~d0 & n5328;
  assign n5330 = ~m & n5329;
  assign n5331 = ~g0 & n5313;
  assign n5332 = ~j0 & n5331;
  assign n5333 = m0 & n5332;
  assign n5334 = ~e & n5333;
  assign n5335 = ~f & n5334;
  assign n5336 = ~g & n5335;
  assign n5337 = ~d0 & n5336;
  assign n5338 = ~m & n5337;
  assign n5339 = ~w & n5169;
  assign n5340 = ~y & n5339;
  assign n5341 = ~a0 & n5340;
  assign n5342 = ~c0 & n5341;
  assign n5343 = ~j0 & n5342;
  assign n5344 = m0 & n5343;
  assign n5345 = ~h0 & n5344;
  assign n5346 = ~e & n5345;
  assign n5347 = ~f & n5346;
  assign n5348 = ~g & n5347;
  assign n5349 = ~i & n5348;
  assign n5350 = t & n5349;
  assign n5351 = ~m & n5350;
  assign n5352 = ~z & n5340;
  assign n5353 = ~a0 & n5352;
  assign n5354 = ~c0 & n5353;
  assign n5355 = ~j0 & n5354;
  assign n5356 = m0 & n5355;
  assign n5357 = ~e & n5356;
  assign n5358 = ~f & n5357;
  assign n5359 = ~g & n5358;
  assign n5360 = ~i & n5359;
  assign n5361 = t & n5360;
  assign n5362 = ~m & n5361;
  assign n5363 = ~g0 & n5342;
  assign n5364 = ~j0 & n5363;
  assign n5365 = m0 & n5364;
  assign n5366 = ~h0 & n5365;
  assign n5367 = ~e & n5366;
  assign n5368 = ~f & n5367;
  assign n5369 = ~g & n5368;
  assign n5370 = t & n5369;
  assign n5371 = ~m & n5370;
  assign n5372 = ~g0 & n5354;
  assign n5373 = ~j0 & n5372;
  assign n5374 = m0 & n5373;
  assign n5375 = ~e & n5374;
  assign n5376 = ~f & n5375;
  assign n5377 = ~g & n5376;
  assign n5378 = t & n5377;
  assign n5379 = ~m & n5378;
  assign n5380 = ~w & n5216;
  assign n5381 = ~y & n5380;
  assign n5382 = ~a0 & n5381;
  assign n5383 = ~c0 & n5382;
  assign n5384 = ~j0 & n5383;
  assign n5385 = m0 & n5384;
  assign n5386 = ~h0 & n5385;
  assign n5387 = ~e & n5386;
  assign n5388 = ~f & n5387;
  assign n5389 = ~g & n5388;
  assign n5390 = ~i & n5389;
  assign n5391 = ~m & n5390;
  assign n5392 = ~z & n5381;
  assign n5393 = ~a0 & n5392;
  assign n5394 = ~c0 & n5393;
  assign n5395 = ~j0 & n5394;
  assign n5396 = m0 & n5395;
  assign n5397 = ~e & n5396;
  assign n5398 = ~f & n5397;
  assign n5399 = ~g & n5398;
  assign n5400 = ~i & n5399;
  assign n5401 = ~m & n5400;
  assign n5402 = ~g0 & n5383;
  assign n5403 = ~j0 & n5402;
  assign n5404 = m0 & n5403;
  assign n5405 = ~h0 & n5404;
  assign n5406 = ~e & n5405;
  assign n5407 = ~f & n5406;
  assign n5408 = ~g & n5407;
  assign n5409 = ~m & n5408;
  assign n5410 = ~g0 & n5394;
  assign n5411 = ~j0 & n5410;
  assign n5412 = m0 & n5411;
  assign n5413 = ~e & n5412;
  assign n5414 = ~f & n5413;
  assign n5415 = ~g & n5414;
  assign n5416 = ~m & n5415;
  assign n5417 = ~b & n4908;
  assign n5418 = ~d & n5417;
  assign n5419 = ~b & n4921;
  assign n5420 = ~d & n5419;
  assign n5421 = ~b & n4933;
  assign n5422 = ~d & n5421;
  assign n5423 = ~b & n4944;
  assign n5424 = ~d & n5423;
  assign n5425 = ~b & n4959;
  assign n5426 = ~d & n5425;
  assign n5427 = ~b & n4971;
  assign n5428 = ~d & n5427;
  assign n5429 = ~b & n4982;
  assign n5430 = ~d & n5429;
  assign n5431 = ~b & n4992;
  assign n5432 = ~d & n5431;
  assign n5433 = ~b & n5005;
  assign n5434 = ~d & n5433;
  assign n5435 = ~b & n5017;
  assign n5436 = ~d & n5435;
  assign n5437 = ~b & n5028;
  assign n5438 = ~d & n5437;
  assign n5439 = ~b & n5038;
  assign n5440 = ~d & n5439;
  assign n5441 = ~b & n5050;
  assign n5442 = ~d & n5441;
  assign n5443 = ~b & n5061;
  assign n5444 = ~d & n5443;
  assign n5445 = ~b & n5071;
  assign n5446 = ~d & n5445;
  assign n5447 = ~b & n5080;
  assign n5448 = ~d & n5447;
  assign n5449 = ~b & n5094;
  assign n5450 = ~d & n5449;
  assign n5451 = ~b & n5106;
  assign n5452 = ~d & n5451;
  assign n5453 = ~b & n5116;
  assign n5454 = ~d & n5453;
  assign n5455 = ~b & n5125;
  assign n5456 = ~d & n5455;
  assign n5457 = ~b & n5138;
  assign n5458 = ~d & n5457;
  assign n5459 = ~b & n5149;
  assign n5460 = ~d & n5459;
  assign n5461 = ~b & n5158;
  assign n5462 = ~d & n5461;
  assign n5463 = ~b & n5166;
  assign n5464 = ~d & n5463;
  assign n5465 = ~b & n5181;
  assign n5466 = ~b & n5193;
  assign n5467 = ~b & n5204;
  assign n5468 = ~b & n5214;
  assign n5469 = ~b & n5227;
  assign n5470 = ~b & n5238;
  assign n5471 = ~b & n5248;
  assign n5472 = ~b & n5257;
  assign n5473 = ~b & n5269;
  assign n5474 = ~b & n5280;
  assign n5475 = ~b & n5290;
  assign n5476 = ~b & n5299;
  assign n5477 = ~b & n5310;
  assign n5478 = ~b & n5320;
  assign n5479 = ~b & n5329;
  assign n5480 = ~b & n5337;
  assign n5481 = ~b & n5350;
  assign n5482 = ~b & n5361;
  assign n5483 = ~b & n5370;
  assign n5484 = ~b & n5378;
  assign n5485 = ~b & n5390;
  assign n5486 = ~b & n5400;
  assign n5487 = ~b & n5408;
  assign n5488 = ~b & n5415;
  assign n5489 = ~c & ~j;
  assign n5490 = ~s & n5489;
  assign n5491 = ~y & n5490;
  assign n5492 = ~c0 & n5491;
  assign n5493 = ~j0 & n5492;
  assign n5494 = m0 & n5493;
  assign n5495 = ~f0 & n5494;
  assign n5496 = ~h0 & n5495;
  assign n5497 = ~e & n5496;
  assign n5498 = ~f & n5497;
  assign n5499 = ~g & n5498;
  assign n5500 = ~i & n5499;
  assign n5501 = ~d0 & n5500;
  assign n5502 = i0 & n5501;
  assign n5503 = d & n5502;
  assign n5504 = ~z & n5491;
  assign n5505 = ~c0 & n5504;
  assign n5506 = ~j0 & n5505;
  assign n5507 = m0 & n5506;
  assign n5508 = ~f0 & n5507;
  assign n5509 = ~e & n5508;
  assign n5510 = ~f & n5509;
  assign n5511 = ~g & n5510;
  assign n5512 = ~i & n5511;
  assign n5513 = ~d0 & n5512;
  assign n5514 = i0 & n5513;
  assign n5515 = d & n5514;
  assign n5516 = ~g0 & n5492;
  assign n5517 = ~j0 & n5516;
  assign n5518 = m0 & n5517;
  assign n5519 = ~f0 & n5518;
  assign n5520 = ~h0 & n5519;
  assign n5521 = ~e & n5520;
  assign n5522 = ~f & n5521;
  assign n5523 = ~g & n5522;
  assign n5524 = ~d0 & n5523;
  assign n5525 = i0 & n5524;
  assign n5526 = d & n5525;
  assign n5527 = ~g0 & n5505;
  assign n5528 = ~j0 & n5527;
  assign n5529 = m0 & n5528;
  assign n5530 = ~f0 & n5529;
  assign n5531 = ~e & n5530;
  assign n5532 = ~f & n5531;
  assign n5533 = ~g & n5532;
  assign n5534 = ~d0 & n5533;
  assign n5535 = i0 & n5534;
  assign n5536 = d & n5535;
  assign n5537 = ~a0 & n5491;
  assign n5538 = ~c0 & n5537;
  assign n5539 = ~j0 & n5538;
  assign n5540 = m0 & n5539;
  assign n5541 = ~f0 & n5540;
  assign n5542 = ~h0 & n5541;
  assign n5543 = ~e & n5542;
  assign n5544 = ~f & n5543;
  assign n5545 = ~g & n5544;
  assign n5546 = ~i & n5545;
  assign n5547 = ~d0 & n5546;
  assign n5548 = d & n5547;
  assign n5549 = ~a0 & n5504;
  assign n5550 = ~c0 & n5549;
  assign n5551 = ~j0 & n5550;
  assign n5552 = m0 & n5551;
  assign n5553 = ~f0 & n5552;
  assign n5554 = ~e & n5553;
  assign n5555 = ~f & n5554;
  assign n5556 = ~g & n5555;
  assign n5557 = ~i & n5556;
  assign n5558 = ~d0 & n5557;
  assign n5559 = d & n5558;
  assign n5560 = ~g0 & n5538;
  assign n5561 = ~j0 & n5560;
  assign n5562 = m0 & n5561;
  assign n5563 = ~f0 & n5562;
  assign n5564 = ~h0 & n5563;
  assign n5565 = ~e & n5564;
  assign n5566 = ~f & n5565;
  assign n5567 = ~g & n5566;
  assign n5568 = ~d0 & n5567;
  assign n5569 = d & n5568;
  assign n5570 = ~g0 & n5550;
  assign n5571 = ~j0 & n5570;
  assign n5572 = m0 & n5571;
  assign n5573 = ~f0 & n5572;
  assign n5574 = ~e & n5573;
  assign n5575 = ~f & n5574;
  assign n5576 = ~g & n5575;
  assign n5577 = ~d0 & n5576;
  assign n5578 = d & n5577;
  assign n5579 = ~w & n5490;
  assign n5580 = ~y & n5579;
  assign n5581 = ~a0 & n5580;
  assign n5582 = ~c0 & n5581;
  assign n5583 = ~j0 & n5582;
  assign n5584 = m0 & n5583;
  assign n5585 = ~f0 & n5584;
  assign n5586 = ~h0 & n5585;
  assign n5587 = ~e & n5586;
  assign n5588 = ~f & n5587;
  assign n5589 = ~g & n5588;
  assign n5590 = ~i & n5589;
  assign n5591 = d & n5590;
  assign n5592 = ~z & n5580;
  assign n5593 = ~a0 & n5592;
  assign n5594 = ~c0 & n5593;
  assign n5595 = ~j0 & n5594;
  assign n5596 = m0 & n5595;
  assign n5597 = ~f0 & n5596;
  assign n5598 = ~e & n5597;
  assign n5599 = ~f & n5598;
  assign n5600 = ~g & n5599;
  assign n5601 = ~i & n5600;
  assign n5602 = d & n5601;
  assign n5603 = ~g0 & n5582;
  assign n5604 = ~j0 & n5603;
  assign n5605 = m0 & n5604;
  assign n5606 = ~f0 & n5605;
  assign n5607 = ~h0 & n5606;
  assign n5608 = ~e & n5607;
  assign n5609 = ~f & n5608;
  assign n5610 = ~g & n5609;
  assign n5611 = d & n5610;
  assign n5612 = ~g0 & n5594;
  assign n5613 = ~j0 & n5612;
  assign n5614 = m0 & n5613;
  assign n5615 = ~f0 & n5614;
  assign n5616 = ~e & n5615;
  assign n5617 = ~f & n5616;
  assign n5618 = ~g & n5617;
  assign n5619 = d & n5618;
  assign n5620 = ~l & n5489;
  assign n5621 = ~y & n5620;
  assign n5622 = ~c0 & n5621;
  assign n5623 = ~j0 & n5622;
  assign n5624 = m0 & n5623;
  assign n5625 = ~f0 & n5624;
  assign n5626 = ~h0 & n5625;
  assign n5627 = ~e & n5626;
  assign n5628 = ~f & n5627;
  assign n5629 = ~g & n5628;
  assign n5630 = ~i & n5629;
  assign n5631 = ~t & n5630;
  assign n5632 = ~d0 & n5631;
  assign n5633 = i0 & n5632;
  assign n5634 = ~z & n5621;
  assign n5635 = ~c0 & n5634;
  assign n5636 = ~j0 & n5635;
  assign n5637 = m0 & n5636;
  assign n5638 = ~f0 & n5637;
  assign n5639 = ~e & n5638;
  assign n5640 = ~f & n5639;
  assign n5641 = ~g & n5640;
  assign n5642 = ~i & n5641;
  assign n5643 = ~t & n5642;
  assign n5644 = ~d0 & n5643;
  assign n5645 = i0 & n5644;
  assign n5646 = ~g0 & n5622;
  assign n5647 = ~j0 & n5646;
  assign n5648 = m0 & n5647;
  assign n5649 = ~f0 & n5648;
  assign n5650 = ~h0 & n5649;
  assign n5651 = ~e & n5650;
  assign n5652 = ~f & n5651;
  assign n5653 = ~g & n5652;
  assign n5654 = ~t & n5653;
  assign n5655 = ~d0 & n5654;
  assign n5656 = i0 & n5655;
  assign n5657 = ~g0 & n5635;
  assign n5658 = ~j0 & n5657;
  assign n5659 = m0 & n5658;
  assign n5660 = ~f0 & n5659;
  assign n5661 = ~e & n5660;
  assign n5662 = ~f & n5661;
  assign n5663 = ~g & n5662;
  assign n5664 = ~t & n5663;
  assign n5665 = ~d0 & n5664;
  assign n5666 = i0 & n5665;
  assign n5667 = ~a0 & n5621;
  assign n5668 = ~c0 & n5667;
  assign n5669 = ~j0 & n5668;
  assign n5670 = m0 & n5669;
  assign n5671 = ~f0 & n5670;
  assign n5672 = ~h0 & n5671;
  assign n5673 = ~e & n5672;
  assign n5674 = ~f & n5673;
  assign n5675 = ~g & n5674;
  assign n5676 = ~i & n5675;
  assign n5677 = ~t & n5676;
  assign n5678 = ~d0 & n5677;
  assign n5679 = ~a0 & n5634;
  assign n5680 = ~c0 & n5679;
  assign n5681 = ~j0 & n5680;
  assign n5682 = m0 & n5681;
  assign n5683 = ~f0 & n5682;
  assign n5684 = ~e & n5683;
  assign n5685 = ~f & n5684;
  assign n5686 = ~g & n5685;
  assign n5687 = ~i & n5686;
  assign n5688 = ~t & n5687;
  assign n5689 = ~d0 & n5688;
  assign n5690 = ~g0 & n5668;
  assign n5691 = ~j0 & n5690;
  assign n5692 = m0 & n5691;
  assign n5693 = ~f0 & n5692;
  assign n5694 = ~h0 & n5693;
  assign n5695 = ~e & n5694;
  assign n5696 = ~f & n5695;
  assign n5697 = ~g & n5696;
  assign n5698 = ~t & n5697;
  assign n5699 = ~d0 & n5698;
  assign n5700 = ~g0 & n5680;
  assign n5701 = ~j0 & n5700;
  assign n5702 = m0 & n5701;
  assign n5703 = ~f0 & n5702;
  assign n5704 = ~e & n5703;
  assign n5705 = ~f & n5704;
  assign n5706 = ~g & n5705;
  assign n5707 = ~t & n5706;
  assign n5708 = ~d0 & n5707;
  assign n5709 = ~w & n5620;
  assign n5710 = ~y & n5709;
  assign n5711 = ~a0 & n5710;
  assign n5712 = ~c0 & n5711;
  assign n5713 = ~j0 & n5712;
  assign n5714 = m0 & n5713;
  assign n5715 = ~f0 & n5714;
  assign n5716 = ~h0 & n5715;
  assign n5717 = ~e & n5716;
  assign n5718 = ~f & n5717;
  assign n5719 = ~g & n5718;
  assign n5720 = ~i & n5719;
  assign n5721 = ~t & n5720;
  assign n5722 = ~z & n5710;
  assign n5723 = ~a0 & n5722;
  assign n5724 = ~c0 & n5723;
  assign n5725 = ~j0 & n5724;
  assign n5726 = m0 & n5725;
  assign n5727 = ~f0 & n5726;
  assign n5728 = ~e & n5727;
  assign n5729 = ~f & n5728;
  assign n5730 = ~g & n5729;
  assign n5731 = ~i & n5730;
  assign n5732 = ~t & n5731;
  assign n5733 = ~g0 & n5712;
  assign n5734 = ~j0 & n5733;
  assign n5735 = m0 & n5734;
  assign n5736 = ~f0 & n5735;
  assign n5737 = ~h0 & n5736;
  assign n5738 = ~e & n5737;
  assign n5739 = ~f & n5738;
  assign n5740 = ~g & n5739;
  assign n5741 = ~t & n5740;
  assign n5742 = ~g0 & n5724;
  assign n5743 = ~j0 & n5742;
  assign n5744 = m0 & n5743;
  assign n5745 = ~f0 & n5744;
  assign n5746 = ~e & n5745;
  assign n5747 = ~f & n5746;
  assign n5748 = ~g & n5747;
  assign n5749 = ~t & n5748;
  assign n5750 = ~y & n4895;
  assign n5751 = ~c0 & n5750;
  assign n5752 = ~j0 & n5751;
  assign n5753 = m0 & n5752;
  assign n5754 = ~h0 & n5753;
  assign n5755 = ~e & n5754;
  assign n5756 = ~f & n5755;
  assign n5757 = ~g & n5756;
  assign n5758 = ~i & n5757;
  assign n5759 = ~d0 & n5758;
  assign n5760 = i0 & n5759;
  assign n5761 = ~m & n5760;
  assign n5762 = ~k & n5761;
  assign n5763 = ~z & n5750;
  assign n5764 = ~c0 & n5763;
  assign n5765 = ~j0 & n5764;
  assign n5766 = m0 & n5765;
  assign n5767 = ~e & n5766;
  assign n5768 = ~f & n5767;
  assign n5769 = ~g & n5768;
  assign n5770 = ~i & n5769;
  assign n5771 = ~d0 & n5770;
  assign n5772 = i0 & n5771;
  assign n5773 = ~m & n5772;
  assign n5774 = ~k & n5773;
  assign n5775 = ~g0 & n5751;
  assign n5776 = ~j0 & n5775;
  assign n5777 = m0 & n5776;
  assign n5778 = ~h0 & n5777;
  assign n5779 = ~e & n5778;
  assign n5780 = ~f & n5779;
  assign n5781 = ~g & n5780;
  assign n5782 = ~d0 & n5781;
  assign n5783 = i0 & n5782;
  assign n5784 = ~m & n5783;
  assign n5785 = ~k & n5784;
  assign n5786 = ~g0 & n5764;
  assign n5787 = ~j0 & n5786;
  assign n5788 = m0 & n5787;
  assign n5789 = ~e & n5788;
  assign n5790 = ~f & n5789;
  assign n5791 = ~g & n5790;
  assign n5792 = ~d0 & n5791;
  assign n5793 = i0 & n5792;
  assign n5794 = ~m & n5793;
  assign n5795 = ~k & n5794;
  assign n5796 = ~a0 & n5750;
  assign n5797 = ~c0 & n5796;
  assign n5798 = ~j0 & n5797;
  assign n5799 = m0 & n5798;
  assign n5800 = ~h0 & n5799;
  assign n5801 = ~e & n5800;
  assign n5802 = ~f & n5801;
  assign n5803 = ~g & n5802;
  assign n5804 = ~i & n5803;
  assign n5805 = ~d0 & n5804;
  assign n5806 = ~m & n5805;
  assign n5807 = ~k & n5806;
  assign n5808 = ~a0 & n5763;
  assign n5809 = ~c0 & n5808;
  assign n5810 = ~j0 & n5809;
  assign n5811 = m0 & n5810;
  assign n5812 = ~e & n5811;
  assign n5813 = ~f & n5812;
  assign n5814 = ~g & n5813;
  assign n5815 = ~i & n5814;
  assign n5816 = ~d0 & n5815;
  assign n5817 = ~m & n5816;
  assign n5818 = ~k & n5817;
  assign n5819 = ~g0 & n5797;
  assign n5820 = ~j0 & n5819;
  assign n5821 = m0 & n5820;
  assign n5822 = ~h0 & n5821;
  assign n5823 = ~e & n5822;
  assign n5824 = ~f & n5823;
  assign n5825 = ~g & n5824;
  assign n5826 = ~d0 & n5825;
  assign n5827 = ~m & n5826;
  assign n5828 = ~k & n5827;
  assign n5829 = ~g0 & n5809;
  assign n5830 = ~j0 & n5829;
  assign n5831 = m0 & n5830;
  assign n5832 = ~e & n5831;
  assign n5833 = ~f & n5832;
  assign n5834 = ~g & n5833;
  assign n5835 = ~d0 & n5834;
  assign n5836 = ~m & n5835;
  assign n5837 = ~k & n5836;
  assign n5838 = ~w & n4895;
  assign n5839 = ~y & n5838;
  assign n5840 = ~a0 & n5839;
  assign n5841 = ~c0 & n5840;
  assign n5842 = ~j0 & n5841;
  assign n5843 = m0 & n5842;
  assign n5844 = ~h0 & n5843;
  assign n5845 = ~e & n5844;
  assign n5846 = ~f & n5845;
  assign n5847 = ~g & n5846;
  assign n5848 = ~i & n5847;
  assign n5849 = ~m & n5848;
  assign n5850 = ~k & n5849;
  assign n5851 = ~z & n5839;
  assign n5852 = ~a0 & n5851;
  assign n5853 = ~c0 & n5852;
  assign n5854 = ~j0 & n5853;
  assign n5855 = m0 & n5854;
  assign n5856 = ~e & n5855;
  assign n5857 = ~f & n5856;
  assign n5858 = ~g & n5857;
  assign n5859 = ~i & n5858;
  assign n5860 = ~m & n5859;
  assign n5861 = ~k & n5860;
  assign n5862 = ~g0 & n5841;
  assign n5863 = ~j0 & n5862;
  assign n5864 = m0 & n5863;
  assign n5865 = ~h0 & n5864;
  assign n5866 = ~e & n5865;
  assign n5867 = ~f & n5866;
  assign n5868 = ~g & n5867;
  assign n5869 = ~m & n5868;
  assign n5870 = ~k & n5869;
  assign n5871 = ~g0 & n5853;
  assign n5872 = ~j0 & n5871;
  assign n5873 = m0 & n5872;
  assign n5874 = ~e & n5873;
  assign n5875 = ~f & n5874;
  assign n5876 = ~g & n5875;
  assign n5877 = ~m & n5876;
  assign n5878 = ~k & n5877;
  assign n5879 = ~b & n5760;
  assign n5880 = ~k & n5879;
  assign n5881 = ~b & n5772;
  assign n5882 = ~k & n5881;
  assign n5883 = ~b & n5783;
  assign n5884 = ~k & n5883;
  assign n5885 = ~b & n5793;
  assign n5886 = ~k & n5885;
  assign n5887 = ~b & n5805;
  assign n5888 = ~k & n5887;
  assign n5889 = ~b & n5816;
  assign n5890 = ~k & n5889;
  assign n5891 = ~b & n5826;
  assign n5892 = ~k & n5891;
  assign n5893 = ~b & n5835;
  assign n5894 = ~k & n5893;
  assign n5895 = ~b & n5848;
  assign n5896 = ~k & n5895;
  assign n5897 = ~b & n5859;
  assign n5898 = ~k & n5897;
  assign n5899 = ~b & n5868;
  assign n5900 = ~k & n5899;
  assign n5901 = ~b & n5876;
  assign n5902 = ~k & n5901;
  assign n5903 = ~y & n5489;
  assign n5904 = ~c0 & n5903;
  assign n5905 = ~j0 & n5904;
  assign n5906 = m0 & n5905;
  assign n5907 = ~f0 & n5906;
  assign n5908 = ~h0 & n5907;
  assign n5909 = ~e & n5908;
  assign n5910 = ~f & n5909;
  assign n5911 = ~g & n5910;
  assign n5912 = ~i & n5911;
  assign n5913 = ~d0 & n5912;
  assign n5914 = i0 & n5913;
  assign n5915 = ~k & n5914;
  assign n5916 = ~z & n5903;
  assign n5917 = ~c0 & n5916;
  assign n5918 = ~j0 & n5917;
  assign n5919 = m0 & n5918;
  assign n5920 = ~f0 & n5919;
  assign n5921 = ~e & n5920;
  assign n5922 = ~f & n5921;
  assign n5923 = ~g & n5922;
  assign n5924 = ~i & n5923;
  assign n5925 = ~d0 & n5924;
  assign n5926 = i0 & n5925;
  assign n5927 = ~k & n5926;
  assign n5928 = ~g0 & n5904;
  assign n5929 = ~j0 & n5928;
  assign n5930 = m0 & n5929;
  assign n5931 = ~f0 & n5930;
  assign n5932 = ~h0 & n5931;
  assign n5933 = ~e & n5932;
  assign n5934 = ~f & n5933;
  assign n5935 = ~g & n5934;
  assign n5936 = ~d0 & n5935;
  assign n5937 = i0 & n5936;
  assign n5938 = ~k & n5937;
  assign n5939 = ~g0 & n5917;
  assign n5940 = ~j0 & n5939;
  assign n5941 = m0 & n5940;
  assign n5942 = ~f0 & n5941;
  assign n5943 = ~e & n5942;
  assign n5944 = ~f & n5943;
  assign n5945 = ~g & n5944;
  assign n5946 = ~d0 & n5945;
  assign n5947 = i0 & n5946;
  assign n5948 = ~k & n5947;
  assign n5949 = ~a0 & n5903;
  assign n5950 = ~c0 & n5949;
  assign n5951 = ~j0 & n5950;
  assign n5952 = m0 & n5951;
  assign n5953 = ~f0 & n5952;
  assign n5954 = ~h0 & n5953;
  assign n5955 = ~e & n5954;
  assign n5956 = ~f & n5955;
  assign n5957 = ~g & n5956;
  assign n5958 = ~i & n5957;
  assign n5959 = ~d0 & n5958;
  assign n5960 = ~k & n5959;
  assign n5961 = ~a0 & n5916;
  assign n5962 = ~c0 & n5961;
  assign n5963 = ~j0 & n5962;
  assign n5964 = m0 & n5963;
  assign n5965 = ~f0 & n5964;
  assign n5966 = ~e & n5965;
  assign n5967 = ~f & n5966;
  assign n5968 = ~g & n5967;
  assign n5969 = ~i & n5968;
  assign n5970 = ~d0 & n5969;
  assign n5971 = ~k & n5970;
  assign n5972 = ~g0 & n5950;
  assign n5973 = ~j0 & n5972;
  assign n5974 = m0 & n5973;
  assign n5975 = ~f0 & n5974;
  assign n5976 = ~h0 & n5975;
  assign n5977 = ~e & n5976;
  assign n5978 = ~f & n5977;
  assign n5979 = ~g & n5978;
  assign n5980 = ~d0 & n5979;
  assign n5981 = ~k & n5980;
  assign n5982 = ~g0 & n5962;
  assign n5983 = ~j0 & n5982;
  assign n5984 = m0 & n5983;
  assign n5985 = ~f0 & n5984;
  assign n5986 = ~e & n5985;
  assign n5987 = ~f & n5986;
  assign n5988 = ~g & n5987;
  assign n5989 = ~d0 & n5988;
  assign n5990 = ~k & n5989;
  assign n5991 = ~w & n5489;
  assign n5992 = ~y & n5991;
  assign n5993 = ~a0 & n5992;
  assign n5994 = ~c0 & n5993;
  assign n5995 = ~j0 & n5994;
  assign n5996 = m0 & n5995;
  assign n5997 = ~f0 & n5996;
  assign n5998 = ~h0 & n5997;
  assign n5999 = ~e & n5998;
  assign n6000 = ~f & n5999;
  assign n6001 = ~g & n6000;
  assign n6002 = ~i & n6001;
  assign n6003 = ~k & n6002;
  assign n6004 = ~z & n5992;
  assign n6005 = ~a0 & n6004;
  assign n6006 = ~c0 & n6005;
  assign n6007 = ~j0 & n6006;
  assign n6008 = m0 & n6007;
  assign n6009 = ~f0 & n6008;
  assign n6010 = ~e & n6009;
  assign n6011 = ~f & n6010;
  assign n6012 = ~g & n6011;
  assign n6013 = ~i & n6012;
  assign n6014 = ~k & n6013;
  assign n6015 = ~g0 & n5994;
  assign n6016 = ~j0 & n6015;
  assign n6017 = m0 & n6016;
  assign n6018 = ~f0 & n6017;
  assign n6019 = ~h0 & n6018;
  assign n6020 = ~e & n6019;
  assign n6021 = ~f & n6020;
  assign n6022 = ~g & n6021;
  assign n6023 = ~k & n6022;
  assign n6024 = ~g0 & n6006;
  assign n6025 = ~j0 & n6024;
  assign n6026 = m0 & n6025;
  assign n6027 = ~f0 & n6026;
  assign n6028 = ~e & n6027;
  assign n6029 = ~f & n6028;
  assign n6030 = ~g & n6029;
  assign n6031 = ~k & n6030;
  assign n6032 = ~n & ~w;
  assign n6033 = ~y & n6032;
  assign n6034 = ~a0 & n6033;
  assign n6035 = ~c0 & n6034;
  assign n6036 = ~e0 & n6035;
  assign n6037 = ~j0 & n6036;
  assign n6038 = m0 & n6037;
  assign n6039 = ~f0 & n6038;
  assign n6040 = ~h0 & n6039;
  assign n6041 = ~i & n6040;
  assign n6042 = t & n6041;
  assign n6043 = ~d & n6042;
  assign n6044 = m & n6043;
  assign n6045 = k & n6044;
  assign n6046 = ~z & n6033;
  assign n6047 = ~a0 & n6046;
  assign n6048 = ~c0 & n6047;
  assign n6049 = ~e0 & n6048;
  assign n6050 = ~j0 & n6049;
  assign n6051 = m0 & n6050;
  assign n6052 = ~f0 & n6051;
  assign n6053 = ~i & n6052;
  assign n6054 = t & n6053;
  assign n6055 = ~d & n6054;
  assign n6056 = m & n6055;
  assign n6057 = k & n6056;
  assign n6058 = ~g0 & n6036;
  assign n6059 = ~j0 & n6058;
  assign n6060 = m0 & n6059;
  assign n6061 = ~f0 & n6060;
  assign n6062 = ~h0 & n6061;
  assign n6063 = t & n6062;
  assign n6064 = ~d & n6063;
  assign n6065 = m & n6064;
  assign n6066 = k & n6065;
  assign n6067 = ~g0 & n6049;
  assign n6068 = ~j0 & n6067;
  assign n6069 = m0 & n6068;
  assign n6070 = ~f0 & n6069;
  assign n6071 = t & n6070;
  assign n6072 = ~d & n6071;
  assign n6073 = m & n6072;
  assign n6074 = k & n6073;
  assign n6075 = l & ~n;
  assign n6076 = ~w & n6075;
  assign n6077 = ~y & n6076;
  assign n6078 = ~a0 & n6077;
  assign n6079 = ~c0 & n6078;
  assign n6080 = ~e0 & n6079;
  assign n6081 = ~j0 & n6080;
  assign n6082 = m0 & n6081;
  assign n6083 = ~f0 & n6082;
  assign n6084 = ~h0 & n6083;
  assign n6085 = ~i & n6084;
  assign n6086 = ~d & n6085;
  assign n6087 = m & n6086;
  assign n6088 = k & n6087;
  assign n6089 = ~z & n6077;
  assign n6090 = ~a0 & n6089;
  assign n6091 = ~c0 & n6090;
  assign n6092 = ~e0 & n6091;
  assign n6093 = ~j0 & n6092;
  assign n6094 = m0 & n6093;
  assign n6095 = ~f0 & n6094;
  assign n6096 = ~i & n6095;
  assign n6097 = ~d & n6096;
  assign n6098 = m & n6097;
  assign n6099 = k & n6098;
  assign n6100 = ~g0 & n6080;
  assign n6101 = ~j0 & n6100;
  assign n6102 = m0 & n6101;
  assign n6103 = ~f0 & n6102;
  assign n6104 = ~h0 & n6103;
  assign n6105 = ~d & n6104;
  assign n6106 = m & n6105;
  assign n6107 = k & n6106;
  assign n6108 = ~g0 & n6092;
  assign n6109 = ~j0 & n6108;
  assign n6110 = m0 & n6109;
  assign n6111 = ~f0 & n6110;
  assign n6112 = ~d & n6111;
  assign n6113 = m & n6112;
  assign n6114 = k & n6113;
  assign n6115 = ~n & s;
  assign n6116 = ~w & n6115;
  assign n6117 = ~y & n6116;
  assign n6118 = ~a0 & n6117;
  assign n6119 = ~c0 & n6118;
  assign n6120 = ~e0 & n6119;
  assign n6121 = ~j0 & n6120;
  assign n6122 = m0 & n6121;
  assign n6123 = ~f0 & n6122;
  assign n6124 = ~h0 & n6123;
  assign n6125 = ~i & n6124;
  assign n6126 = t & n6125;
  assign n6127 = m & n6126;
  assign n6128 = k & n6127;
  assign n6129 = ~z & n6117;
  assign n6130 = ~a0 & n6129;
  assign n6131 = ~c0 & n6130;
  assign n6132 = ~e0 & n6131;
  assign n6133 = ~j0 & n6132;
  assign n6134 = m0 & n6133;
  assign n6135 = ~f0 & n6134;
  assign n6136 = ~i & n6135;
  assign n6137 = t & n6136;
  assign n6138 = m & n6137;
  assign n6139 = k & n6138;
  assign n6140 = ~g0 & n6120;
  assign n6141 = ~j0 & n6140;
  assign n6142 = m0 & n6141;
  assign n6143 = ~f0 & n6142;
  assign n6144 = ~h0 & n6143;
  assign n6145 = t & n6144;
  assign n6146 = m & n6145;
  assign n6147 = k & n6146;
  assign n6148 = ~g0 & n6132;
  assign n6149 = ~j0 & n6148;
  assign n6150 = m0 & n6149;
  assign n6151 = ~f0 & n6150;
  assign n6152 = t & n6151;
  assign n6153 = m & n6152;
  assign n6154 = k & n6153;
  assign n6155 = s & n6075;
  assign n6156 = ~w & n6155;
  assign n6157 = ~y & n6156;
  assign n6158 = ~a0 & n6157;
  assign n6159 = ~c0 & n6158;
  assign n6160 = ~e0 & n6159;
  assign n6161 = ~j0 & n6160;
  assign n6162 = m0 & n6161;
  assign n6163 = ~f0 & n6162;
  assign n6164 = ~h0 & n6163;
  assign n6165 = ~i & n6164;
  assign n6166 = m & n6165;
  assign n6167 = k & n6166;
  assign n6168 = ~z & n6157;
  assign n6169 = ~a0 & n6168;
  assign n6170 = ~c0 & n6169;
  assign n6171 = ~e0 & n6170;
  assign n6172 = ~j0 & n6171;
  assign n6173 = m0 & n6172;
  assign n6174 = ~f0 & n6173;
  assign n6175 = ~i & n6174;
  assign n6176 = m & n6175;
  assign n6177 = k & n6176;
  assign n6178 = ~g0 & n6160;
  assign n6179 = ~j0 & n6178;
  assign n6180 = m0 & n6179;
  assign n6181 = ~f0 & n6180;
  assign n6182 = ~h0 & n6181;
  assign n6183 = m & n6182;
  assign n6184 = k & n6183;
  assign n6185 = ~g0 & n6171;
  assign n6186 = ~j0 & n6185;
  assign n6187 = m0 & n6186;
  assign n6188 = ~f0 & n6187;
  assign n6189 = m & n6188;
  assign n6190 = k & n6189;
  assign n6191 = ~c0 & n5490;
  assign n6192 = j0 & n6191;
  assign n6193 = m0 & n6192;
  assign n6194 = ~h0 & n6193;
  assign n6195 = ~e & n6194;
  assign n6196 = ~f & n6195;
  assign n6197 = ~g & n6196;
  assign n6198 = ~h & n6197;
  assign n6199 = ~i & n6198;
  assign n6200 = ~d0 & n6199;
  assign n6201 = ~i0 & n6200;
  assign n6202 = d & n6201;
  assign n6203 = ~z & n5490;
  assign n6204 = ~c0 & n6203;
  assign n6205 = j0 & n6204;
  assign n6206 = m0 & n6205;
  assign n6207 = ~e & n6206;
  assign n6208 = ~f & n6207;
  assign n6209 = ~g & n6208;
  assign n6210 = ~h & n6209;
  assign n6211 = ~i & n6210;
  assign n6212 = ~d0 & n6211;
  assign n6213 = ~i0 & n6212;
  assign n6214 = d & n6213;
  assign n6215 = ~g0 & n6191;
  assign n6216 = j0 & n6215;
  assign n6217 = m0 & n6216;
  assign n6218 = ~h0 & n6217;
  assign n6219 = ~e & n6218;
  assign n6220 = ~f & n6219;
  assign n6221 = ~g & n6220;
  assign n6222 = ~h & n6221;
  assign n6223 = ~d0 & n6222;
  assign n6224 = ~i0 & n6223;
  assign n6225 = d & n6224;
  assign n6226 = ~g0 & n6204;
  assign n6227 = j0 & n6226;
  assign n6228 = m0 & n6227;
  assign n6229 = ~e & n6228;
  assign n6230 = ~f & n6229;
  assign n6231 = ~g & n6230;
  assign n6232 = ~h & n6231;
  assign n6233 = ~d0 & n6232;
  assign n6234 = ~i0 & n6233;
  assign n6235 = d & n6234;
  assign n6236 = m0 & n5492;
  assign n6237 = ~h0 & n6236;
  assign n6238 = ~e & n6237;
  assign n6239 = ~f & n6238;
  assign n6240 = ~g & n6239;
  assign n6241 = ~h & n6240;
  assign n6242 = ~i & n6241;
  assign n6243 = ~d0 & n6242;
  assign n6244 = i0 & n6243;
  assign n6245 = d & n6244;
  assign n6246 = m0 & n5505;
  assign n6247 = ~e & n6246;
  assign n6248 = ~f & n6247;
  assign n6249 = ~g & n6248;
  assign n6250 = ~h & n6249;
  assign n6251 = ~i & n6250;
  assign n6252 = ~d0 & n6251;
  assign n6253 = i0 & n6252;
  assign n6254 = d & n6253;
  assign n6255 = m0 & n5516;
  assign n6256 = ~h0 & n6255;
  assign n6257 = ~e & n6256;
  assign n6258 = ~f & n6257;
  assign n6259 = ~g & n6258;
  assign n6260 = ~h & n6259;
  assign n6261 = ~d0 & n6260;
  assign n6262 = i0 & n6261;
  assign n6263 = d & n6262;
  assign n6264 = m0 & n5527;
  assign n6265 = ~e & n6264;
  assign n6266 = ~f & n6265;
  assign n6267 = ~g & n6266;
  assign n6268 = ~h & n6267;
  assign n6269 = ~d0 & n6268;
  assign n6270 = i0 & n6269;
  assign n6271 = d & n6270;
  assign n6272 = m0 & n5538;
  assign n6273 = ~h0 & n6272;
  assign n6274 = ~e & n6273;
  assign n6275 = ~f & n6274;
  assign n6276 = ~g & n6275;
  assign n6277 = ~h & n6276;
  assign n6278 = ~i & n6277;
  assign n6279 = ~d0 & n6278;
  assign n6280 = d & n6279;
  assign n6281 = m0 & n5550;
  assign n6282 = ~e & n6281;
  assign n6283 = ~f & n6282;
  assign n6284 = ~g & n6283;
  assign n6285 = ~h & n6284;
  assign n6286 = ~i & n6285;
  assign n6287 = ~d0 & n6286;
  assign n6288 = d & n6287;
  assign n6289 = m0 & n5560;
  assign n6290 = ~h0 & n6289;
  assign n6291 = ~e & n6290;
  assign n6292 = ~f & n6291;
  assign n6293 = ~g & n6292;
  assign n6294 = ~h & n6293;
  assign n6295 = ~d0 & n6294;
  assign n6296 = d & n6295;
  assign n6297 = m0 & n5570;
  assign n6298 = ~e & n6297;
  assign n6299 = ~f & n6298;
  assign n6300 = ~g & n6299;
  assign n6301 = ~h & n6300;
  assign n6302 = ~d0 & n6301;
  assign n6303 = d & n6302;
  assign n6304 = m0 & n5582;
  assign n6305 = ~h0 & n6304;
  assign n6306 = ~e & n6305;
  assign n6307 = ~f & n6306;
  assign n6308 = ~g & n6307;
  assign n6309 = ~h & n6308;
  assign n6310 = ~i & n6309;
  assign n6311 = d & n6310;
  assign n6312 = m0 & n5594;
  assign n6313 = ~e & n6312;
  assign n6314 = ~f & n6313;
  assign n6315 = ~g & n6314;
  assign n6316 = ~h & n6315;
  assign n6317 = ~i & n6316;
  assign n6318 = d & n6317;
  assign n6319 = m0 & n5603;
  assign n6320 = ~h0 & n6319;
  assign n6321 = ~e & n6320;
  assign n6322 = ~f & n6321;
  assign n6323 = ~g & n6322;
  assign n6324 = ~h & n6323;
  assign n6325 = d & n6324;
  assign n6326 = m0 & n5612;
  assign n6327 = ~e & n6326;
  assign n6328 = ~f & n6327;
  assign n6329 = ~g & n6328;
  assign n6330 = ~h & n6329;
  assign n6331 = d & n6330;
  assign n6332 = ~c0 & n5620;
  assign n6333 = j0 & n6332;
  assign n6334 = m0 & n6333;
  assign n6335 = ~h0 & n6334;
  assign n6336 = ~e & n6335;
  assign n6337 = ~f & n6336;
  assign n6338 = ~g & n6337;
  assign n6339 = ~h & n6338;
  assign n6340 = ~i & n6339;
  assign n6341 = ~t & n6340;
  assign n6342 = ~d0 & n6341;
  assign n6343 = ~i0 & n6342;
  assign n6344 = ~z & n5620;
  assign n6345 = ~c0 & n6344;
  assign n6346 = j0 & n6345;
  assign n6347 = m0 & n6346;
  assign n6348 = ~e & n6347;
  assign n6349 = ~f & n6348;
  assign n6350 = ~g & n6349;
  assign n6351 = ~h & n6350;
  assign n6352 = ~i & n6351;
  assign n6353 = ~t & n6352;
  assign n6354 = ~d0 & n6353;
  assign n6355 = ~i0 & n6354;
  assign n6356 = ~g0 & n6332;
  assign n6357 = j0 & n6356;
  assign n6358 = m0 & n6357;
  assign n6359 = ~h0 & n6358;
  assign n6360 = ~e & n6359;
  assign n6361 = ~f & n6360;
  assign n6362 = ~g & n6361;
  assign n6363 = ~h & n6362;
  assign n6364 = ~t & n6363;
  assign n6365 = ~d0 & n6364;
  assign n6366 = ~i0 & n6365;
  assign n6367 = ~g0 & n6345;
  assign n6368 = j0 & n6367;
  assign n6369 = m0 & n6368;
  assign n6370 = ~e & n6369;
  assign n6371 = ~f & n6370;
  assign n6372 = ~g & n6371;
  assign n6373 = ~h & n6372;
  assign n6374 = ~t & n6373;
  assign n6375 = ~d0 & n6374;
  assign n6376 = ~i0 & n6375;
  assign n6377 = m0 & n5622;
  assign n6378 = ~h0 & n6377;
  assign n6379 = ~e & n6378;
  assign n6380 = ~f & n6379;
  assign n6381 = ~g & n6380;
  assign n6382 = ~h & n6381;
  assign n6383 = ~i & n6382;
  assign n6384 = ~t & n6383;
  assign n6385 = ~d0 & n6384;
  assign n6386 = i0 & n6385;
  assign n6387 = m0 & n5635;
  assign n6388 = ~e & n6387;
  assign n6389 = ~f & n6388;
  assign n6390 = ~g & n6389;
  assign n6391 = ~h & n6390;
  assign n6392 = ~i & n6391;
  assign n6393 = ~t & n6392;
  assign n6394 = ~d0 & n6393;
  assign n6395 = i0 & n6394;
  assign n6396 = m0 & n5646;
  assign n6397 = ~h0 & n6396;
  assign n6398 = ~e & n6397;
  assign n6399 = ~f & n6398;
  assign n6400 = ~g & n6399;
  assign n6401 = ~h & n6400;
  assign n6402 = ~t & n6401;
  assign n6403 = ~d0 & n6402;
  assign n6404 = i0 & n6403;
  assign n6405 = m0 & n5657;
  assign n6406 = ~e & n6405;
  assign n6407 = ~f & n6406;
  assign n6408 = ~g & n6407;
  assign n6409 = ~h & n6408;
  assign n6410 = ~t & n6409;
  assign n6411 = ~d0 & n6410;
  assign n6412 = i0 & n6411;
  assign n6413 = n & n5489;
  assign n6414 = ~y & n6413;
  assign n6415 = ~c0 & n6414;
  assign n6416 = ~j0 & n6415;
  assign n6417 = m0 & n6416;
  assign n6418 = ~f0 & n6417;
  assign n6419 = ~h0 & n6418;
  assign n6420 = ~e & n6419;
  assign n6421 = ~f & n6420;
  assign n6422 = ~g & n6421;
  assign n6423 = ~i & n6422;
  assign n6424 = ~d0 & n6423;
  assign n6425 = i0 & n6424;
  assign n6426 = ~z & n6414;
  assign n6427 = ~c0 & n6426;
  assign n6428 = ~j0 & n6427;
  assign n6429 = m0 & n6428;
  assign n6430 = ~f0 & n6429;
  assign n6431 = ~e & n6430;
  assign n6432 = ~f & n6431;
  assign n6433 = ~g & n6432;
  assign n6434 = ~i & n6433;
  assign n6435 = ~d0 & n6434;
  assign n6436 = i0 & n6435;
  assign n6437 = ~g0 & n6415;
  assign n6438 = ~j0 & n6437;
  assign n6439 = m0 & n6438;
  assign n6440 = ~f0 & n6439;
  assign n6441 = ~h0 & n6440;
  assign n6442 = ~e & n6441;
  assign n6443 = ~f & n6442;
  assign n6444 = ~g & n6443;
  assign n6445 = ~d0 & n6444;
  assign n6446 = i0 & n6445;
  assign n6447 = ~g0 & n6427;
  assign n6448 = ~j0 & n6447;
  assign n6449 = m0 & n6448;
  assign n6450 = ~f0 & n6449;
  assign n6451 = ~e & n6450;
  assign n6452 = ~f & n6451;
  assign n6453 = ~g & n6452;
  assign n6454 = ~d0 & n6453;
  assign n6455 = i0 & n6454;
  assign n6456 = m0 & n5668;
  assign n6457 = ~h0 & n6456;
  assign n6458 = ~e & n6457;
  assign n6459 = ~f & n6458;
  assign n6460 = ~g & n6459;
  assign n6461 = ~h & n6460;
  assign n6462 = ~i & n6461;
  assign n6463 = ~t & n6462;
  assign n6464 = ~d0 & n6463;
  assign n6465 = m0 & n5680;
  assign n6466 = ~e & n6465;
  assign n6467 = ~f & n6466;
  assign n6468 = ~g & n6467;
  assign n6469 = ~h & n6468;
  assign n6470 = ~i & n6469;
  assign n6471 = ~t & n6470;
  assign n6472 = ~d0 & n6471;
  assign n6473 = m0 & n5690;
  assign n6474 = ~h0 & n6473;
  assign n6475 = ~e & n6474;
  assign n6476 = ~f & n6475;
  assign n6477 = ~g & n6476;
  assign n6478 = ~h & n6477;
  assign n6479 = ~t & n6478;
  assign n6480 = ~d0 & n6479;
  assign n6481 = m0 & n5700;
  assign n6482 = ~e & n6481;
  assign n6483 = ~f & n6482;
  assign n6484 = ~g & n6483;
  assign n6485 = ~h & n6484;
  assign n6486 = ~t & n6485;
  assign n6487 = ~d0 & n6486;
  assign n6488 = ~a0 & n6414;
  assign n6489 = ~c0 & n6488;
  assign n6490 = ~j0 & n6489;
  assign n6491 = m0 & n6490;
  assign n6492 = ~f0 & n6491;
  assign n6493 = ~h0 & n6492;
  assign n6494 = ~e & n6493;
  assign n6495 = ~f & n6494;
  assign n6496 = ~g & n6495;
  assign n6497 = ~i & n6496;
  assign n6498 = ~d0 & n6497;
  assign n6499 = ~a0 & n6426;
  assign n6500 = ~c0 & n6499;
  assign n6501 = ~j0 & n6500;
  assign n6502 = m0 & n6501;
  assign n6503 = ~f0 & n6502;
  assign n6504 = ~e & n6503;
  assign n6505 = ~f & n6504;
  assign n6506 = ~g & n6505;
  assign n6507 = ~i & n6506;
  assign n6508 = ~d0 & n6507;
  assign n6509 = ~g0 & n6489;
  assign n6510 = ~j0 & n6509;
  assign n6511 = m0 & n6510;
  assign n6512 = ~f0 & n6511;
  assign n6513 = ~h0 & n6512;
  assign n6514 = ~e & n6513;
  assign n6515 = ~f & n6514;
  assign n6516 = ~g & n6515;
  assign n6517 = ~d0 & n6516;
  assign n6518 = ~g0 & n6500;
  assign n6519 = ~j0 & n6518;
  assign n6520 = m0 & n6519;
  assign n6521 = ~f0 & n6520;
  assign n6522 = ~e & n6521;
  assign n6523 = ~f & n6522;
  assign n6524 = ~g & n6523;
  assign n6525 = ~d0 & n6524;
  assign n6526 = m0 & n5712;
  assign n6527 = ~h0 & n6526;
  assign n6528 = ~e & n6527;
  assign n6529 = ~f & n6528;
  assign n6530 = ~g & n6529;
  assign n6531 = ~h & n6530;
  assign n6532 = ~i & n6531;
  assign n6533 = ~t & n6532;
  assign n6534 = m0 & n5724;
  assign n6535 = ~e & n6534;
  assign n6536 = ~f & n6535;
  assign n6537 = ~g & n6536;
  assign n6538 = ~h & n6537;
  assign n6539 = ~i & n6538;
  assign n6540 = ~t & n6539;
  assign n6541 = m0 & n5733;
  assign n6542 = ~h0 & n6541;
  assign n6543 = ~e & n6542;
  assign n6544 = ~f & n6543;
  assign n6545 = ~g & n6544;
  assign n6546 = ~h & n6545;
  assign n6547 = ~t & n6546;
  assign n6548 = m0 & n5742;
  assign n6549 = ~e & n6548;
  assign n6550 = ~f & n6549;
  assign n6551 = ~g & n6550;
  assign n6552 = ~h & n6551;
  assign n6553 = ~t & n6552;
  assign n6554 = ~w & n6413;
  assign n6555 = ~y & n6554;
  assign n6556 = ~a0 & n6555;
  assign n6557 = ~c0 & n6556;
  assign n6558 = ~j0 & n6557;
  assign n6559 = m0 & n6558;
  assign n6560 = ~f0 & n6559;
  assign n6561 = ~h0 & n6560;
  assign n6562 = ~e & n6561;
  assign n6563 = ~f & n6562;
  assign n6564 = ~g & n6563;
  assign n6565 = ~i & n6564;
  assign n6566 = ~z & n6555;
  assign n6567 = ~a0 & n6566;
  assign n6568 = ~c0 & n6567;
  assign n6569 = ~j0 & n6568;
  assign n6570 = m0 & n6569;
  assign n6571 = ~f0 & n6570;
  assign n6572 = ~e & n6571;
  assign n6573 = ~f & n6572;
  assign n6574 = ~g & n6573;
  assign n6575 = ~i & n6574;
  assign n6576 = ~g0 & n6557;
  assign n6577 = ~j0 & n6576;
  assign n6578 = m0 & n6577;
  assign n6579 = ~f0 & n6578;
  assign n6580 = ~h0 & n6579;
  assign n6581 = ~e & n6580;
  assign n6582 = ~f & n6581;
  assign n6583 = ~g & n6582;
  assign n6584 = ~g0 & n6568;
  assign n6585 = ~j0 & n6584;
  assign n6586 = m0 & n6585;
  assign n6587 = ~f0 & n6586;
  assign n6588 = ~e & n6587;
  assign n6589 = ~f & n6588;
  assign n6590 = ~g & n6589;
  assign n6591 = ~c0 & n5489;
  assign n6592 = j0 & n6591;
  assign n6593 = m0 & n6592;
  assign n6594 = ~h0 & n6593;
  assign n6595 = ~e & n6594;
  assign n6596 = ~f & n6595;
  assign n6597 = ~g & n6596;
  assign n6598 = ~h & n6597;
  assign n6599 = ~i & n6598;
  assign n6600 = ~d0 & n6599;
  assign n6601 = ~i0 & n6600;
  assign n6602 = ~k & n6601;
  assign n6603 = ~z & n5489;
  assign n6604 = ~c0 & n6603;
  assign n6605 = j0 & n6604;
  assign n6606 = m0 & n6605;
  assign n6607 = ~e & n6606;
  assign n6608 = ~f & n6607;
  assign n6609 = ~g & n6608;
  assign n6610 = ~h & n6609;
  assign n6611 = ~i & n6610;
  assign n6612 = ~d0 & n6611;
  assign n6613 = ~i0 & n6612;
  assign n6614 = ~k & n6613;
  assign n6615 = ~g0 & n6591;
  assign n6616 = j0 & n6615;
  assign n6617 = m0 & n6616;
  assign n6618 = ~h0 & n6617;
  assign n6619 = ~e & n6618;
  assign n6620 = ~f & n6619;
  assign n6621 = ~g & n6620;
  assign n6622 = ~h & n6621;
  assign n6623 = ~d0 & n6622;
  assign n6624 = ~i0 & n6623;
  assign n6625 = ~k & n6624;
  assign n6626 = ~g0 & n6604;
  assign n6627 = j0 & n6626;
  assign n6628 = m0 & n6627;
  assign n6629 = ~e & n6628;
  assign n6630 = ~f & n6629;
  assign n6631 = ~g & n6630;
  assign n6632 = ~h & n6631;
  assign n6633 = ~d0 & n6632;
  assign n6634 = ~i0 & n6633;
  assign n6635 = ~k & n6634;
  assign n6636 = m0 & n5904;
  assign n6637 = ~h0 & n6636;
  assign n6638 = ~e & n6637;
  assign n6639 = ~f & n6638;
  assign n6640 = ~g & n6639;
  assign n6641 = ~h & n6640;
  assign n6642 = ~i & n6641;
  assign n6643 = ~d0 & n6642;
  assign n6644 = i0 & n6643;
  assign n6645 = ~k & n6644;
  assign n6646 = m0 & n5917;
  assign n6647 = ~e & n6646;
  assign n6648 = ~f & n6647;
  assign n6649 = ~g & n6648;
  assign n6650 = ~h & n6649;
  assign n6651 = ~i & n6650;
  assign n6652 = ~d0 & n6651;
  assign n6653 = i0 & n6652;
  assign n6654 = ~k & n6653;
  assign n6655 = m0 & n5928;
  assign n6656 = ~h0 & n6655;
  assign n6657 = ~e & n6656;
  assign n6658 = ~f & n6657;
  assign n6659 = ~g & n6658;
  assign n6660 = ~h & n6659;
  assign n6661 = ~d0 & n6660;
  assign n6662 = i0 & n6661;
  assign n6663 = ~k & n6662;
  assign n6664 = m0 & n5939;
  assign n6665 = ~e & n6664;
  assign n6666 = ~f & n6665;
  assign n6667 = ~g & n6666;
  assign n6668 = ~h & n6667;
  assign n6669 = ~d0 & n6668;
  assign n6670 = i0 & n6669;
  assign n6671 = ~k & n6670;
  assign n6672 = m0 & n5950;
  assign n6673 = ~h0 & n6672;
  assign n6674 = ~e & n6673;
  assign n6675 = ~f & n6674;
  assign n6676 = ~g & n6675;
  assign n6677 = ~h & n6676;
  assign n6678 = ~i & n6677;
  assign n6679 = ~d0 & n6678;
  assign n6680 = ~k & n6679;
  assign n6681 = m0 & n5962;
  assign n6682 = ~e & n6681;
  assign n6683 = ~f & n6682;
  assign n6684 = ~g & n6683;
  assign n6685 = ~h & n6684;
  assign n6686 = ~i & n6685;
  assign n6687 = ~d0 & n6686;
  assign n6688 = ~k & n6687;
  assign n6689 = m0 & n5972;
  assign n6690 = ~h0 & n6689;
  assign n6691 = ~e & n6690;
  assign n6692 = ~f & n6691;
  assign n6693 = ~g & n6692;
  assign n6694 = ~h & n6693;
  assign n6695 = ~d0 & n6694;
  assign n6696 = ~k & n6695;
  assign n6697 = m0 & n5982;
  assign n6698 = ~e & n6697;
  assign n6699 = ~f & n6698;
  assign n6700 = ~g & n6699;
  assign n6701 = ~h & n6700;
  assign n6702 = ~d0 & n6701;
  assign n6703 = ~k & n6702;
  assign n6704 = m0 & n5994;
  assign n6705 = ~h0 & n6704;
  assign n6706 = ~e & n6705;
  assign n6707 = ~f & n6706;
  assign n6708 = ~g & n6707;
  assign n6709 = ~h & n6708;
  assign n6710 = ~i & n6709;
  assign n6711 = ~k & n6710;
  assign n6712 = m0 & n6006;
  assign n6713 = ~e & n6712;
  assign n6714 = ~f & n6713;
  assign n6715 = ~g & n6714;
  assign n6716 = ~h & n6715;
  assign n6717 = ~i & n6716;
  assign n6718 = ~k & n6717;
  assign n6719 = m0 & n6015;
  assign n6720 = ~h0 & n6719;
  assign n6721 = ~e & n6720;
  assign n6722 = ~f & n6721;
  assign n6723 = ~g & n6722;
  assign n6724 = ~h & n6723;
  assign n6725 = ~k & n6724;
  assign n6726 = m0 & n6024;
  assign n6727 = ~e & n6726;
  assign n6728 = ~f & n6727;
  assign n6729 = ~g & n6728;
  assign n6730 = ~h & n6729;
  assign n6731 = ~k & n6730;
  assign n6732 = m0 & n6036;
  assign n6733 = ~h0 & n6732;
  assign n6734 = ~h & n6733;
  assign n6735 = ~i & n6734;
  assign n6736 = t & n6735;
  assign n6737 = ~d & n6736;
  assign n6738 = m & n6737;
  assign n6739 = k & n6738;
  assign n6740 = m0 & n6049;
  assign n6741 = ~h & n6740;
  assign n6742 = ~i & n6741;
  assign n6743 = t & n6742;
  assign n6744 = ~d & n6743;
  assign n6745 = m & n6744;
  assign n6746 = k & n6745;
  assign n6747 = m0 & n6058;
  assign n6748 = ~h0 & n6747;
  assign n6749 = ~h & n6748;
  assign n6750 = t & n6749;
  assign n6751 = ~d & n6750;
  assign n6752 = m & n6751;
  assign n6753 = k & n6752;
  assign n6754 = m0 & n6067;
  assign n6755 = ~h & n6754;
  assign n6756 = t & n6755;
  assign n6757 = ~d & n6756;
  assign n6758 = m & n6757;
  assign n6759 = k & n6758;
  assign n6760 = m0 & n6080;
  assign n6761 = ~h0 & n6760;
  assign n6762 = ~h & n6761;
  assign n6763 = ~i & n6762;
  assign n6764 = ~d & n6763;
  assign n6765 = m & n6764;
  assign n6766 = k & n6765;
  assign n6767 = m0 & n6092;
  assign n6768 = ~h & n6767;
  assign n6769 = ~i & n6768;
  assign n6770 = ~d & n6769;
  assign n6771 = m & n6770;
  assign n6772 = k & n6771;
  assign n6773 = m0 & n6100;
  assign n6774 = ~h0 & n6773;
  assign n6775 = ~h & n6774;
  assign n6776 = ~d & n6775;
  assign n6777 = m & n6776;
  assign n6778 = k & n6777;
  assign n6779 = m0 & n6108;
  assign n6780 = ~h & n6779;
  assign n6781 = ~d & n6780;
  assign n6782 = m & n6781;
  assign n6783 = k & n6782;
  assign n6784 = m0 & n6120;
  assign n6785 = ~h0 & n6784;
  assign n6786 = ~h & n6785;
  assign n6787 = ~i & n6786;
  assign n6788 = t & n6787;
  assign n6789 = m & n6788;
  assign n6790 = k & n6789;
  assign n6791 = m0 & n6132;
  assign n6792 = ~h & n6791;
  assign n6793 = ~i & n6792;
  assign n6794 = t & n6793;
  assign n6795 = m & n6794;
  assign n6796 = k & n6795;
  assign n6797 = m0 & n6140;
  assign n6798 = ~h0 & n6797;
  assign n6799 = ~h & n6798;
  assign n6800 = t & n6799;
  assign n6801 = m & n6800;
  assign n6802 = k & n6801;
  assign n6803 = m0 & n6148;
  assign n6804 = ~h & n6803;
  assign n6805 = t & n6804;
  assign n6806 = m & n6805;
  assign n6807 = k & n6806;
  assign n6808 = m0 & n6160;
  assign n6809 = ~h0 & n6808;
  assign n6810 = ~h & n6809;
  assign n6811 = ~i & n6810;
  assign n6812 = m & n6811;
  assign n6813 = k & n6812;
  assign n6814 = m0 & n6171;
  assign n6815 = ~h & n6814;
  assign n6816 = ~i & n6815;
  assign n6817 = m & n6816;
  assign n6818 = k & n6817;
  assign n6819 = m0 & n6178;
  assign n6820 = ~h0 & n6819;
  assign n6821 = ~h & n6820;
  assign n6822 = m & n6821;
  assign n6823 = k & n6822;
  assign n6824 = m0 & n6185;
  assign n6825 = ~h & n6824;
  assign n6826 = m & n6825;
  assign n6827 = k & n6826;
  assign n6828 = ~c & ~y;
  assign n6829 = ~c0 & n6828;
  assign n6830 = ~j0 & n6829;
  assign n6831 = m0 & n6830;
  assign n6832 = ~f0 & n6831;
  assign n6833 = ~h0 & n6832;
  assign n6834 = ~e & n6833;
  assign n6835 = ~f & n6834;
  assign n6836 = ~g & n6835;
  assign n6837 = ~i & n6836;
  assign n6838 = ~d0 & n6837;
  assign n6839 = i0 & n6838;
  assign n6840 = ~m & n6839;
  assign n6841 = ~z & n6828;
  assign n6842 = ~c0 & n6841;
  assign n6843 = ~j0 & n6842;
  assign n6844 = m0 & n6843;
  assign n6845 = ~f0 & n6844;
  assign n6846 = ~e & n6845;
  assign n6847 = ~f & n6846;
  assign n6848 = ~g & n6847;
  assign n6849 = ~i & n6848;
  assign n6850 = ~d0 & n6849;
  assign n6851 = i0 & n6850;
  assign n6852 = ~m & n6851;
  assign n6853 = ~g0 & n6829;
  assign n6854 = ~j0 & n6853;
  assign n6855 = m0 & n6854;
  assign n6856 = ~f0 & n6855;
  assign n6857 = ~h0 & n6856;
  assign n6858 = ~e & n6857;
  assign n6859 = ~f & n6858;
  assign n6860 = ~g & n6859;
  assign n6861 = ~d0 & n6860;
  assign n6862 = i0 & n6861;
  assign n6863 = ~m & n6862;
  assign n6864 = ~g0 & n6842;
  assign n6865 = ~j0 & n6864;
  assign n6866 = m0 & n6865;
  assign n6867 = ~f0 & n6866;
  assign n6868 = ~e & n6867;
  assign n6869 = ~f & n6868;
  assign n6870 = ~g & n6869;
  assign n6871 = ~d0 & n6870;
  assign n6872 = i0 & n6871;
  assign n6873 = ~m & n6872;
  assign n6874 = ~a0 & n6828;
  assign n6875 = ~c0 & n6874;
  assign n6876 = ~j0 & n6875;
  assign n6877 = m0 & n6876;
  assign n6878 = ~f0 & n6877;
  assign n6879 = ~h0 & n6878;
  assign n6880 = ~e & n6879;
  assign n6881 = ~f & n6880;
  assign n6882 = ~g & n6881;
  assign n6883 = ~i & n6882;
  assign n6884 = ~d0 & n6883;
  assign n6885 = ~m & n6884;
  assign n6886 = ~a0 & n6841;
  assign n6887 = ~c0 & n6886;
  assign n6888 = ~j0 & n6887;
  assign n6889 = m0 & n6888;
  assign n6890 = ~f0 & n6889;
  assign n6891 = ~e & n6890;
  assign n6892 = ~f & n6891;
  assign n6893 = ~g & n6892;
  assign n6894 = ~i & n6893;
  assign n6895 = ~d0 & n6894;
  assign n6896 = ~m & n6895;
  assign n6897 = ~g0 & n6875;
  assign n6898 = ~j0 & n6897;
  assign n6899 = m0 & n6898;
  assign n6900 = ~f0 & n6899;
  assign n6901 = ~h0 & n6900;
  assign n6902 = ~e & n6901;
  assign n6903 = ~f & n6902;
  assign n6904 = ~g & n6903;
  assign n6905 = ~d0 & n6904;
  assign n6906 = ~m & n6905;
  assign n6907 = ~g0 & n6887;
  assign n6908 = ~j0 & n6907;
  assign n6909 = m0 & n6908;
  assign n6910 = ~f0 & n6909;
  assign n6911 = ~e & n6910;
  assign n6912 = ~f & n6911;
  assign n6913 = ~g & n6912;
  assign n6914 = ~d0 & n6913;
  assign n6915 = ~m & n6914;
  assign n6916 = ~c & ~w;
  assign n6917 = ~y & n6916;
  assign n6918 = ~a0 & n6917;
  assign n6919 = ~c0 & n6918;
  assign n6920 = ~j0 & n6919;
  assign n6921 = m0 & n6920;
  assign n6922 = ~f0 & n6921;
  assign n6923 = ~h0 & n6922;
  assign n6924 = ~e & n6923;
  assign n6925 = ~f & n6924;
  assign n6926 = ~g & n6925;
  assign n6927 = ~i & n6926;
  assign n6928 = ~m & n6927;
  assign n6929 = ~z & n6917;
  assign n6930 = ~a0 & n6929;
  assign n6931 = ~c0 & n6930;
  assign n6932 = ~j0 & n6931;
  assign n6933 = m0 & n6932;
  assign n6934 = ~f0 & n6933;
  assign n6935 = ~e & n6934;
  assign n6936 = ~f & n6935;
  assign n6937 = ~g & n6936;
  assign n6938 = ~i & n6937;
  assign n6939 = ~m & n6938;
  assign n6940 = ~g0 & n6919;
  assign n6941 = ~j0 & n6940;
  assign n6942 = m0 & n6941;
  assign n6943 = ~f0 & n6942;
  assign n6944 = ~h0 & n6943;
  assign n6945 = ~e & n6944;
  assign n6946 = ~f & n6945;
  assign n6947 = ~g & n6946;
  assign n6948 = ~m & n6947;
  assign n6949 = ~g0 & n6931;
  assign n6950 = ~j0 & n6949;
  assign n6951 = m0 & n6950;
  assign n6952 = ~f0 & n6951;
  assign n6953 = ~e & n6952;
  assign n6954 = ~f & n6953;
  assign n6955 = ~g & n6954;
  assign n6956 = ~m & n6955;
  assign n6957 = j & ~n;
  assign n6958 = ~w & n6957;
  assign n6959 = ~y & n6958;
  assign n6960 = ~a0 & n6959;
  assign n6961 = ~c0 & n6960;
  assign n6962 = ~e0 & n6961;
  assign n6963 = ~j0 & n6962;
  assign n6964 = m0 & n6963;
  assign n6965 = ~h0 & n6964;
  assign n6966 = ~i & n6965;
  assign n6967 = t & n6966;
  assign n6968 = ~d & n6967;
  assign n6969 = m & n6968;
  assign n6970 = ~z & n6959;
  assign n6971 = ~a0 & n6970;
  assign n6972 = ~c0 & n6971;
  assign n6973 = ~e0 & n6972;
  assign n6974 = ~j0 & n6973;
  assign n6975 = m0 & n6974;
  assign n6976 = ~i & n6975;
  assign n6977 = t & n6976;
  assign n6978 = ~d & n6977;
  assign n6979 = m & n6978;
  assign n6980 = ~g0 & n6962;
  assign n6981 = ~j0 & n6980;
  assign n6982 = m0 & n6981;
  assign n6983 = ~h0 & n6982;
  assign n6984 = t & n6983;
  assign n6985 = ~d & n6984;
  assign n6986 = m & n6985;
  assign n6987 = ~g0 & n6973;
  assign n6988 = ~j0 & n6987;
  assign n6989 = m0 & n6988;
  assign n6990 = t & n6989;
  assign n6991 = ~d & n6990;
  assign n6992 = m & n6991;
  assign n6993 = j & l;
  assign n6994 = ~n & n6993;
  assign n6995 = ~w & n6994;
  assign n6996 = ~y & n6995;
  assign n6997 = ~a0 & n6996;
  assign n6998 = ~c0 & n6997;
  assign n6999 = ~e0 & n6998;
  assign n7000 = ~j0 & n6999;
  assign n7001 = m0 & n7000;
  assign n7002 = ~h0 & n7001;
  assign n7003 = ~i & n7002;
  assign n7004 = ~d & n7003;
  assign n7005 = m & n7004;
  assign n7006 = ~z & n6996;
  assign n7007 = ~a0 & n7006;
  assign n7008 = ~c0 & n7007;
  assign n7009 = ~e0 & n7008;
  assign n7010 = ~j0 & n7009;
  assign n7011 = m0 & n7010;
  assign n7012 = ~i & n7011;
  assign n7013 = ~d & n7012;
  assign n7014 = m & n7013;
  assign n7015 = ~g0 & n6999;
  assign n7016 = ~j0 & n7015;
  assign n7017 = m0 & n7016;
  assign n7018 = ~h0 & n7017;
  assign n7019 = ~d & n7018;
  assign n7020 = m & n7019;
  assign n7021 = ~g0 & n7009;
  assign n7022 = ~j0 & n7021;
  assign n7023 = m0 & n7022;
  assign n7024 = ~d & n7023;
  assign n7025 = m & n7024;
  assign n7026 = s & n6957;
  assign n7027 = ~w & n7026;
  assign n7028 = ~y & n7027;
  assign n7029 = ~a0 & n7028;
  assign n7030 = ~c0 & n7029;
  assign n7031 = ~e0 & n7030;
  assign n7032 = ~j0 & n7031;
  assign n7033 = m0 & n7032;
  assign n7034 = ~h0 & n7033;
  assign n7035 = ~i & n7034;
  assign n7036 = t & n7035;
  assign n7037 = m & n7036;
  assign n7038 = ~z & n7028;
  assign n7039 = ~a0 & n7038;
  assign n7040 = ~c0 & n7039;
  assign n7041 = ~e0 & n7040;
  assign n7042 = ~j0 & n7041;
  assign n7043 = m0 & n7042;
  assign n7044 = ~i & n7043;
  assign n7045 = t & n7044;
  assign n7046 = m & n7045;
  assign n7047 = ~g0 & n7031;
  assign n7048 = ~j0 & n7047;
  assign n7049 = m0 & n7048;
  assign n7050 = ~h0 & n7049;
  assign n7051 = t & n7050;
  assign n7052 = m & n7051;
  assign n7053 = ~g0 & n7041;
  assign n7054 = ~j0 & n7053;
  assign n7055 = m0 & n7054;
  assign n7056 = t & n7055;
  assign n7057 = m & n7056;
  assign n7058 = s & n6994;
  assign n7059 = ~w & n7058;
  assign n7060 = ~y & n7059;
  assign n7061 = ~a0 & n7060;
  assign n7062 = ~c0 & n7061;
  assign n7063 = ~e0 & n7062;
  assign n7064 = ~j0 & n7063;
  assign n7065 = m0 & n7064;
  assign n7066 = ~h0 & n7065;
  assign n7067 = ~i & n7066;
  assign n7068 = m & n7067;
  assign n7069 = ~z & n7060;
  assign n7070 = ~a0 & n7069;
  assign n7071 = ~c0 & n7070;
  assign n7072 = ~e0 & n7071;
  assign n7073 = ~j0 & n7072;
  assign n7074 = m0 & n7073;
  assign n7075 = ~i & n7074;
  assign n7076 = m & n7075;
  assign n7077 = ~g0 & n7063;
  assign n7078 = ~j0 & n7077;
  assign n7079 = m0 & n7078;
  assign n7080 = ~h0 & n7079;
  assign n7081 = m & n7080;
  assign n7082 = ~g0 & n7072;
  assign n7083 = ~j0 & n7082;
  assign n7084 = m0 & n7083;
  assign n7085 = m & n7084;
  assign n7086 = ~e0 & n5086;
  assign n7087 = ~j0 & n7086;
  assign n7088 = m0 & n7087;
  assign n7089 = ~h0 & n7088;
  assign n7090 = ~i & n7089;
  assign n7091 = t & n7090;
  assign n7092 = ~d & n7091;
  assign n7093 = ~e0 & n5099;
  assign n7094 = ~j0 & n7093;
  assign n7095 = m0 & n7094;
  assign n7096 = ~i & n7095;
  assign n7097 = t & n7096;
  assign n7098 = ~d & n7097;
  assign n7099 = ~g0 & n7086;
  assign n7100 = ~j0 & n7099;
  assign n7101 = m0 & n7100;
  assign n7102 = ~h0 & n7101;
  assign n7103 = t & n7102;
  assign n7104 = ~d & n7103;
  assign n7105 = ~g0 & n7093;
  assign n7106 = ~j0 & n7105;
  assign n7107 = m0 & n7106;
  assign n7108 = t & n7107;
  assign n7109 = ~d & n7108;
  assign n7110 = ~e0 & n5131;
  assign n7111 = ~j0 & n7110;
  assign n7112 = m0 & n7111;
  assign n7113 = ~h0 & n7112;
  assign n7114 = ~i & n7113;
  assign n7115 = ~d & n7114;
  assign n7116 = ~e0 & n5143;
  assign n7117 = ~j0 & n7116;
  assign n7118 = m0 & n7117;
  assign n7119 = ~i & n7118;
  assign n7120 = ~d & n7119;
  assign n7121 = ~g0 & n7110;
  assign n7122 = ~j0 & n7121;
  assign n7123 = m0 & n7122;
  assign n7124 = ~h0 & n7123;
  assign n7125 = ~d & n7124;
  assign n7126 = ~g0 & n7116;
  assign n7127 = ~j0 & n7126;
  assign n7128 = m0 & n7127;
  assign n7129 = ~d & n7128;
  assign n7130 = ~b & n6839;
  assign n7131 = ~b & n6851;
  assign n7132 = ~b & n6862;
  assign n7133 = ~b & n6872;
  assign n7134 = ~b & n6884;
  assign n7135 = ~b & n6895;
  assign n7136 = ~b & n6905;
  assign n7137 = ~b & n6914;
  assign n7138 = ~b & n6927;
  assign n7139 = ~b & n6938;
  assign n7140 = ~b & n6947;
  assign n7141 = ~b & n6955;
  assign n7142 = ~c0 & n6413;
  assign n7143 = j0 & n7142;
  assign n7144 = m0 & n7143;
  assign n7145 = ~h0 & n7144;
  assign n7146 = ~e & n7145;
  assign n7147 = ~f & n7146;
  assign n7148 = ~g & n7147;
  assign n7149 = ~h & n7148;
  assign n7150 = ~i & n7149;
  assign n7151 = ~d0 & n7150;
  assign n7152 = ~i0 & n7151;
  assign n7153 = ~z & n6413;
  assign n7154 = ~c0 & n7153;
  assign n7155 = j0 & n7154;
  assign n7156 = m0 & n7155;
  assign n7157 = ~e & n7156;
  assign n7158 = ~f & n7157;
  assign n7159 = ~g & n7158;
  assign n7160 = ~h & n7159;
  assign n7161 = ~i & n7160;
  assign n7162 = ~d0 & n7161;
  assign n7163 = ~i0 & n7162;
  assign n7164 = ~g0 & n7142;
  assign n7165 = j0 & n7164;
  assign n7166 = m0 & n7165;
  assign n7167 = ~h0 & n7166;
  assign n7168 = ~e & n7167;
  assign n7169 = ~f & n7168;
  assign n7170 = ~g & n7169;
  assign n7171 = ~h & n7170;
  assign n7172 = ~d0 & n7171;
  assign n7173 = ~i0 & n7172;
  assign n7174 = ~g0 & n7154;
  assign n7175 = j0 & n7174;
  assign n7176 = m0 & n7175;
  assign n7177 = ~e & n7176;
  assign n7178 = ~f & n7177;
  assign n7179 = ~g & n7178;
  assign n7180 = ~h & n7179;
  assign n7181 = ~d0 & n7180;
  assign n7182 = ~i0 & n7181;
  assign n7183 = m0 & n6415;
  assign n7184 = ~h0 & n7183;
  assign n7185 = ~e & n7184;
  assign n7186 = ~f & n7185;
  assign n7187 = ~g & n7186;
  assign n7188 = ~h & n7187;
  assign n7189 = ~i & n7188;
  assign n7190 = ~d0 & n7189;
  assign n7191 = i0 & n7190;
  assign n7192 = m0 & n6427;
  assign n7193 = ~e & n7192;
  assign n7194 = ~f & n7193;
  assign n7195 = ~g & n7194;
  assign n7196 = ~h & n7195;
  assign n7197 = ~i & n7196;
  assign n7198 = ~d0 & n7197;
  assign n7199 = i0 & n7198;
  assign n7200 = m0 & n6437;
  assign n7201 = ~h0 & n7200;
  assign n7202 = ~e & n7201;
  assign n7203 = ~f & n7202;
  assign n7204 = ~g & n7203;
  assign n7205 = ~h & n7204;
  assign n7206 = ~d0 & n7205;
  assign n7207 = i0 & n7206;
  assign n7208 = m0 & n6447;
  assign n7209 = ~e & n7208;
  assign n7210 = ~f & n7209;
  assign n7211 = ~g & n7210;
  assign n7212 = ~h & n7211;
  assign n7213 = ~d0 & n7212;
  assign n7214 = i0 & n7213;
  assign n7215 = m0 & n6489;
  assign n7216 = ~h0 & n7215;
  assign n7217 = ~e & n7216;
  assign n7218 = ~f & n7217;
  assign n7219 = ~g & n7218;
  assign n7220 = ~h & n7219;
  assign n7221 = ~i & n7220;
  assign n7222 = ~d0 & n7221;
  assign n7223 = m0 & n6500;
  assign n7224 = ~e & n7223;
  assign n7225 = ~f & n7224;
  assign n7226 = ~g & n7225;
  assign n7227 = ~h & n7226;
  assign n7228 = ~i & n7227;
  assign n7229 = ~d0 & n7228;
  assign n7230 = m0 & n6509;
  assign n7231 = ~h0 & n7230;
  assign n7232 = ~e & n7231;
  assign n7233 = ~f & n7232;
  assign n7234 = ~g & n7233;
  assign n7235 = ~h & n7234;
  assign n7236 = ~d0 & n7235;
  assign n7237 = m0 & n6518;
  assign n7238 = ~e & n7237;
  assign n7239 = ~f & n7238;
  assign n7240 = ~g & n7239;
  assign n7241 = ~h & n7240;
  assign n7242 = ~d0 & n7241;
  assign n7243 = ~e0 & n5342;
  assign n7244 = ~j0 & n7243;
  assign n7245 = m0 & n7244;
  assign n7246 = ~h0 & n7245;
  assign n7247 = ~i & n7246;
  assign n7248 = t & n7247;
  assign n7249 = ~e0 & n5354;
  assign n7250 = ~j0 & n7249;
  assign n7251 = m0 & n7250;
  assign n7252 = ~i & n7251;
  assign n7253 = t & n7252;
  assign n7254 = ~g0 & n7243;
  assign n7255 = ~j0 & n7254;
  assign n7256 = m0 & n7255;
  assign n7257 = ~h0 & n7256;
  assign n7258 = t & n7257;
  assign n7259 = ~g0 & n7249;
  assign n7260 = ~j0 & n7259;
  assign n7261 = m0 & n7260;
  assign n7262 = t & n7261;
  assign n7263 = m0 & n6557;
  assign n7264 = ~h0 & n7263;
  assign n7265 = ~e & n7264;
  assign n7266 = ~f & n7265;
  assign n7267 = ~g & n7266;
  assign n7268 = ~h & n7267;
  assign n7269 = ~i & n7268;
  assign n7270 = m0 & n6568;
  assign n7271 = ~e & n7270;
  assign n7272 = ~f & n7271;
  assign n7273 = ~g & n7272;
  assign n7274 = ~h & n7273;
  assign n7275 = ~i & n7274;
  assign n7276 = ~e0 & n5383;
  assign n7277 = ~j0 & n7276;
  assign n7278 = m0 & n7277;
  assign n7279 = ~h0 & n7278;
  assign n7280 = ~i & n7279;
  assign n7281 = ~e0 & n5394;
  assign n7282 = ~j0 & n7281;
  assign n7283 = m0 & n7282;
  assign n7284 = ~i & n7283;
  assign n7285 = m0 & n6576;
  assign n7286 = ~h0 & n7285;
  assign n7287 = ~e & n7286;
  assign n7288 = ~f & n7287;
  assign n7289 = ~g & n7288;
  assign n7290 = ~h & n7289;
  assign n7291 = m0 & n6584;
  assign n7292 = ~e & n7291;
  assign n7293 = ~f & n7292;
  assign n7294 = ~g & n7293;
  assign n7295 = ~h & n7294;
  assign n7296 = ~g0 & n7276;
  assign n7297 = ~j0 & n7296;
  assign n7298 = m0 & n7297;
  assign n7299 = ~h0 & n7298;
  assign n7300 = ~g0 & n7281;
  assign n7301 = ~j0 & n7300;
  assign n7302 = m0 & n7301;
  assign n7303 = ~c & ~c0;
  assign n7304 = j0 & n7303;
  assign n7305 = m0 & n7304;
  assign n7306 = ~h0 & n7305;
  assign n7307 = ~e & n7306;
  assign n7308 = ~f & n7307;
  assign n7309 = ~g & n7308;
  assign n7310 = ~h & n7309;
  assign n7311 = ~i & n7310;
  assign n7312 = ~d0 & n7311;
  assign n7313 = ~i0 & n7312;
  assign n7314 = ~m & n7313;
  assign n7315 = ~c & ~z;
  assign n7316 = ~c0 & n7315;
  assign n7317 = j0 & n7316;
  assign n7318 = m0 & n7317;
  assign n7319 = ~e & n7318;
  assign n7320 = ~f & n7319;
  assign n7321 = ~g & n7320;
  assign n7322 = ~h & n7321;
  assign n7323 = ~i & n7322;
  assign n7324 = ~d0 & n7323;
  assign n7325 = ~i0 & n7324;
  assign n7326 = ~m & n7325;
  assign n7327 = ~g0 & n7303;
  assign n7328 = j0 & n7327;
  assign n7329 = m0 & n7328;
  assign n7330 = ~h0 & n7329;
  assign n7331 = ~e & n7330;
  assign n7332 = ~f & n7331;
  assign n7333 = ~g & n7332;
  assign n7334 = ~h & n7333;
  assign n7335 = ~d0 & n7334;
  assign n7336 = ~i0 & n7335;
  assign n7337 = ~m & n7336;
  assign n7338 = ~g0 & n7316;
  assign n7339 = j0 & n7338;
  assign n7340 = m0 & n7339;
  assign n7341 = ~e & n7340;
  assign n7342 = ~f & n7341;
  assign n7343 = ~g & n7342;
  assign n7344 = ~h & n7343;
  assign n7345 = ~d0 & n7344;
  assign n7346 = ~i0 & n7345;
  assign n7347 = ~m & n7346;
  assign n7348 = m0 & n6829;
  assign n7349 = ~h0 & n7348;
  assign n7350 = ~e & n7349;
  assign n7351 = ~f & n7350;
  assign n7352 = ~g & n7351;
  assign n7353 = ~h & n7352;
  assign n7354 = ~i & n7353;
  assign n7355 = ~d0 & n7354;
  assign n7356 = i0 & n7355;
  assign n7357 = ~m & n7356;
  assign n7358 = m0 & n6842;
  assign n7359 = ~e & n7358;
  assign n7360 = ~f & n7359;
  assign n7361 = ~g & n7360;
  assign n7362 = ~h & n7361;
  assign n7363 = ~i & n7362;
  assign n7364 = ~d0 & n7363;
  assign n7365 = i0 & n7364;
  assign n7366 = ~m & n7365;
  assign n7367 = m0 & n6853;
  assign n7368 = ~h0 & n7367;
  assign n7369 = ~e & n7368;
  assign n7370 = ~f & n7369;
  assign n7371 = ~g & n7370;
  assign n7372 = ~h & n7371;
  assign n7373 = ~d0 & n7372;
  assign n7374 = i0 & n7373;
  assign n7375 = ~m & n7374;
  assign n7376 = m0 & n6864;
  assign n7377 = ~e & n7376;
  assign n7378 = ~f & n7377;
  assign n7379 = ~g & n7378;
  assign n7380 = ~h & n7379;
  assign n7381 = ~d0 & n7380;
  assign n7382 = i0 & n7381;
  assign n7383 = ~m & n7382;
  assign n7384 = m0 & n6875;
  assign n7385 = ~h0 & n7384;
  assign n7386 = ~e & n7385;
  assign n7387 = ~f & n7386;
  assign n7388 = ~g & n7387;
  assign n7389 = ~h & n7388;
  assign n7390 = ~i & n7389;
  assign n7391 = ~d0 & n7390;
  assign n7392 = ~m & n7391;
  assign n7393 = m0 & n6887;
  assign n7394 = ~e & n7393;
  assign n7395 = ~f & n7394;
  assign n7396 = ~g & n7395;
  assign n7397 = ~h & n7396;
  assign n7398 = ~i & n7397;
  assign n7399 = ~d0 & n7398;
  assign n7400 = ~m & n7399;
  assign n7401 = m0 & n6897;
  assign n7402 = ~h0 & n7401;
  assign n7403 = ~e & n7402;
  assign n7404 = ~f & n7403;
  assign n7405 = ~g & n7404;
  assign n7406 = ~h & n7405;
  assign n7407 = ~d0 & n7406;
  assign n7408 = ~m & n7407;
  assign n7409 = m0 & n6907;
  assign n7410 = ~e & n7409;
  assign n7411 = ~f & n7410;
  assign n7412 = ~g & n7411;
  assign n7413 = ~h & n7412;
  assign n7414 = ~d0 & n7413;
  assign n7415 = ~m & n7414;
  assign n7416 = m0 & n6919;
  assign n7417 = ~h0 & n7416;
  assign n7418 = ~e & n7417;
  assign n7419 = ~f & n7418;
  assign n7420 = ~g & n7419;
  assign n7421 = ~h & n7420;
  assign n7422 = ~i & n7421;
  assign n7423 = ~m & n7422;
  assign n7424 = m0 & n6931;
  assign n7425 = ~e & n7424;
  assign n7426 = ~f & n7425;
  assign n7427 = ~g & n7426;
  assign n7428 = ~h & n7427;
  assign n7429 = ~i & n7428;
  assign n7430 = ~m & n7429;
  assign n7431 = m0 & n6940;
  assign n7432 = ~h0 & n7431;
  assign n7433 = ~e & n7432;
  assign n7434 = ~f & n7433;
  assign n7435 = ~g & n7434;
  assign n7436 = ~h & n7435;
  assign n7437 = ~m & n7436;
  assign n7438 = m0 & n6949;
  assign n7439 = ~e & n7438;
  assign n7440 = ~f & n7439;
  assign n7441 = ~g & n7440;
  assign n7442 = ~h & n7441;
  assign n7443 = ~m & n7442;
  assign n7444 = ~y & n6957;
  assign n7445 = ~c0 & n7444;
  assign n7446 = ~e0 & n7445;
  assign n7447 = ~j0 & n7446;
  assign n7448 = m0 & n7447;
  assign n7449 = ~h0 & n7448;
  assign n7450 = ~i & n7449;
  assign n7451 = t & n7450;
  assign n7452 = ~d0 & n7451;
  assign n7453 = i0 & n7452;
  assign n7454 = ~d & n7453;
  assign n7455 = ~z & n7444;
  assign n7456 = ~c0 & n7455;
  assign n7457 = ~e0 & n7456;
  assign n7458 = ~j0 & n7457;
  assign n7459 = m0 & n7458;
  assign n7460 = ~i & n7459;
  assign n7461 = t & n7460;
  assign n7462 = ~d0 & n7461;
  assign n7463 = i0 & n7462;
  assign n7464 = ~d & n7463;
  assign n7465 = ~g0 & n7446;
  assign n7466 = ~j0 & n7465;
  assign n7467 = m0 & n7466;
  assign n7468 = ~h0 & n7467;
  assign n7469 = t & n7468;
  assign n7470 = ~d0 & n7469;
  assign n7471 = i0 & n7470;
  assign n7472 = ~d & n7471;
  assign n7473 = ~g0 & n7457;
  assign n7474 = ~j0 & n7473;
  assign n7475 = m0 & n7474;
  assign n7476 = t & n7475;
  assign n7477 = ~d0 & n7476;
  assign n7478 = i0 & n7477;
  assign n7479 = ~d & n7478;
  assign n7480 = ~y & n6994;
  assign n7481 = ~c0 & n7480;
  assign n7482 = ~e0 & n7481;
  assign n7483 = ~j0 & n7482;
  assign n7484 = m0 & n7483;
  assign n7485 = ~h0 & n7484;
  assign n7486 = ~i & n7485;
  assign n7487 = ~d0 & n7486;
  assign n7488 = i0 & n7487;
  assign n7489 = ~d & n7488;
  assign n7490 = ~z & n7480;
  assign n7491 = ~c0 & n7490;
  assign n7492 = ~e0 & n7491;
  assign n7493 = ~j0 & n7492;
  assign n7494 = m0 & n7493;
  assign n7495 = ~i & n7494;
  assign n7496 = ~d0 & n7495;
  assign n7497 = i0 & n7496;
  assign n7498 = ~d & n7497;
  assign n7499 = ~g0 & n7482;
  assign n7500 = ~j0 & n7499;
  assign n7501 = m0 & n7500;
  assign n7502 = ~h0 & n7501;
  assign n7503 = ~d0 & n7502;
  assign n7504 = i0 & n7503;
  assign n7505 = ~d & n7504;
  assign n7506 = ~g0 & n7492;
  assign n7507 = ~j0 & n7506;
  assign n7508 = m0 & n7507;
  assign n7509 = ~d0 & n7508;
  assign n7510 = i0 & n7509;
  assign n7511 = ~d & n7510;
  assign n7512 = ~a0 & n7444;
  assign n7513 = ~c0 & n7512;
  assign n7514 = ~e0 & n7513;
  assign n7515 = ~j0 & n7514;
  assign n7516 = m0 & n7515;
  assign n7517 = ~h0 & n7516;
  assign n7518 = ~i & n7517;
  assign n7519 = t & n7518;
  assign n7520 = ~d0 & n7519;
  assign n7521 = ~d & n7520;
  assign n7522 = ~a0 & n7455;
  assign n7523 = ~c0 & n7522;
  assign n7524 = ~e0 & n7523;
  assign n7525 = ~j0 & n7524;
  assign n7526 = m0 & n7525;
  assign n7527 = ~i & n7526;
  assign n7528 = t & n7527;
  assign n7529 = ~d0 & n7528;
  assign n7530 = ~d & n7529;
  assign n7531 = ~g0 & n7514;
  assign n7532 = ~j0 & n7531;
  assign n7533 = m0 & n7532;
  assign n7534 = ~h0 & n7533;
  assign n7535 = t & n7534;
  assign n7536 = ~d0 & n7535;
  assign n7537 = ~d & n7536;
  assign n7538 = ~g0 & n7524;
  assign n7539 = ~j0 & n7538;
  assign n7540 = m0 & n7539;
  assign n7541 = t & n7540;
  assign n7542 = ~d0 & n7541;
  assign n7543 = ~d & n7542;
  assign n7544 = ~a0 & n7480;
  assign n7545 = ~c0 & n7544;
  assign n7546 = ~e0 & n7545;
  assign n7547 = ~j0 & n7546;
  assign n7548 = m0 & n7547;
  assign n7549 = ~h0 & n7548;
  assign n7550 = ~i & n7549;
  assign n7551 = ~d0 & n7550;
  assign n7552 = ~d & n7551;
  assign n7553 = ~a0 & n7490;
  assign n7554 = ~c0 & n7553;
  assign n7555 = ~e0 & n7554;
  assign n7556 = ~j0 & n7555;
  assign n7557 = m0 & n7556;
  assign n7558 = ~i & n7557;
  assign n7559 = ~d0 & n7558;
  assign n7560 = ~d & n7559;
  assign n7561 = ~g0 & n7546;
  assign n7562 = ~j0 & n7561;
  assign n7563 = m0 & n7562;
  assign n7564 = ~h0 & n7563;
  assign n7565 = ~d0 & n7564;
  assign n7566 = ~d & n7565;
  assign n7567 = ~g0 & n7555;
  assign n7568 = ~j0 & n7567;
  assign n7569 = m0 & n7568;
  assign n7570 = ~d0 & n7569;
  assign n7571 = ~d & n7570;
  assign n7572 = ~b & n7313;
  assign n7573 = ~b & n7325;
  assign n7574 = ~b & n7336;
  assign n7575 = ~b & n7346;
  assign n7576 = ~b & n7356;
  assign n7577 = ~b & n7365;
  assign n7578 = ~b & n7374;
  assign n7579 = ~b & n7382;
  assign n7580 = ~b & n7391;
  assign n7581 = ~b & n7399;
  assign n7582 = ~b & n7407;
  assign n7583 = ~b & n7414;
  assign n7584 = ~b & n7422;
  assign n7585 = ~b & n7429;
  assign n7586 = ~b & n7436;
  assign n7587 = ~b & n7442;
  assign n7588 = ~y & n7026;
  assign n7589 = ~c0 & n7588;
  assign n7590 = ~e0 & n7589;
  assign n7591 = ~j0 & n7590;
  assign n7592 = m0 & n7591;
  assign n7593 = ~h0 & n7592;
  assign n7594 = ~i & n7593;
  assign n7595 = t & n7594;
  assign n7596 = ~d0 & n7595;
  assign n7597 = i0 & n7596;
  assign n7598 = ~z & n7588;
  assign n7599 = ~c0 & n7598;
  assign n7600 = ~e0 & n7599;
  assign n7601 = ~j0 & n7600;
  assign n7602 = m0 & n7601;
  assign n7603 = ~i & n7602;
  assign n7604 = t & n7603;
  assign n7605 = ~d0 & n7604;
  assign n7606 = i0 & n7605;
  assign n7607 = ~g0 & n7590;
  assign n7608 = ~j0 & n7607;
  assign n7609 = m0 & n7608;
  assign n7610 = ~h0 & n7609;
  assign n7611 = t & n7610;
  assign n7612 = ~d0 & n7611;
  assign n7613 = i0 & n7612;
  assign n7614 = ~g0 & n7600;
  assign n7615 = ~j0 & n7614;
  assign n7616 = m0 & n7615;
  assign n7617 = t & n7616;
  assign n7618 = ~d0 & n7617;
  assign n7619 = i0 & n7618;
  assign n7620 = ~y & n7058;
  assign n7621 = ~c0 & n7620;
  assign n7622 = ~e0 & n7621;
  assign n7623 = ~j0 & n7622;
  assign n7624 = m0 & n7623;
  assign n7625 = ~h0 & n7624;
  assign n7626 = ~i & n7625;
  assign n7627 = ~d0 & n7626;
  assign n7628 = i0 & n7627;
  assign n7629 = ~z & n7620;
  assign n7630 = ~c0 & n7629;
  assign n7631 = ~e0 & n7630;
  assign n7632 = ~j0 & n7631;
  assign n7633 = m0 & n7632;
  assign n7634 = ~i & n7633;
  assign n7635 = ~d0 & n7634;
  assign n7636 = i0 & n7635;
  assign n7637 = ~g0 & n7622;
  assign n7638 = ~j0 & n7637;
  assign n7639 = m0 & n7638;
  assign n7640 = ~h0 & n7639;
  assign n7641 = ~d0 & n7640;
  assign n7642 = i0 & n7641;
  assign n7643 = ~g0 & n7631;
  assign n7644 = ~j0 & n7643;
  assign n7645 = m0 & n7644;
  assign n7646 = ~d0 & n7645;
  assign n7647 = i0 & n7646;
  assign n7648 = ~a0 & n7588;
  assign n7649 = ~c0 & n7648;
  assign n7650 = ~e0 & n7649;
  assign n7651 = ~j0 & n7650;
  assign n7652 = m0 & n7651;
  assign n7653 = ~h0 & n7652;
  assign n7654 = ~i & n7653;
  assign n7655 = t & n7654;
  assign n7656 = ~d0 & n7655;
  assign n7657 = ~a0 & n7598;
  assign n7658 = ~c0 & n7657;
  assign n7659 = ~e0 & n7658;
  assign n7660 = ~j0 & n7659;
  assign n7661 = m0 & n7660;
  assign n7662 = ~i & n7661;
  assign n7663 = t & n7662;
  assign n7664 = ~d0 & n7663;
  assign n7665 = ~g0 & n7650;
  assign n7666 = ~j0 & n7665;
  assign n7667 = m0 & n7666;
  assign n7668 = ~h0 & n7667;
  assign n7669 = t & n7668;
  assign n7670 = ~d0 & n7669;
  assign n7671 = ~g0 & n7659;
  assign n7672 = ~j0 & n7671;
  assign n7673 = m0 & n7672;
  assign n7674 = t & n7673;
  assign n7675 = ~d0 & n7674;
  assign n7676 = ~a0 & n7620;
  assign n7677 = ~c0 & n7676;
  assign n7678 = ~e0 & n7677;
  assign n7679 = ~j0 & n7678;
  assign n7680 = m0 & n7679;
  assign n7681 = ~h0 & n7680;
  assign n7682 = ~i & n7681;
  assign n7683 = ~d0 & n7682;
  assign n7684 = ~a0 & n7629;
  assign n7685 = ~c0 & n7684;
  assign n7686 = ~e0 & n7685;
  assign n7687 = ~j0 & n7686;
  assign n7688 = m0 & n7687;
  assign n7689 = ~i & n7688;
  assign n7690 = ~d0 & n7689;
  assign n7691 = ~g0 & n7678;
  assign n7692 = ~j0 & n7691;
  assign n7693 = m0 & n7692;
  assign n7694 = ~h0 & n7693;
  assign n7695 = ~d0 & n7694;
  assign n7696 = ~g0 & n7686;
  assign n7697 = ~j0 & n7696;
  assign n7698 = m0 & n7697;
  assign n7699 = ~d0 & n7698;
  assign n7700 = j & ~w;
  assign n7701 = ~y & n7700;
  assign n7702 = ~a0 & n7701;
  assign n7703 = ~c0 & n7702;
  assign n7704 = ~e0 & n7703;
  assign n7705 = ~j0 & n7704;
  assign n7706 = m0 & n7705;
  assign n7707 = ~h0 & n7706;
  assign n7708 = ~i & n7707;
  assign n7709 = m & n7708;
  assign n7710 = ~k & n7709;
  assign n7711 = ~z & n7701;
  assign n7712 = ~a0 & n7711;
  assign n7713 = ~c0 & n7712;
  assign n7714 = ~e0 & n7713;
  assign n7715 = ~j0 & n7714;
  assign n7716 = m0 & n7715;
  assign n7717 = ~i & n7716;
  assign n7718 = m & n7717;
  assign n7719 = ~k & n7718;
  assign n7720 = ~g0 & n7704;
  assign n7721 = ~j0 & n7720;
  assign n7722 = m0 & n7721;
  assign n7723 = ~h0 & n7722;
  assign n7724 = m & n7723;
  assign n7725 = ~k & n7724;
  assign n7726 = ~g0 & n7714;
  assign n7727 = ~j0 & n7726;
  assign n7728 = m0 & n7727;
  assign n7729 = m & n7728;
  assign n7730 = ~k & n7729;
  assign n7731 = ~e0 & n5841;
  assign n7732 = ~j0 & n7731;
  assign n7733 = m0 & n7732;
  assign n7734 = ~h0 & n7733;
  assign n7735 = ~i & n7734;
  assign n7736 = ~k & n7735;
  assign n7737 = ~e0 & n5853;
  assign n7738 = ~j0 & n7737;
  assign n7739 = m0 & n7738;
  assign n7740 = ~i & n7739;
  assign n7741 = ~k & n7740;
  assign n7742 = ~g0 & n7731;
  assign n7743 = ~j0 & n7742;
  assign n7744 = m0 & n7743;
  assign n7745 = ~h0 & n7744;
  assign n7746 = ~k & n7745;
  assign n7747 = ~g0 & n7737;
  assign n7748 = ~j0 & n7747;
  assign n7749 = m0 & n7748;
  assign n7750 = ~k & n7749;
  assign n7751 = ~f0 & n7706;
  assign n7752 = ~h0 & n7751;
  assign n7753 = ~i & n7752;
  assign n7754 = m & n7753;
  assign n7755 = ~f0 & n7716;
  assign n7756 = ~i & n7755;
  assign n7757 = m & n7756;
  assign n7758 = ~f0 & n7722;
  assign n7759 = ~h0 & n7758;
  assign n7760 = m & n7759;
  assign n7761 = ~f0 & n7728;
  assign n7762 = m & n7761;
  assign n7763 = j & ~y;
  assign n7764 = ~c0 & n7763;
  assign n7765 = ~e0 & n7764;
  assign n7766 = ~j0 & n7765;
  assign n7767 = m0 & n7766;
  assign n7768 = ~h0 & n7767;
  assign n7769 = ~i & n7768;
  assign n7770 = ~d0 & n7769;
  assign n7771 = i0 & n7770;
  assign n7772 = ~k & n7771;
  assign n7773 = ~z & n7763;
  assign n7774 = ~c0 & n7773;
  assign n7775 = ~e0 & n7774;
  assign n7776 = ~j0 & n7775;
  assign n7777 = m0 & n7776;
  assign n7778 = ~i & n7777;
  assign n7779 = ~d0 & n7778;
  assign n7780 = i0 & n7779;
  assign n7781 = ~k & n7780;
  assign n7782 = ~g0 & n7765;
  assign n7783 = ~j0 & n7782;
  assign n7784 = m0 & n7783;
  assign n7785 = ~h0 & n7784;
  assign n7786 = ~d0 & n7785;
  assign n7787 = i0 & n7786;
  assign n7788 = ~k & n7787;
  assign n7789 = ~g0 & n7775;
  assign n7790 = ~j0 & n7789;
  assign n7791 = m0 & n7790;
  assign n7792 = ~d0 & n7791;
  assign n7793 = i0 & n7792;
  assign n7794 = ~k & n7793;
  assign n7795 = ~a0 & n7763;
  assign n7796 = ~c0 & n7795;
  assign n7797 = ~e0 & n7796;
  assign n7798 = ~j0 & n7797;
  assign n7799 = m0 & n7798;
  assign n7800 = ~h0 & n7799;
  assign n7801 = ~i & n7800;
  assign n7802 = ~d0 & n7801;
  assign n7803 = ~k & n7802;
  assign n7804 = ~a0 & n7773;
  assign n7805 = ~c0 & n7804;
  assign n7806 = ~e0 & n7805;
  assign n7807 = ~j0 & n7806;
  assign n7808 = m0 & n7807;
  assign n7809 = ~i & n7808;
  assign n7810 = ~d0 & n7809;
  assign n7811 = ~k & n7810;
  assign n7812 = ~g0 & n7797;
  assign n7813 = ~j0 & n7812;
  assign n7814 = m0 & n7813;
  assign n7815 = ~h0 & n7814;
  assign n7816 = ~d0 & n7815;
  assign n7817 = ~k & n7816;
  assign n7818 = ~g0 & n7806;
  assign n7819 = ~j0 & n7818;
  assign n7820 = m0 & n7819;
  assign n7821 = ~d0 & n7820;
  assign n7822 = ~k & n7821;
  assign n7823 = m0 & n7704;
  assign n7824 = ~h0 & n7823;
  assign n7825 = ~h & n7824;
  assign n7826 = ~i & n7825;
  assign n7827 = m & n7826;
  assign n7828 = m0 & n7714;
  assign n7829 = ~h & n7828;
  assign n7830 = ~i & n7829;
  assign n7831 = m & n7830;
  assign n7832 = m0 & n7720;
  assign n7833 = ~h0 & n7832;
  assign n7834 = ~h & n7833;
  assign n7835 = m & n7834;
  assign n7836 = m0 & n7726;
  assign n7837 = ~h & n7836;
  assign n7838 = m & n7837;
  assign n7839 = ~e0 & n6919;
  assign n7840 = ~j0 & n7839;
  assign n7841 = m0 & n7840;
  assign n7842 = ~f0 & n7841;
  assign n7843 = ~h0 & n7842;
  assign n7844 = ~i & n7843;
  assign n7845 = ~e0 & n6931;
  assign n7846 = ~j0 & n7845;
  assign n7847 = m0 & n7846;
  assign n7848 = ~f0 & n7847;
  assign n7849 = ~i & n7848;
  assign n7850 = ~g0 & n7839;
  assign n7851 = ~j0 & n7850;
  assign n7852 = m0 & n7851;
  assign n7853 = ~f0 & n7852;
  assign n7854 = ~h0 & n7853;
  assign n7855 = ~g0 & n7845;
  assign n7856 = ~j0 & n7855;
  assign n7857 = m0 & n7856;
  assign n7858 = ~f0 & n7857;
  assign n7859 = ~y & ~c0;
  assign n7860 = ~e0 & n7859;
  assign n7861 = ~j0 & n7860;
  assign n7862 = m0 & n7861;
  assign n7863 = ~f0 & n7862;
  assign n7864 = ~h0 & n7863;
  assign n7865 = ~i & n7864;
  assign n7866 = ~d0 & n7865;
  assign n7867 = i0 & n7866;
  assign n7868 = ~y & ~z;
  assign n7869 = ~c0 & n7868;
  assign n7870 = ~e0 & n7869;
  assign n7871 = ~j0 & n7870;
  assign n7872 = m0 & n7871;
  assign n7873 = ~f0 & n7872;
  assign n7874 = ~i & n7873;
  assign n7875 = ~d0 & n7874;
  assign n7876 = i0 & n7875;
  assign n7877 = ~g0 & n7860;
  assign n7878 = ~j0 & n7877;
  assign n7879 = m0 & n7878;
  assign n7880 = ~f0 & n7879;
  assign n7881 = ~h0 & n7880;
  assign n7882 = ~d0 & n7881;
  assign n7883 = i0 & n7882;
  assign n7884 = ~g0 & n7870;
  assign n7885 = ~j0 & n7884;
  assign n7886 = m0 & n7885;
  assign n7887 = ~f0 & n7886;
  assign n7888 = ~d0 & n7887;
  assign n7889 = i0 & n7888;
  assign n7890 = ~e0 & n4346;
  assign n7891 = ~j0 & n7890;
  assign n7892 = m0 & n7891;
  assign n7893 = ~f0 & n7892;
  assign n7894 = ~h0 & n7893;
  assign n7895 = ~i & n7894;
  assign n7896 = ~d0 & n7895;
  assign n7897 = ~a0 & n7868;
  assign n7898 = ~c0 & n7897;
  assign n7899 = ~e0 & n7898;
  assign n7900 = ~j0 & n7899;
  assign n7901 = m0 & n7900;
  assign n7902 = ~f0 & n7901;
  assign n7903 = ~i & n7902;
  assign n7904 = ~d0 & n7903;
  assign n7905 = ~g0 & n7890;
  assign n7906 = ~j0 & n7905;
  assign n7907 = m0 & n7906;
  assign n7908 = ~f0 & n7907;
  assign n7909 = ~h0 & n7908;
  assign n7910 = ~d0 & n7909;
  assign n7911 = ~g0 & n7899;
  assign n7912 = ~j0 & n7911;
  assign n7913 = m0 & n7912;
  assign n7914 = ~f0 & n7913;
  assign n7915 = ~d0 & n7914;
  assign n7916 = m0 & n7839;
  assign n7917 = ~h0 & n7916;
  assign n7918 = ~h & n7917;
  assign n7919 = ~i & n7918;
  assign n7920 = m0 & n7845;
  assign n7921 = ~h & n7920;
  assign n7922 = ~i & n7921;
  assign n7923 = m0 & n7850;
  assign n7924 = ~h0 & n7923;
  assign n7925 = ~h & n7924;
  assign n7926 = m0 & n7855;
  assign n7927 = ~h & n7926;
  assign n7928 = ~c0 & ~e0;
  assign n7929 = j0 & n7928;
  assign n7930 = m0 & n7929;
  assign n7931 = ~h0 & n7930;
  assign n7932 = ~h & n7931;
  assign n7933 = ~i & n7932;
  assign n7934 = ~d0 & n7933;
  assign n7935 = ~i0 & n7934;
  assign n7936 = ~z & ~c0;
  assign n7937 = ~e0 & n7936;
  assign n7938 = j0 & n7937;
  assign n7939 = m0 & n7938;
  assign n7940 = ~h & n7939;
  assign n7941 = ~i & n7940;
  assign n7942 = ~d0 & n7941;
  assign n7943 = ~i0 & n7942;
  assign n7944 = ~g0 & n7928;
  assign n7945 = j0 & n7944;
  assign n7946 = m0 & n7945;
  assign n7947 = ~h0 & n7946;
  assign n7948 = ~h & n7947;
  assign n7949 = ~d0 & n7948;
  assign n7950 = ~i0 & n7949;
  assign n7951 = ~g0 & n7937;
  assign n7952 = j0 & n7951;
  assign n7953 = m0 & n7952;
  assign n7954 = ~h & n7953;
  assign n7955 = ~d0 & n7954;
  assign n7956 = ~i0 & n7955;
  assign n7957 = m0 & n7860;
  assign n7958 = ~h0 & n7957;
  assign n7959 = ~h & n7958;
  assign n7960 = ~i & n7959;
  assign n7961 = ~d0 & n7960;
  assign n7962 = i0 & n7961;
  assign n7963 = m0 & n7870;
  assign n7964 = ~h & n7963;
  assign n7965 = ~i & n7964;
  assign n7966 = ~d0 & n7965;
  assign n7967 = i0 & n7966;
  assign n7968 = m0 & n7877;
  assign n7969 = ~h0 & n7968;
  assign n7970 = ~h & n7969;
  assign n7971 = ~d0 & n7970;
  assign n7972 = i0 & n7971;
  assign n7973 = m0 & n7884;
  assign n7974 = ~h & n7973;
  assign n7975 = ~d0 & n7974;
  assign n7976 = i0 & n7975;
  assign n7977 = m0 & n7890;
  assign n7978 = ~h0 & n7977;
  assign n7979 = ~h & n7978;
  assign n7980 = ~i & n7979;
  assign n7981 = ~d0 & n7980;
  assign n7982 = m0 & n7899;
  assign n7983 = ~h & n7982;
  assign n7984 = ~i & n7983;
  assign n7985 = ~d0 & n7984;
  assign n7986 = m0 & n7905;
  assign n7987 = ~h0 & n7986;
  assign n7988 = ~h & n7987;
  assign n7989 = ~d0 & n7988;
  assign n7990 = m0 & n7911;
  assign n7991 = ~h & n7990;
  assign n7992 = ~d0 & n7991;
  assign n7993 = j0 & ~c0;
  assign n7994 = f0 & n7993;
  assign n7995 = ~d0 & n7994;
  assign n7996 = ~i0 & n7995;
  assign n7997 = m & n7996;
  assign n7998 = r & n7997;
  assign n7999 = g0 & ~c0;
  assign n8000 = j0 & n7999;
  assign n8001 = ~d0 & n8000;
  assign n8002 = ~i0 & n8001;
  assign n8003 = m & n8002;
  assign n8004 = r & n8003;
  assign n8005 = ~c0 & e0;
  assign n8006 = j0 & n8005;
  assign n8007 = ~d0 & n8006;
  assign n8008 = ~i0 & n8007;
  assign n8009 = m & n8008;
  assign n8010 = r & n8009;
  assign n8011 = j0 & n102;
  assign n8012 = f0 & n8011;
  assign n8013 = ~i0 & n8012;
  assign n8014 = m & n8013;
  assign n8015 = r & n8014;
  assign n8016 = g0 & n102;
  assign n8017 = j0 & n8016;
  assign n8018 = ~i0 & n8017;
  assign n8019 = m & n8018;
  assign n8020 = r & n8019;
  assign n8021 = e0 & n102;
  assign n8022 = j0 & n8021;
  assign n8023 = ~i0 & n8022;
  assign n8024 = m & n8023;
  assign n8025 = r & n8024;
  assign n8026 = f0 & n7859;
  assign n8027 = ~d0 & n8026;
  assign n8028 = i0 & n8027;
  assign n8029 = m & n8028;
  assign n8030 = r & n8029;
  assign n8031 = g0 & n7859;
  assign n8032 = ~d0 & n8031;
  assign n8033 = i0 & n8032;
  assign n8034 = m & n8033;
  assign n8035 = r & n8034;
  assign n8036 = e0 & n7859;
  assign n8037 = ~d0 & n8036;
  assign n8038 = i0 & n8037;
  assign n8039 = m & n8038;
  assign n8040 = r & n8039;
  assign n8041 = ~c0 & n68;
  assign n8042 = f0 & n8041;
  assign n8043 = i0 & n8042;
  assign n8044 = m & n8043;
  assign n8045 = r & n8044;
  assign n8046 = g0 & n8041;
  assign n8047 = i0 & n8046;
  assign n8048 = m & n8047;
  assign n8049 = r & n8048;
  assign n8050 = e0 & n8041;
  assign n8051 = i0 & n8050;
  assign n8052 = m & n8051;
  assign n8053 = r & n8052;
  assign n8054 = ~w & ~y;
  assign n8055 = ~a0 & n8054;
  assign n8056 = ~c0 & n8055;
  assign n8057 = d0 & n8056;
  assign n8058 = m & n8057;
  assign n8059 = r & n8058;
  assign n8060 = n & ~c0;
  assign n8061 = j0 & n8060;
  assign n8062 = f0 & n8061;
  assign n8063 = o & n8062;
  assign n8064 = ~d0 & n8063;
  assign n8065 = ~i0 & n8064;
  assign n8066 = g0 & n8060;
  assign n8067 = j0 & n8066;
  assign n8068 = o & n8067;
  assign n8069 = ~d0 & n8068;
  assign n8070 = ~i0 & n8069;
  assign n8071 = e0 & n8060;
  assign n8072 = j0 & n8071;
  assign n8073 = o & n8072;
  assign n8074 = ~d0 & n8073;
  assign n8075 = ~i0 & n8074;
  assign n8076 = n & w;
  assign n8077 = ~c0 & n8076;
  assign n8078 = j0 & n8077;
  assign n8079 = f0 & n8078;
  assign n8080 = o & n8079;
  assign n8081 = ~i0 & n8080;
  assign n8082 = g0 & n8077;
  assign n8083 = j0 & n8082;
  assign n8084 = o & n8083;
  assign n8085 = ~i0 & n8084;
  assign n8086 = e0 & n8077;
  assign n8087 = j0 & n8086;
  assign n8088 = o & n8087;
  assign n8089 = ~i0 & n8088;
  assign n8090 = n & ~y;
  assign n8091 = ~c0 & n8090;
  assign n8092 = f0 & n8091;
  assign n8093 = o & n8092;
  assign n8094 = ~d0 & n8093;
  assign n8095 = i0 & n8094;
  assign n8096 = g0 & n8091;
  assign n8097 = o & n8096;
  assign n8098 = ~d0 & n8097;
  assign n8099 = i0 & n8098;
  assign n8100 = e0 & n8091;
  assign n8101 = o & n8100;
  assign n8102 = ~d0 & n8101;
  assign n8103 = i0 & n8102;
  assign n8104 = ~y & n8076;
  assign n8105 = ~c0 & n8104;
  assign n8106 = f0 & n8105;
  assign n8107 = o & n8106;
  assign n8108 = i0 & n8107;
  assign n8109 = g0 & n8105;
  assign n8110 = o & n8109;
  assign n8111 = i0 & n8110;
  assign n8112 = e0 & n8105;
  assign n8113 = o & n8112;
  assign n8114 = i0 & n8113;
  assign n8115 = n & ~w;
  assign n8116 = ~y & n8115;
  assign n8117 = ~a0 & n8116;
  assign n8118 = ~c0 & n8117;
  assign n8119 = o & n8118;
  assign n8120 = d0 & n8119;
  assign n8121 = ~w & ~c0;
  assign n8122 = j0 & n8121;
  assign n8123 = d0 & n8122;
  assign n8124 = ~i0 & n8123;
  assign n8125 = v & n8124;
  assign n8126 = ~c0 & n8054;
  assign n8127 = d0 & n8126;
  assign n8128 = i0 & n8127;
  assign n8129 = v & n8128;
  assign n8130 = u & n8124;
  assign n8131 = u & n8128;
  assign n8132 = f0 & n4346;
  assign n8133 = m & n8132;
  assign n8134 = r & n8133;
  assign n8135 = g0 & n4346;
  assign n8136 = m & n8135;
  assign n8137 = r & n8136;
  assign n8138 = e0 & n4346;
  assign n8139 = m & n8138;
  assign n8140 = r & n8139;
  assign n8141 = b0 & n7996;
  assign n8142 = b0 & n8002;
  assign n8143 = b0 & n8008;
  assign n8144 = b0 & n8013;
  assign n8145 = b0 & n8018;
  assign n8146 = b0 & n8023;
  assign n8147 = b0 & n8028;
  assign n8148 = b0 & n8033;
  assign n8149 = b0 & n8038;
  assign n8150 = b0 & n8043;
  assign n8151 = b0 & n8047;
  assign n8152 = b0 & n8051;
  assign n8153 = b0 & n8057;
  assign n8154 = q & n7996;
  assign n8155 = q & n8002;
  assign n8156 = q & n8008;
  assign n8157 = q & n8013;
  assign n8158 = q & n8018;
  assign n8159 = q & n8023;
  assign n8160 = q & n8028;
  assign n8161 = q & n8033;
  assign n8162 = q & n8038;
  assign n8163 = q & n8043;
  assign n8164 = q & n8047;
  assign n8165 = q & n8051;
  assign n8166 = q & n8057;
  assign n8167 = x & n7993;
  assign n8168 = f0 & n8167;
  assign n8169 = ~d0 & n8168;
  assign n8170 = ~i0 & n8169;
  assign n8171 = x & n8000;
  assign n8172 = ~d0 & n8171;
  assign n8173 = ~i0 & n8172;
  assign n8174 = x & n8006;
  assign n8175 = ~d0 & n8174;
  assign n8176 = ~i0 & n8175;
  assign n8177 = o & n8011;
  assign n8178 = h0 & n8177;
  assign n8179 = ~i0 & n8178;
  assign n8180 = x & n8011;
  assign n8181 = f0 & n8180;
  assign n8182 = ~i0 & n8181;
  assign n8183 = x & n8017;
  assign n8184 = ~i0 & n8183;
  assign n8185 = x & n8022;
  assign n8186 = ~i0 & n8185;
  assign n8187 = o & n8041;
  assign n8188 = h0 & n8187;
  assign n8189 = i0 & n8188;
  assign n8190 = x & n8056;
  assign n8191 = d0 & n8190;
  assign n8192 = ~a0 & n8090;
  assign n8193 = ~c0 & n8192;
  assign n8194 = f0 & n8193;
  assign n8195 = o & n8194;
  assign n8196 = g0 & n8193;
  assign n8197 = o & n8196;
  assign n8198 = e0 & n8193;
  assign n8199 = o & n8198;
  assign n8200 = b0 & n8132;
  assign n8201 = b0 & n8135;
  assign n8202 = b0 & n8138;
  assign n8203 = q & n8132;
  assign n8204 = q & n8135;
  assign n8205 = q & n8138;
  assign n8206 = x & n7859;
  assign n8207 = ~d0 & n8206;
  assign n8208 = i0 & n8207;
  assign n8209 = x & n8041;
  assign n8210 = i0 & n8209;
  assign n8211 = o & n4346;
  assign n8212 = h0 & n8211;
  assign n8213 = x & n4346;
  assign n8214 = f0 & n8213;
  assign n8215 = x & n8135;
  assign n8216 = x & n8138;
  assign n8217 = ~n261 & ~n270;
  assign n8218 = ~n252 & n8217;
  assign n8219 = ~n243 & n8218;
  assign n8220 = ~n234 & n8219;
  assign n8221 = ~n228 & n8220;
  assign n8222 = ~n2536 & n8221;
  assign n8223 = ~n2528 & n8222;
  assign n8224 = ~n2520 & n8223;
  assign n8225 = ~n166 & n8224;
  assign n8226 = ~n158 & n8225;
  assign n8227 = ~n2512 & n8226;
  assign n8228 = ~n149 & n8227;
  assign n8229 = ~n124 & n8228;
  assign n8230 = ~n8216 & n8229;
  assign n8231 = ~n8215 & n8230;
  assign n8232 = ~n8214 & n8231;
  assign n8233 = ~n8212 & n8232;
  assign n8234 = ~n8210 & n8233;
  assign n8235 = ~n8208 & n8234;
  assign n8236 = ~n8205 & n8235;
  assign n8237 = ~n8204 & n8236;
  assign n8238 = ~n8203 & n8237;
  assign n8239 = ~n8202 & n8238;
  assign n8240 = ~n8201 & n8239;
  assign n8241 = ~n8200 & n8240;
  assign n8242 = ~n8199 & n8241;
  assign n8243 = ~n8197 & n8242;
  assign n8244 = ~n8195 & n8243;
  assign n8245 = ~n8191 & n8244;
  assign n8246 = ~n8189 & n8245;
  assign n8247 = ~n8186 & n8246;
  assign n8248 = ~n8184 & n8247;
  assign n8249 = ~n8182 & n8248;
  assign n8250 = ~n8179 & n8249;
  assign n8251 = ~n8176 & n8250;
  assign n8252 = ~n8173 & n8251;
  assign n8253 = ~n8170 & n8252;
  assign n8254 = ~n8166 & n8253;
  assign n8255 = ~n8165 & n8254;
  assign n8256 = ~n8164 & n8255;
  assign n8257 = ~n8163 & n8256;
  assign n8258 = ~n8162 & n8257;
  assign n8259 = ~n8161 & n8258;
  assign n8260 = ~n8160 & n8259;
  assign n8261 = ~n8159 & n8260;
  assign n8262 = ~n8158 & n8261;
  assign n8263 = ~n8157 & n8262;
  assign n8264 = ~n8156 & n8263;
  assign n8265 = ~n8155 & n8264;
  assign n8266 = ~n8154 & n8265;
  assign n8267 = ~n8153 & n8266;
  assign n8268 = ~n8152 & n8267;
  assign n8269 = ~n8151 & n8268;
  assign n8270 = ~n8150 & n8269;
  assign n8271 = ~n8149 & n8270;
  assign n8272 = ~n8148 & n8271;
  assign n8273 = ~n8147 & n8272;
  assign n8274 = ~n8146 & n8273;
  assign n8275 = ~n8145 & n8274;
  assign n8276 = ~n8144 & n8275;
  assign n8277 = ~n8143 & n8276;
  assign n8278 = ~n8142 & n8277;
  assign n8279 = ~n8141 & n8278;
  assign n8280 = ~n8140 & n8279;
  assign n8281 = ~n8137 & n8280;
  assign n8282 = ~n8134 & n8281;
  assign n8283 = ~n8131 & n8282;
  assign n8284 = ~n8130 & n8283;
  assign n8285 = ~n8129 & n8284;
  assign n8286 = ~n8125 & n8285;
  assign n8287 = ~n8120 & n8286;
  assign n8288 = ~n8114 & n8287;
  assign n8289 = ~n8111 & n8288;
  assign n8290 = ~n8108 & n8289;
  assign n8291 = ~n8103 & n8290;
  assign n8292 = ~n8099 & n8291;
  assign n8293 = ~n8095 & n8292;
  assign n8294 = ~n8089 & n8293;
  assign n8295 = ~n8085 & n8294;
  assign n8296 = ~n8081 & n8295;
  assign n8297 = ~n8075 & n8296;
  assign n8298 = ~n8070 & n8297;
  assign n8299 = ~n8065 & n8298;
  assign n8300 = ~n8059 & n8299;
  assign n8301 = ~n8053 & n8300;
  assign n8302 = ~n8049 & n8301;
  assign n8303 = ~n8045 & n8302;
  assign n8304 = ~n8040 & n8303;
  assign n8305 = ~n8035 & n8304;
  assign n8306 = ~n8030 & n8305;
  assign n8307 = ~n8025 & n8306;
  assign n8308 = ~n8020 & n8307;
  assign n8309 = ~n8015 & n8308;
  assign n8310 = ~n8010 & n8309;
  assign n8311 = ~n8004 & n8310;
  assign n8312 = ~n7998 & n8311;
  assign n8313 = ~n7992 & n8312;
  assign n8314 = ~n7989 & n8313;
  assign n8315 = ~n7985 & n8314;
  assign n8316 = ~n7981 & n8315;
  assign n8317 = ~n7976 & n8316;
  assign n8318 = ~n7972 & n8317;
  assign n8319 = ~n7967 & n8318;
  assign n8320 = ~n7962 & n8319;
  assign n8321 = ~n7956 & n8320;
  assign n8322 = ~n7950 & n8321;
  assign n8323 = ~n7943 & n8322;
  assign n8324 = ~n7935 & n8323;
  assign n8325 = ~n7927 & n8324;
  assign n8326 = ~n7925 & n8325;
  assign n8327 = ~n7922 & n8326;
  assign n8328 = ~n7919 & n8327;
  assign n8329 = ~n7915 & n8328;
  assign n8330 = ~n7910 & n8329;
  assign n8331 = ~n7904 & n8330;
  assign n8332 = ~n7896 & n8331;
  assign n8333 = ~n7889 & n8332;
  assign n8334 = ~n7883 & n8333;
  assign n8335 = ~n7876 & n8334;
  assign n8336 = ~n7867 & n8335;
  assign n8337 = ~n7858 & n8336;
  assign n8338 = ~n7854 & n8337;
  assign n8339 = ~n7849 & n8338;
  assign n8340 = ~n7844 & n8339;
  assign n8341 = ~n7838 & n8340;
  assign n8342 = ~n7835 & n8341;
  assign n8343 = ~n7831 & n8342;
  assign n8344 = ~n7827 & n8343;
  assign n8345 = ~n7822 & n8344;
  assign n8346 = ~n7817 & n8345;
  assign n8347 = ~n7811 & n8346;
  assign n8348 = ~n7803 & n8347;
  assign n8349 = ~n7794 & n8348;
  assign n8350 = ~n7788 & n8349;
  assign n8351 = ~n7781 & n8350;
  assign n8352 = ~n7772 & n8351;
  assign n8353 = ~n7762 & n8352;
  assign n8354 = ~n7760 & n8353;
  assign n8355 = ~n7757 & n8354;
  assign n8356 = ~n7754 & n8355;
  assign n8357 = ~n7750 & n8356;
  assign n8358 = ~n7746 & n8357;
  assign n8359 = ~n7741 & n8358;
  assign n8360 = ~n7736 & n8359;
  assign n8361 = ~n7730 & n8360;
  assign n8362 = ~n7725 & n8361;
  assign n8363 = ~n7719 & n8362;
  assign n8364 = ~n7710 & n8363;
  assign n8365 = ~n7699 & n8364;
  assign n8366 = ~n7695 & n8365;
  assign n8367 = ~n7690 & n8366;
  assign n8368 = ~n7683 & n8367;
  assign n8369 = ~n7675 & n8368;
  assign n8370 = ~n7670 & n8369;
  assign n8371 = ~n7664 & n8370;
  assign n8372 = ~n7656 & n8371;
  assign n8373 = ~n7647 & n8372;
  assign n8374 = ~n7642 & n8373;
  assign n8375 = ~n7636 & n8374;
  assign n8376 = ~n7628 & n8375;
  assign n8377 = ~n7619 & n8376;
  assign n8378 = ~n7613 & n8377;
  assign n8379 = ~n7606 & n8378;
  assign n8380 = ~n7597 & n8379;
  assign n8381 = ~n7587 & n8380;
  assign n8382 = ~n7586 & n8381;
  assign n8383 = ~n7585 & n8382;
  assign n8384 = ~n7584 & n8383;
  assign n8385 = ~n7583 & n8384;
  assign n8386 = ~n7582 & n8385;
  assign n8387 = ~n7581 & n8386;
  assign n8388 = ~n7580 & n8387;
  assign n8389 = ~n7579 & n8388;
  assign n8390 = ~n7578 & n8389;
  assign n8391 = ~n7577 & n8390;
  assign n8392 = ~n7576 & n8391;
  assign n8393 = ~n7575 & n8392;
  assign n8394 = ~n7574 & n8393;
  assign n8395 = ~n7573 & n8394;
  assign n8396 = ~n7572 & n8395;
  assign n8397 = ~n7571 & n8396;
  assign n8398 = ~n7566 & n8397;
  assign n8399 = ~n7560 & n8398;
  assign n8400 = ~n7552 & n8399;
  assign n8401 = ~n7543 & n8400;
  assign n8402 = ~n7537 & n8401;
  assign n8403 = ~n7530 & n8402;
  assign n8404 = ~n7521 & n8403;
  assign n8405 = ~n7511 & n8404;
  assign n8406 = ~n7505 & n8405;
  assign n8407 = ~n7498 & n8406;
  assign n8408 = ~n7489 & n8407;
  assign n8409 = ~n7479 & n8408;
  assign n8410 = ~n7472 & n8409;
  assign n8411 = ~n7464 & n8410;
  assign n8412 = ~n7454 & n8411;
  assign n8413 = ~n7443 & n8412;
  assign n8414 = ~n7437 & n8413;
  assign n8415 = ~n7430 & n8414;
  assign n8416 = ~n7423 & n8415;
  assign n8417 = ~n7415 & n8416;
  assign n8418 = ~n7408 & n8417;
  assign n8419 = ~n7400 & n8418;
  assign n8420 = ~n7392 & n8419;
  assign n8421 = ~n7383 & n8420;
  assign n8422 = ~n7375 & n8421;
  assign n8423 = ~n7366 & n8422;
  assign n8424 = ~n7357 & n8423;
  assign n8425 = ~n7347 & n8424;
  assign n8426 = ~n7337 & n8425;
  assign n8427 = ~n7326 & n8426;
  assign n8428 = ~n7314 & n8427;
  assign n8429 = ~n7302 & n8428;
  assign n8430 = ~n7299 & n8429;
  assign n8431 = ~n7295 & n8430;
  assign n8432 = ~n7290 & n8431;
  assign n8433 = ~n7284 & n8432;
  assign n8434 = ~n7280 & n8433;
  assign n8435 = ~n7275 & n8434;
  assign n8436 = ~n7269 & n8435;
  assign n8437 = ~n7262 & n8436;
  assign n8438 = ~n7258 & n8437;
  assign n8439 = ~n7253 & n8438;
  assign n8440 = ~n7248 & n8439;
  assign n8441 = ~n7242 & n8440;
  assign n8442 = ~n7236 & n8441;
  assign n8443 = ~n7229 & n8442;
  assign n8444 = ~n7222 & n8443;
  assign n8445 = ~n7214 & n8444;
  assign n8446 = ~n7207 & n8445;
  assign n8447 = ~n7199 & n8446;
  assign n8448 = ~n7191 & n8447;
  assign n8449 = ~n7182 & n8448;
  assign n8450 = ~n7173 & n8449;
  assign n8451 = ~n7163 & n8450;
  assign n8452 = ~n7152 & n8451;
  assign n8453 = ~n7141 & n8452;
  assign n8454 = ~n7140 & n8453;
  assign n8455 = ~n7139 & n8454;
  assign n8456 = ~n7138 & n8455;
  assign n8457 = ~n7137 & n8456;
  assign n8458 = ~n7136 & n8457;
  assign n8459 = ~n7135 & n8458;
  assign n8460 = ~n7134 & n8459;
  assign n8461 = ~n7133 & n8460;
  assign n8462 = ~n7132 & n8461;
  assign n8463 = ~n7131 & n8462;
  assign n8464 = ~n7130 & n8463;
  assign n8465 = ~n7129 & n8464;
  assign n8466 = ~n7125 & n8465;
  assign n8467 = ~n7120 & n8466;
  assign n8468 = ~n7115 & n8467;
  assign n8469 = ~n7109 & n8468;
  assign n8470 = ~n7104 & n8469;
  assign n8471 = ~n7098 & n8470;
  assign n8472 = ~n7092 & n8471;
  assign n8473 = ~n7085 & n8472;
  assign n8474 = ~n7081 & n8473;
  assign n8475 = ~n7076 & n8474;
  assign n8476 = ~n7068 & n8475;
  assign n8477 = ~n7057 & n8476;
  assign n8478 = ~n7052 & n8477;
  assign n8479 = ~n7046 & n8478;
  assign n8480 = ~n7037 & n8479;
  assign n8481 = ~n7025 & n8480;
  assign n8482 = ~n7020 & n8481;
  assign n8483 = ~n7014 & n8482;
  assign n8484 = ~n7005 & n8483;
  assign n8485 = ~n6992 & n8484;
  assign n8486 = ~n6986 & n8485;
  assign n8487 = ~n6979 & n8486;
  assign n8488 = ~n6969 & n8487;
  assign n8489 = ~n6956 & n8488;
  assign n8490 = ~n6948 & n8489;
  assign n8491 = ~n6939 & n8490;
  assign n8492 = ~n6928 & n8491;
  assign n8493 = ~n6915 & n8492;
  assign n8494 = ~n6906 & n8493;
  assign n8495 = ~n6896 & n8494;
  assign n8496 = ~n6885 & n8495;
  assign n8497 = ~n6873 & n8496;
  assign n8498 = ~n6863 & n8497;
  assign n8499 = ~n6852 & n8498;
  assign n8500 = ~n6840 & n8499;
  assign n8501 = ~n6827 & n8500;
  assign n8502 = ~n6823 & n8501;
  assign n8503 = ~n6818 & n8502;
  assign n8504 = ~n6813 & n8503;
  assign n8505 = ~n6807 & n8504;
  assign n8506 = ~n6802 & n8505;
  assign n8507 = ~n6796 & n8506;
  assign n8508 = ~n6790 & n8507;
  assign n8509 = ~n6783 & n8508;
  assign n8510 = ~n6778 & n8509;
  assign n8511 = ~n6772 & n8510;
  assign n8512 = ~n6766 & n8511;
  assign n8513 = ~n6759 & n8512;
  assign n8514 = ~n6753 & n8513;
  assign n8515 = ~n6746 & n8514;
  assign n8516 = ~n6739 & n8515;
  assign n8517 = ~n6731 & n8516;
  assign n8518 = ~n6725 & n8517;
  assign n8519 = ~n6718 & n8518;
  assign n8520 = ~n6711 & n8519;
  assign n8521 = ~n6703 & n8520;
  assign n8522 = ~n6696 & n8521;
  assign n8523 = ~n6688 & n8522;
  assign n8524 = ~n6680 & n8523;
  assign n8525 = ~n6671 & n8524;
  assign n8526 = ~n6663 & n8525;
  assign n8527 = ~n6654 & n8526;
  assign n8528 = ~n6645 & n8527;
  assign n8529 = ~n6635 & n8528;
  assign n8530 = ~n6625 & n8529;
  assign n8531 = ~n6614 & n8530;
  assign n8532 = ~n6602 & n8531;
  assign n8533 = ~n6590 & n8532;
  assign n8534 = ~n6583 & n8533;
  assign n8535 = ~n6575 & n8534;
  assign n8536 = ~n6565 & n8535;
  assign n8537 = ~n6553 & n8536;
  assign n8538 = ~n6547 & n8537;
  assign n8539 = ~n6540 & n8538;
  assign n8540 = ~n6533 & n8539;
  assign n8541 = ~n6525 & n8540;
  assign n8542 = ~n6517 & n8541;
  assign n8543 = ~n6508 & n8542;
  assign n8544 = ~n6498 & n8543;
  assign n8545 = ~n6487 & n8544;
  assign n8546 = ~n6480 & n8545;
  assign n8547 = ~n6472 & n8546;
  assign n8548 = ~n6464 & n8547;
  assign n8549 = ~n6455 & n8548;
  assign n8550 = ~n6446 & n8549;
  assign n8551 = ~n6436 & n8550;
  assign n8552 = ~n6425 & n8551;
  assign n8553 = ~n6412 & n8552;
  assign n8554 = ~n6404 & n8553;
  assign n8555 = ~n6395 & n8554;
  assign n8556 = ~n6386 & n8555;
  assign n8557 = ~n6376 & n8556;
  assign n8558 = ~n6366 & n8557;
  assign n8559 = ~n6355 & n8558;
  assign n8560 = ~n6343 & n8559;
  assign n8561 = ~n6331 & n8560;
  assign n8562 = ~n6325 & n8561;
  assign n8563 = ~n6318 & n8562;
  assign n8564 = ~n6311 & n8563;
  assign n8565 = ~n6303 & n8564;
  assign n8566 = ~n6296 & n8565;
  assign n8567 = ~n6288 & n8566;
  assign n8568 = ~n6280 & n8567;
  assign n8569 = ~n6271 & n8568;
  assign n8570 = ~n6263 & n8569;
  assign n8571 = ~n6254 & n8570;
  assign n8572 = ~n6245 & n8571;
  assign n8573 = ~n6235 & n8572;
  assign n8574 = ~n6225 & n8573;
  assign n8575 = ~n6214 & n8574;
  assign n8576 = ~n6202 & n8575;
  assign n8577 = ~n6190 & n8576;
  assign n8578 = ~n6184 & n8577;
  assign n8579 = ~n6177 & n8578;
  assign n8580 = ~n6167 & n8579;
  assign n8581 = ~n6154 & n8580;
  assign n8582 = ~n6147 & n8581;
  assign n8583 = ~n6139 & n8582;
  assign n8584 = ~n6128 & n8583;
  assign n8585 = ~n6114 & n8584;
  assign n8586 = ~n6107 & n8585;
  assign n8587 = ~n6099 & n8586;
  assign n8588 = ~n6088 & n8587;
  assign n8589 = ~n6074 & n8588;
  assign n8590 = ~n6066 & n8589;
  assign n8591 = ~n6057 & n8590;
  assign n8592 = ~n6045 & n8591;
  assign n8593 = ~n6031 & n8592;
  assign n8594 = ~n6023 & n8593;
  assign n8595 = ~n6014 & n8594;
  assign n8596 = ~n6003 & n8595;
  assign n8597 = ~n5990 & n8596;
  assign n8598 = ~n5981 & n8597;
  assign n8599 = ~n5971 & n8598;
  assign n8600 = ~n5960 & n8599;
  assign n8601 = ~n5948 & n8600;
  assign n8602 = ~n5938 & n8601;
  assign n8603 = ~n5927 & n8602;
  assign n8604 = ~n5915 & n8603;
  assign n8605 = ~n5902 & n8604;
  assign n8606 = ~n5900 & n8605;
  assign n8607 = ~n5898 & n8606;
  assign n8608 = ~n5896 & n8607;
  assign n8609 = ~n5894 & n8608;
  assign n8610 = ~n5892 & n8609;
  assign n8611 = ~n5890 & n8610;
  assign n8612 = ~n5888 & n8611;
  assign n8613 = ~n5886 & n8612;
  assign n8614 = ~n5884 & n8613;
  assign n8615 = ~n5882 & n8614;
  assign n8616 = ~n5880 & n8615;
  assign n8617 = ~n5878 & n8616;
  assign n8618 = ~n5870 & n8617;
  assign n8619 = ~n5861 & n8618;
  assign n8620 = ~n5850 & n8619;
  assign n8621 = ~n5837 & n8620;
  assign n8622 = ~n5828 & n8621;
  assign n8623 = ~n5818 & n8622;
  assign n8624 = ~n5807 & n8623;
  assign n8625 = ~n5795 & n8624;
  assign n8626 = ~n5785 & n8625;
  assign n8627 = ~n5774 & n8626;
  assign n8628 = ~n5762 & n8627;
  assign n8629 = ~n5749 & n8628;
  assign n8630 = ~n5741 & n8629;
  assign n8631 = ~n5732 & n8630;
  assign n8632 = ~n5721 & n8631;
  assign n8633 = ~n5708 & n8632;
  assign n8634 = ~n5699 & n8633;
  assign n8635 = ~n5689 & n8634;
  assign n8636 = ~n5678 & n8635;
  assign n8637 = ~n5666 & n8636;
  assign n8638 = ~n5656 & n8637;
  assign n8639 = ~n5645 & n8638;
  assign n8640 = ~n5633 & n8639;
  assign n8641 = ~n5619 & n8640;
  assign n8642 = ~n5611 & n8641;
  assign n8643 = ~n5602 & n8642;
  assign n8644 = ~n5591 & n8643;
  assign n8645 = ~n5578 & n8644;
  assign n8646 = ~n5569 & n8645;
  assign n8647 = ~n5559 & n8646;
  assign n8648 = ~n5548 & n8647;
  assign n8649 = ~n5536 & n8648;
  assign n8650 = ~n5526 & n8649;
  assign n8651 = ~n5515 & n8650;
  assign n8652 = ~n5503 & n8651;
  assign n8653 = ~n5488 & n8652;
  assign n8654 = ~n5487 & n8653;
  assign n8655 = ~n5486 & n8654;
  assign n8656 = ~n5485 & n8655;
  assign n8657 = ~n5484 & n8656;
  assign n8658 = ~n5483 & n8657;
  assign n8659 = ~n5482 & n8658;
  assign n8660 = ~n5481 & n8659;
  assign n8661 = ~n5480 & n8660;
  assign n8662 = ~n5479 & n8661;
  assign n8663 = ~n5478 & n8662;
  assign n8664 = ~n5477 & n8663;
  assign n8665 = ~n5476 & n8664;
  assign n8666 = ~n5475 & n8665;
  assign n8667 = ~n5474 & n8666;
  assign n8668 = ~n5473 & n8667;
  assign n8669 = ~n5472 & n8668;
  assign n8670 = ~n5471 & n8669;
  assign n8671 = ~n5470 & n8670;
  assign n8672 = ~n5469 & n8671;
  assign n8673 = ~n5468 & n8672;
  assign n8674 = ~n5467 & n8673;
  assign n8675 = ~n5466 & n8674;
  assign n8676 = ~n5465 & n8675;
  assign n8677 = ~n5464 & n8676;
  assign n8678 = ~n5462 & n8677;
  assign n8679 = ~n5460 & n8678;
  assign n8680 = ~n5458 & n8679;
  assign n8681 = ~n5456 & n8680;
  assign n8682 = ~n5454 & n8681;
  assign n8683 = ~n5452 & n8682;
  assign n8684 = ~n5450 & n8683;
  assign n8685 = ~n5448 & n8684;
  assign n8686 = ~n5446 & n8685;
  assign n8687 = ~n5444 & n8686;
  assign n8688 = ~n5442 & n8687;
  assign n8689 = ~n5440 & n8688;
  assign n8690 = ~n5438 & n8689;
  assign n8691 = ~n5436 & n8690;
  assign n8692 = ~n5434 & n8691;
  assign n8693 = ~n5432 & n8692;
  assign n8694 = ~n5430 & n8693;
  assign n8695 = ~n5428 & n8694;
  assign n8696 = ~n5426 & n8695;
  assign n8697 = ~n5424 & n8696;
  assign n8698 = ~n5422 & n8697;
  assign n8699 = ~n5420 & n8698;
  assign n8700 = ~n5418 & n8699;
  assign n8701 = ~n5416 & n8700;
  assign n8702 = ~n5409 & n8701;
  assign n8703 = ~n5401 & n8702;
  assign n8704 = ~n5391 & n8703;
  assign n8705 = ~n5379 & n8704;
  assign n8706 = ~n5371 & n8705;
  assign n8707 = ~n5362 & n8706;
  assign n8708 = ~n5351 & n8707;
  assign n8709 = ~n5338 & n8708;
  assign n8710 = ~n5330 & n8709;
  assign n8711 = ~n5321 & n8710;
  assign n8712 = ~n5311 & n8711;
  assign n8713 = ~n5300 & n8712;
  assign n8714 = ~n5291 & n8713;
  assign n8715 = ~n5281 & n8714;
  assign n8716 = ~n5270 & n8715;
  assign n8717 = ~n5258 & n8716;
  assign n8718 = ~n5249 & n8717;
  assign n8719 = ~n5239 & n8718;
  assign n8720 = ~n5228 & n8719;
  assign n8721 = ~n5215 & n8720;
  assign n8722 = ~n5205 & n8721;
  assign n8723 = ~n5194 & n8722;
  assign n8724 = ~n5182 & n8723;
  assign n8725 = ~n5168 & n8724;
  assign n8726 = ~n5160 & n8725;
  assign n8727 = ~n5151 & n8726;
  assign n8728 = ~n5140 & n8727;
  assign n8729 = ~n5127 & n8728;
  assign n8730 = ~n5118 & n8729;
  assign n8731 = ~n5108 & n8730;
  assign n8732 = ~n5096 & n8731;
  assign n8733 = ~n5082 & n8732;
  assign n8734 = ~n5073 & n8733;
  assign n8735 = ~n5063 & n8734;
  assign n8736 = ~n5052 & n8735;
  assign n8737 = ~n5040 & n8736;
  assign n8738 = ~n5030 & n8737;
  assign n8739 = ~n5019 & n8738;
  assign n8740 = ~n5007 & n8739;
  assign n8741 = ~n4994 & n8740;
  assign n8742 = ~n4984 & n8741;
  assign n8743 = ~n4973 & n8742;
  assign n8744 = ~n4961 & n8743;
  assign n8745 = ~n4946 & n8744;
  assign n8746 = ~n4935 & n8745;
  assign n8747 = ~n4923 & n8746;
  assign p0 = n4910 | ~n8747;
endmodule


