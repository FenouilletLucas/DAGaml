// Benchmark "i2" written by ABC on Tue May 16 16:07:50 2017

module i2 ( 
    \V126(17) , \V144(21) , \V30(29) , \V126(1) , \V126(16) , \V144(20) ,
    \V30(28) , \V126(0) , \V126(19) , \V144(23) , \V126(18) , \V144(22) ,
    \V62(13) , \V144(25) , \V62(12) , \V191(31) , \V144(24) , \V62(15) ,
    \V94(31) , \V62(14) , \V126(7) , \V94(30) , \V126(6) , \V144(19) ,
    \V30(31) , \V201(3) , \V126(9) , \V144(18) , \V62(11) , \V30(30) ,
    \V201(2) , \V126(8) , \V126(11) , \V62(10) , \V201(5) , \V126(10) ,
    \V201(4) , \V126(13) , \V176(31) , \V126(12) , \V176(30) , \V94(2) ,
    \V126(15) , \V63(0) , \V201(1) , \V94(3) , \V126(14) , \V62(17) ,
    \V201(0) , \V94(4) , \V193(1) , \V62(16) , \V94(5) , \V193(0) ,
    \V62(19) , \V94(6) , \V62(18) , \V176(3) , \V94(7) , \V62(23) ,
    \V176(2) , \V94(8) , \V129(0) , \V62(22) , \V176(5) , \V201(7) ,
    \V94(9) , \V62(25) , \V176(4) , \V201(6) , \V62(24) , \V176(27) ,
    \V176(26) , \V176(1) , \V176(29) , \V62(21) , \V176(0) , \V176(28) ,
    \V62(20) , \V188(31) , \V176(7) , \V62(0) , \V188(30) , \V62(27) ,
    \V176(6) , \V62(1) , \V62(26) , \V176(9) , \V176(21) , \V62(2) ,
    \V62(29) , \V176(8) , \V176(20) , \V62(3) , \V62(28) , \V176(23) ,
    \V62(4) , \V176(22) , \V62(5) , \V94(13) , \V128(0) , \V176(25) ,
    \V62(6) , \V94(12) , \V176(24) , \V62(7) , \V94(15) , \V30(13) ,
    \V130(0) , \V176(17) , \V62(8) , \V94(14) , \V30(12) , \V176(16) ,
    \V62(9) , \V188(27) , \V30(15) , \V176(19) , \V188(26) , \V62(31) ,
    \V30(14) , \V126(31) , \V176(18) , \V94(11) , \V188(29) , \V62(30) ,
    \V126(30) , \V94(10) , \V188(28) , \V30(11) , \V30(10) , \V144(31) ,
    \V94(17) , \V176(11) , \V144(30) , \V94(16) , \V176(10) , \V94(19) ,
    \V30(17) , \V176(13) , \V94(18) , \V30(16) , \V176(12) , \V126(27) ,
    \V94(23) , \V188(23) , \V30(2) , \V30(19) , \V176(15) , \V126(26) ,
    \V94(22) , \V188(22) , \V30(3) , \V127(0) , \V30(18) , \V176(14) ,
    \V126(29) , \V94(25) , \V188(25) , \V30(4) , \V30(23) , \V126(28) ,
    \V94(24) , \V188(24) , \V30(5) , \V30(22) , \V30(6) , \V30(25) ,
    \V30(7) , \V30(24) , \V144(27) , \V94(21) , \V30(8) , \V144(26) ,
    \V94(20) , \V30(9) , \V178(1) , \V144(29) , \V178(0) , \V30(21) ,
    \V144(28) , \V30(20) , \V126(21) , \V126(3) , \V126(20) , \V126(2) ,
    \V126(23) , \V94(27) , \V126(5) , \V126(22) , \V94(26) , \V64(0) ,
    \V126(4) , \V126(25) , \V94(29) , \V190(1) , \V30(27) , \V126(24) ,
    \V94(28) , \V190(0) , \V30(26) ,
    \V202(0)   );
  input  \V126(17) , \V144(21) , \V30(29) , \V126(1) , \V126(16) ,
    \V144(20) , \V30(28) , \V126(0) , \V126(19) , \V144(23) , \V126(18) ,
    \V144(22) , \V62(13) , \V144(25) , \V62(12) , \V191(31) , \V144(24) ,
    \V62(15) , \V94(31) , \V62(14) , \V126(7) , \V94(30) , \V126(6) ,
    \V144(19) , \V30(31) , \V201(3) , \V126(9) , \V144(18) , \V62(11) ,
    \V30(30) , \V201(2) , \V126(8) , \V126(11) , \V62(10) , \V201(5) ,
    \V126(10) , \V201(4) , \V126(13) , \V176(31) , \V126(12) , \V176(30) ,
    \V94(2) , \V126(15) , \V63(0) , \V201(1) , \V94(3) , \V126(14) ,
    \V62(17) , \V201(0) , \V94(4) , \V193(1) , \V62(16) , \V94(5) ,
    \V193(0) , \V62(19) , \V94(6) , \V62(18) , \V176(3) , \V94(7) ,
    \V62(23) , \V176(2) , \V94(8) , \V129(0) , \V62(22) , \V176(5) ,
    \V201(7) , \V94(9) , \V62(25) , \V176(4) , \V201(6) , \V62(24) ,
    \V176(27) , \V176(26) , \V176(1) , \V176(29) , \V62(21) , \V176(0) ,
    \V176(28) , \V62(20) , \V188(31) , \V176(7) , \V62(0) , \V188(30) ,
    \V62(27) , \V176(6) , \V62(1) , \V62(26) , \V176(9) , \V176(21) ,
    \V62(2) , \V62(29) , \V176(8) , \V176(20) , \V62(3) , \V62(28) ,
    \V176(23) , \V62(4) , \V176(22) , \V62(5) , \V94(13) , \V128(0) ,
    \V176(25) , \V62(6) , \V94(12) , \V176(24) , \V62(7) , \V94(15) ,
    \V30(13) , \V130(0) , \V176(17) , \V62(8) , \V94(14) , \V30(12) ,
    \V176(16) , \V62(9) , \V188(27) , \V30(15) , \V176(19) , \V188(26) ,
    \V62(31) , \V30(14) , \V126(31) , \V176(18) , \V94(11) , \V188(29) ,
    \V62(30) , \V126(30) , \V94(10) , \V188(28) , \V30(11) , \V30(10) ,
    \V144(31) , \V94(17) , \V176(11) , \V144(30) , \V94(16) , \V176(10) ,
    \V94(19) , \V30(17) , \V176(13) , \V94(18) , \V30(16) , \V176(12) ,
    \V126(27) , \V94(23) , \V188(23) , \V30(2) , \V30(19) , \V176(15) ,
    \V126(26) , \V94(22) , \V188(22) , \V30(3) , \V127(0) , \V30(18) ,
    \V176(14) , \V126(29) , \V94(25) , \V188(25) , \V30(4) , \V30(23) ,
    \V126(28) , \V94(24) , \V188(24) , \V30(5) , \V30(22) , \V30(6) ,
    \V30(25) , \V30(7) , \V30(24) , \V144(27) , \V94(21) , \V30(8) ,
    \V144(26) , \V94(20) , \V30(9) , \V178(1) , \V144(29) , \V178(0) ,
    \V30(21) , \V144(28) , \V30(20) , \V126(21) , \V126(3) , \V126(20) ,
    \V126(2) , \V126(23) , \V94(27) , \V126(5) , \V126(22) , \V94(26) ,
    \V64(0) , \V126(4) , \V126(25) , \V94(29) , \V190(1) , \V30(27) ,
    \V126(24) , \V94(28) , \V190(0) , \V30(26) ;
  output \V202(0) ;
  wire n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432;
  assign n203 = \V193(1)  & \V201(6) ;
  assign n204 = \V201(7)  & n203;
  assign n205 = \V191(31)  & \V201(7) ;
  assign n206 = \V201(6)  & n205;
  assign n207 = ~\V188(31)  & ~\V190(1) ;
  assign n208 = ~\V188(30)  & n207;
  assign n209 = ~\V190(0)  & n208;
  assign n210 = \V201(4)  & ~n209;
  assign n211 = \V201(5)  & n210;
  assign n212 = ~\V188(23)  & ~\V188(25) ;
  assign n213 = ~\V188(22)  & n212;
  assign n214 = ~\V188(24)  & n213;
  assign n215 = \V201(5)  & ~n214;
  assign n216 = \V201(4)  & n215;
  assign n217 = ~\V176(31)  & ~\V178(1) ;
  assign n218 = ~\V176(29)  & n217;
  assign n219 = ~\V176(27)  & n218;
  assign n220 = ~\V176(25)  & n219;
  assign n221 = ~\V176(23)  & n220;
  assign n222 = ~\V176(21)  & n221;
  assign n223 = ~\V176(19)  & n222;
  assign n224 = ~\V176(18)  & n223;
  assign n225 = ~\V176(20)  & n224;
  assign n226 = ~\V176(22)  & n225;
  assign n227 = ~\V176(24)  & n226;
  assign n228 = ~\V176(26)  & n227;
  assign n229 = ~\V176(28)  & n228;
  assign n230 = ~\V176(30)  & n229;
  assign n231 = ~\V178(0)  & n230;
  assign n232 = \V201(2)  & ~n231;
  assign n233 = \V201(3)  & n232;
  assign n234 = ~\V176(1)  & ~\V144(31) ;
  assign n235 = ~\V144(29)  & n234;
  assign n236 = ~\V144(27)  & n235;
  assign n237 = ~\V144(25)  & n236;
  assign n238 = ~\V144(23)  & n237;
  assign n239 = ~\V144(21)  & n238;
  assign n240 = ~\V144(19)  & n239;
  assign n241 = ~\V144(18)  & n240;
  assign n242 = ~\V144(20)  & n241;
  assign n243 = ~\V144(22)  & n242;
  assign n244 = ~\V144(24)  & n243;
  assign n245 = ~\V144(26)  & n244;
  assign n246 = ~\V144(28)  & n245;
  assign n247 = ~\V144(30)  & n246;
  assign n248 = ~\V176(0)  & n247;
  assign n249 = \V201(3)  & ~n248;
  assign n250 = \V201(2)  & n249;
  assign n251 = ~\V126(1)  & ~\V94(31) ;
  assign n252 = ~\V94(29)  & n251;
  assign n253 = ~\V94(27)  & n252;
  assign n254 = ~\V94(25)  & n253;
  assign n255 = ~\V94(23)  & n254;
  assign n256 = ~\V94(21)  & n255;
  assign n257 = ~\V94(19)  & n256;
  assign n258 = ~\V94(17)  & n257;
  assign n259 = ~\V94(15)  & n258;
  assign n260 = ~\V94(13)  & n259;
  assign n261 = ~\V94(11)  & n260;
  assign n262 = ~\V94(9)  & n261;
  assign n263 = ~\V94(7)  & n262;
  assign n264 = ~\V94(5)  & n263;
  assign n265 = ~\V94(3)  & n264;
  assign n266 = ~\V94(2)  & n265;
  assign n267 = ~\V94(4)  & n266;
  assign n268 = ~\V94(6)  & n267;
  assign n269 = ~\V94(8)  & n268;
  assign n270 = ~\V94(10)  & n269;
  assign n271 = ~\V94(12)  & n270;
  assign n272 = ~\V94(14)  & n271;
  assign n273 = ~\V94(16)  & n272;
  assign n274 = ~\V94(18)  & n273;
  assign n275 = ~\V94(20)  & n274;
  assign n276 = ~\V94(22)  & n275;
  assign n277 = ~\V94(24)  & n276;
  assign n278 = ~\V94(26)  & n277;
  assign n279 = ~\V94(28)  & n278;
  assign n280 = ~\V94(30)  & n279;
  assign n281 = ~\V126(0)  & n280;
  assign n282 = \V201(1)  & ~n281;
  assign n283 = \V201(0)  & n282;
  assign n284 = ~\V62(31)  & ~\V64(0) ;
  assign n285 = ~\V62(29)  & n284;
  assign n286 = ~\V62(27)  & n285;
  assign n287 = ~\V62(25)  & n286;
  assign n288 = ~\V62(23)  & n287;
  assign n289 = ~\V62(21)  & n288;
  assign n290 = ~\V62(19)  & n289;
  assign n291 = ~\V62(17)  & n290;
  assign n292 = ~\V62(15)  & n291;
  assign n293 = ~\V62(13)  & n292;
  assign n294 = ~\V62(11)  & n293;
  assign n295 = ~\V62(9)  & n294;
  assign n296 = ~\V62(7)  & n295;
  assign n297 = ~\V62(5)  & n296;
  assign n298 = ~\V62(3)  & n297;
  assign n299 = ~\V62(2)  & n298;
  assign n300 = ~\V62(4)  & n299;
  assign n301 = ~\V62(6)  & n300;
  assign n302 = ~\V62(8)  & n301;
  assign n303 = ~\V62(10)  & n302;
  assign n304 = ~\V62(12)  & n303;
  assign n305 = ~\V62(14)  & n304;
  assign n306 = ~\V62(16)  & n305;
  assign n307 = ~\V62(18)  & n306;
  assign n308 = ~\V62(20)  & n307;
  assign n309 = ~\V62(22)  & n308;
  assign n310 = ~\V62(24)  & n309;
  assign n311 = ~\V62(26)  & n310;
  assign n312 = ~\V62(28)  & n311;
  assign n313 = ~\V62(30)  & n312;
  assign n314 = ~\V63(0)  & n313;
  assign n315 = \V201(1)  & ~\V201(0) ;
  assign n316 = ~n314 & n315;
  assign n317 = ~\V201(0)  & \V129(0) ;
  assign n318 = ~\V30(31)  & ~\V62(1) ;
  assign n319 = ~\V30(29)  & n318;
  assign n320 = ~\V30(27)  & n319;
  assign n321 = ~\V30(25)  & n320;
  assign n322 = ~\V30(23)  & n321;
  assign n323 = ~\V30(21)  & n322;
  assign n324 = ~\V30(19)  & n323;
  assign n325 = ~\V30(17)  & n324;
  assign n326 = ~\V30(15)  & n325;
  assign n327 = ~\V30(13)  & n326;
  assign n328 = ~\V30(11)  & n327;
  assign n329 = ~\V30(9)  & n328;
  assign n330 = ~\V30(7)  & n329;
  assign n331 = ~\V30(5)  & n330;
  assign n332 = ~\V30(3)  & n331;
  assign n333 = ~\V30(2)  & n332;
  assign n334 = ~\V30(4)  & n333;
  assign n335 = ~\V30(6)  & n334;
  assign n336 = ~\V30(8)  & n335;
  assign n337 = ~\V30(10)  & n336;
  assign n338 = ~\V30(12)  & n337;
  assign n339 = ~\V30(14)  & n338;
  assign n340 = ~\V30(16)  & n339;
  assign n341 = ~\V30(18)  & n340;
  assign n342 = ~\V30(20)  & n341;
  assign n343 = ~\V30(22)  & n342;
  assign n344 = ~\V30(24)  & n343;
  assign n345 = ~\V30(26)  & n344;
  assign n346 = ~\V30(28)  & n345;
  assign n347 = ~\V30(30)  & n346;
  assign n348 = ~\V62(0)  & n347;
  assign n349 = n315 & ~n348;
  assign n350 = \V201(0)  & \V130(0) ;
  assign n351 = ~\V128(0)  & ~\V126(31) ;
  assign n352 = ~\V126(29)  & n351;
  assign n353 = ~\V126(27)  & n352;
  assign n354 = ~\V126(25)  & n353;
  assign n355 = ~\V126(23)  & n354;
  assign n356 = ~\V126(21)  & n355;
  assign n357 = ~\V126(19)  & n356;
  assign n358 = ~\V126(17)  & n357;
  assign n359 = ~\V126(15)  & n358;
  assign n360 = ~\V126(13)  & n359;
  assign n361 = ~\V126(11)  & n360;
  assign n362 = ~\V126(9)  & n361;
  assign n363 = ~\V126(7)  & n362;
  assign n364 = ~\V126(5)  & n363;
  assign n365 = ~\V126(3)  & n364;
  assign n366 = ~\V126(2)  & n365;
  assign n367 = ~\V126(4)  & n366;
  assign n368 = ~\V126(6)  & n367;
  assign n369 = ~\V126(8)  & n368;
  assign n370 = ~\V126(10)  & n369;
  assign n371 = ~\V126(12)  & n370;
  assign n372 = ~\V126(14)  & n371;
  assign n373 = ~\V126(16)  & n372;
  assign n374 = ~\V126(18)  & n373;
  assign n375 = ~\V126(20)  & n374;
  assign n376 = ~\V126(22)  & n375;
  assign n377 = ~\V126(24)  & n376;
  assign n378 = ~\V126(26)  & n377;
  assign n379 = ~\V126(28)  & n378;
  assign n380 = ~\V126(30)  & n379;
  assign n381 = ~\V127(0)  & n380;
  assign n382 = \V201(1)  & ~n381;
  assign n383 = \V201(0)  & n382;
  assign n384 = ~\V176(17)  & ~\V176(15) ;
  assign n385 = ~\V176(13)  & n384;
  assign n386 = ~\V176(11)  & n385;
  assign n387 = ~\V176(9)  & n386;
  assign n388 = ~\V176(7)  & n387;
  assign n389 = ~\V176(5)  & n388;
  assign n390 = ~\V176(3)  & n389;
  assign n391 = ~\V176(2)  & n390;
  assign n392 = ~\V176(4)  & n391;
  assign n393 = ~\V176(6)  & n392;
  assign n394 = ~\V176(8)  & n393;
  assign n395 = ~\V176(10)  & n394;
  assign n396 = ~\V176(12)  & n395;
  assign n397 = ~\V176(14)  & n396;
  assign n398 = ~\V176(16)  & n397;
  assign n399 = \V201(2)  & ~n398;
  assign n400 = \V201(3)  & n399;
  assign n401 = \V201(3)  & ~n231;
  assign n402 = ~\V188(27)  & ~\V188(29) ;
  assign n403 = ~\V188(26)  & n402;
  assign n404 = ~\V188(28)  & n403;
  assign n405 = \V201(4)  & ~n404;
  assign n406 = \V201(5)  & n405;
  assign n407 = \V201(5)  & ~n209;
  assign n408 = \V193(0)  & \V201(6) ;
  assign n409 = \V201(7)  & n408;
  assign n410 = \V193(1)  & \V201(7) ;
  assign n411 = ~n408 & ~n410;
  assign n412 = ~n409 & n411;
  assign n413 = ~n407 & n412;
  assign n414 = ~n405 & n413;
  assign n415 = ~n406 & n414;
  assign n416 = ~n401 & n415;
  assign n417 = ~n399 & n416;
  assign n418 = ~n400 & n417;
  assign n419 = ~n383 & n418;
  assign n420 = ~n350 & n419;
  assign n421 = ~n349 & n420;
  assign n422 = ~n317 & n421;
  assign n423 = ~n316 & n422;
  assign n424 = ~n283 & n423;
  assign n425 = ~n250 & n424;
  assign n426 = ~n233 & n425;
  assign n427 = ~n232 & n426;
  assign n428 = ~n216 & n427;
  assign n429 = ~n211 & n428;
  assign n430 = ~n210 & n429;
  assign n431 = ~n206 & n430;
  assign n432 = ~n204 & n431;
  assign \V202(0)  = n203 | ~n432;
endmodule


