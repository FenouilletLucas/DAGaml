// Benchmark "i9" written by ABC on Tue May 16 16:07:51 2017

module i9 ( 
    \V9(10) , \V56(0) , \V56(1) , \V56(2) , \V56(3) , \V56(4) , \V56(5) ,
    \V56(6) , \V56(7) , \V56(8) , \V56(9) , \V24(13) , \V24(12) ,
    \V24(14) , \V24(11) , \V24(10) , \V9(0) , \V9(1) , \V9(2) , \V9(3) ,
    \V9(5) , \V9(6) , \V9(7) , \V9(8) , \V88(13) , \V88(12) , \V88(15) ,
    \V88(14) , \V88(11) , \V88(10) , \V88(0) , \V88(1) , \V88(2) ,
    \V88(3) , \V88(17) , \V88(4) , \V88(16) , \V88(5) , \V88(19) ,
    \V88(6) , \V88(18) , \V88(7) , \V88(23) , \V88(8) , \V88(22) ,
    \V88(9) , \V88(25) , \V88(24) , \V88(21) , \V88(20) , \V88(27) ,
    \V88(26) , \V88(29) , \V88(28) , \V88(31) , \V88(30) , \V56(13) ,
    \V56(12) , \V56(15) , \V56(14) , \V24(0) , \V56(11) , \V24(1) ,
    \V56(10) , \V24(2) , \V24(3) , \V24(4) , \V24(5) , \V24(6) , \V56(17) ,
    \V24(7) , \V56(16) , \V24(8) , \V56(19) , \V24(9) , \V56(18) ,
    \V56(23) , \V56(22) , \V56(25) , \V56(24) , \V56(21) , \V56(20) ,
    \V56(27) , \V56(26) , \V56(29) , \V56(28) , \V56(31) , \V56(30) ,
    \V151(27) , \V151(26) , \V151(29) , \V151(28) , \V151(21) , \V151(20) ,
    \V151(23) , \V151(22) , \V119(27) , \V151(25) , \V119(26) , \V151(24) ,
    \V119(29) , \V151(17) , \V119(28) , \V151(16) , \V151(19) , \V151(18) ,
    \V119(21) , \V119(20) , \V119(23) , \V151(11) , \V119(22) , \V151(10) ,
    \V119(25) , \V151(3) , \V151(13) , \V119(24) , \V151(2) , \V151(12) ,
    \V119(17) , \V151(5) , \V151(15) , \V119(16) , \V151(4) , \V151(14) ,
    \V119(19) , \V119(18) , \V151(1) , \V151(0) , \V119(11) , \V151(7) ,
    \V119(10) , \V151(6) , \V119(13) , \V151(9) , \V119(12) , \V151(8) ,
    \V119(15) , \V119(14) , \V151(31) , \V151(30) , \V119(30) , \V119(3) ,
    \V119(2) , \V119(5) , \V119(4) , \V119(1) , \V119(0) , \V119(7) ,
    \V119(6) , \V119(9) , \V119(8)   );
  input  \V9(10) , \V56(0) , \V56(1) , \V56(2) , \V56(3) , \V56(4) ,
    \V56(5) , \V56(6) , \V56(7) , \V56(8) , \V56(9) , \V24(13) , \V24(12) ,
    \V24(14) , \V24(11) , \V24(10) , \V9(0) , \V9(1) , \V9(2) , \V9(3) ,
    \V9(5) , \V9(6) , \V9(7) , \V9(8) , \V88(13) , \V88(12) , \V88(15) ,
    \V88(14) , \V88(11) , \V88(10) , \V88(0) , \V88(1) , \V88(2) ,
    \V88(3) , \V88(17) , \V88(4) , \V88(16) , \V88(5) , \V88(19) ,
    \V88(6) , \V88(18) , \V88(7) , \V88(23) , \V88(8) , \V88(22) ,
    \V88(9) , \V88(25) , \V88(24) , \V88(21) , \V88(20) , \V88(27) ,
    \V88(26) , \V88(29) , \V88(28) , \V88(31) , \V88(30) , \V56(13) ,
    \V56(12) , \V56(15) , \V56(14) , \V24(0) , \V56(11) , \V24(1) ,
    \V56(10) , \V24(2) , \V24(3) , \V24(4) , \V24(5) , \V24(6) , \V56(17) ,
    \V24(7) , \V56(16) , \V24(8) , \V56(19) , \V24(9) , \V56(18) ,
    \V56(23) , \V56(22) , \V56(25) , \V56(24) , \V56(21) , \V56(20) ,
    \V56(27) , \V56(26) , \V56(29) , \V56(28) , \V56(31) , \V56(30) ;
  output \V151(27) , \V151(26) , \V151(29) , \V151(28) , \V151(21) ,
    \V151(20) , \V151(23) , \V151(22) , \V119(27) , \V151(25) , \V119(26) ,
    \V151(24) , \V119(29) , \V151(17) , \V119(28) , \V151(16) , \V151(19) ,
    \V151(18) , \V119(21) , \V119(20) , \V119(23) , \V151(11) , \V119(22) ,
    \V151(10) , \V119(25) , \V151(3) , \V151(13) , \V119(24) , \V151(2) ,
    \V151(12) , \V119(17) , \V151(5) , \V151(15) , \V119(16) , \V151(4) ,
    \V151(14) , \V119(19) , \V119(18) , \V151(1) , \V151(0) , \V119(11) ,
    \V151(7) , \V119(10) , \V151(6) , \V119(13) , \V151(9) , \V119(12) ,
    \V151(8) , \V119(15) , \V119(14) , \V151(31) , \V151(30) , \V119(30) ,
    \V119(3) , \V119(2) , \V119(5) , \V119(4) , \V119(1) , \V119(0) ,
    \V119(7) , \V119(6) , \V119(9) , \V119(8) ;
  wire n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n414, n415,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n951, n952, n953, n954, n955, n956, n957, n958, n960,
    n961, n962, n963, n964, n965, n966, n967, n969, n970, n971, n972, n973,
    n974, n975, n976, n978, n979, n980, n981, n982, n983, n984, n985, n987,
    n988, n989, n990, n991, n992, n993, n994, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  assign n152 = ~\V9(10)  & \V9(2) ;
  assign n153 = ~\V9(1)  & n152;
  assign n154 = \V9(8)  & n153;
  assign n155 = ~\V9(10)  & ~\V9(5) ;
  assign n156 = ~\V9(1)  & n155;
  assign n157 = \V9(0)  & n156;
  assign n158 = \V9(2)  & n157;
  assign n159 = ~\V9(6)  & n158;
  assign n160 = \V9(1)  & n152;
  assign n161 = ~\V9(3)  & n160;
  assign n162 = ~\V9(10)  & \V9(1) ;
  assign n163 = \V9(8)  & n162;
  assign n164 = \V9(1)  & n155;
  assign n165 = ~\V9(2)  & n164;
  assign n166 = ~\V9(6)  & n165;
  assign n167 = ~\V9(10)  & ~\V9(0) ;
  assign n168 = ~\V9(5)  & n167;
  assign n169 = \V9(7)  & n167;
  assign n170 = \V9(1)  & \V9(3) ;
  assign n171 = \V9(2)  & n170;
  assign n172 = \V9(10)  & \V9(1) ;
  assign n173 = \V9(10)  & \V9(2) ;
  assign n174 = ~\V9(2)  & ~\V9(6) ;
  assign n175 = ~\V9(1)  & n174;
  assign n176 = ~\V9(5)  & n175;
  assign n177 = ~\V9(1)  & \V9(7) ;
  assign n178 = ~\V9(2)  & n177;
  assign n179 = \V9(10)  & ~\V9(1) ;
  assign n180 = ~\V9(2)  & n179;
  assign n181 = ~n178 & ~n180;
  assign n182 = ~n176 & n181;
  assign n183 = ~n173 & n182;
  assign n184 = ~n172 & n183;
  assign n185 = ~n171 & n184;
  assign n186 = ~n169 & n185;
  assign n187 = ~n168 & n186;
  assign n188 = ~n166 & n187;
  assign n189 = ~n163 & n188;
  assign n190 = ~n161 & n189;
  assign n191 = ~n159 & n190;
  assign n192 = ~n154 & n191;
  assign n193 = ~n154 & ~n159;
  assign n194 = ~n161 & n193;
  assign n195 = ~n178 & n194;
  assign n196 = ~n176 & n195;
  assign n197 = ~n180 & n196;
  assign n198 = ~n163 & ~n169;
  assign n199 = ~n168 & n198;
  assign n200 = ~n166 & n199;
  assign n201 = ~n178 & n200;
  assign n202 = ~n176 & n201;
  assign n203 = ~n180 & n202;
  assign n204 = \V88(12)  & ~n203;
  assign n205 = ~n197 & n204;
  assign n206 = ~n192 & n205;
  assign n207 = \V88(16)  & n203;
  assign n208 = ~n197 & n207;
  assign n209 = ~n192 & n208;
  assign n210 = \V88(19)  & ~n203;
  assign n211 = n197 & n210;
  assign n212 = ~n192 & n211;
  assign n213 = \V88(27)  & n203;
  assign n214 = n197 & n213;
  assign n215 = ~n192 & n214;
  assign n216 = n192 & ~n197;
  assign n217 = ~n203 & n216;
  assign n218 = n203 & n216;
  assign n219 = n192 & n197;
  assign n220 = ~n203 & n219;
  assign n221 = n203 & n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~n218 & n222;
  assign n224 = ~n217 & n223;
  assign n225 = ~n215 & n224;
  assign n226 = ~n212 & n225;
  assign n227 = ~n209 & n226;
  assign \V151(27)  = n206 | ~n227;
  assign n229 = \V88(11)  & ~n203;
  assign n230 = ~n197 & n229;
  assign n231 = ~n192 & n230;
  assign n232 = \V88(15)  & n203;
  assign n233 = ~n197 & n232;
  assign n234 = ~n192 & n233;
  assign n235 = \V88(18)  & ~n203;
  assign n236 = n197 & n235;
  assign n237 = ~n192 & n236;
  assign n238 = \V88(26)  & n203;
  assign n239 = n197 & n238;
  assign n240 = ~n192 & n239;
  assign n241 = n224 & ~n240;
  assign n242 = ~n237 & n241;
  assign n243 = ~n234 & n242;
  assign \V151(26)  = n231 | ~n243;
  assign n245 = \V88(14)  & ~n203;
  assign n246 = ~n197 & n245;
  assign n247 = ~n192 & n246;
  assign n248 = \V88(18)  & n203;
  assign n249 = ~n197 & n248;
  assign n250 = ~n192 & n249;
  assign n251 = \V88(21)  & ~n203;
  assign n252 = n197 & n251;
  assign n253 = ~n192 & n252;
  assign n254 = \V88(29)  & n203;
  assign n255 = n197 & n254;
  assign n256 = ~n192 & n255;
  assign n257 = n224 & ~n256;
  assign n258 = ~n253 & n257;
  assign n259 = ~n250 & n258;
  assign \V151(29)  = n247 | ~n259;
  assign n261 = \V88(13)  & ~n203;
  assign n262 = ~n197 & n261;
  assign n263 = ~n192 & n262;
  assign n264 = \V88(17)  & n203;
  assign n265 = ~n197 & n264;
  assign n266 = ~n192 & n265;
  assign n267 = \V88(20)  & ~n203;
  assign n268 = n197 & n267;
  assign n269 = ~n192 & n268;
  assign n270 = \V88(28)  & n203;
  assign n271 = n197 & n270;
  assign n272 = ~n192 & n271;
  assign n273 = n224 & ~n272;
  assign n274 = ~n269 & n273;
  assign n275 = ~n266 & n274;
  assign \V151(28)  = n263 | ~n275;
  assign n277 = \V88(6)  & ~n203;
  assign n278 = ~n197 & n277;
  assign n279 = ~n192 & n278;
  assign n280 = \V88(10)  & n203;
  assign n281 = ~n197 & n280;
  assign n282 = ~n192 & n281;
  assign n283 = n197 & n261;
  assign n284 = ~n192 & n283;
  assign n285 = \V88(21)  & n203;
  assign n286 = n197 & n285;
  assign n287 = ~n192 & n286;
  assign n288 = n224 & ~n287;
  assign n289 = ~n284 & n288;
  assign n290 = ~n282 & n289;
  assign \V151(21)  = n279 | ~n290;
  assign n292 = \V88(5)  & ~n203;
  assign n293 = ~n197 & n292;
  assign n294 = ~n192 & n293;
  assign n295 = \V88(9)  & n203;
  assign n296 = ~n197 & n295;
  assign n297 = ~n192 & n296;
  assign n298 = n197 & n204;
  assign n299 = ~n192 & n298;
  assign n300 = \V88(20)  & n203;
  assign n301 = n197 & n300;
  assign n302 = ~n192 & n301;
  assign n303 = n224 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~n297 & n304;
  assign \V151(20)  = n294 | ~n305;
  assign n307 = \V88(8)  & ~n203;
  assign n308 = ~n197 & n307;
  assign n309 = ~n192 & n308;
  assign n310 = \V88(12)  & n203;
  assign n311 = ~n197 & n310;
  assign n312 = ~n192 & n311;
  assign n313 = \V88(15)  & ~n203;
  assign n314 = n197 & n313;
  assign n315 = ~n192 & n314;
  assign n316 = \V88(23)  & n203;
  assign n317 = n197 & n316;
  assign n318 = ~n192 & n317;
  assign n319 = n224 & ~n318;
  assign n320 = ~n315 & n319;
  assign n321 = ~n312 & n320;
  assign \V151(23)  = n309 | ~n321;
  assign n323 = \V88(7)  & ~n203;
  assign n324 = ~n197 & n323;
  assign n325 = ~n192 & n324;
  assign n326 = \V88(11)  & n203;
  assign n327 = ~n197 & n326;
  assign n328 = ~n192 & n327;
  assign n329 = n197 & n245;
  assign n330 = ~n192 & n329;
  assign n331 = \V88(22)  & n203;
  assign n332 = n197 & n331;
  assign n333 = ~n192 & n332;
  assign n334 = n224 & ~n333;
  assign n335 = ~n330 & n334;
  assign n336 = ~n328 & n335;
  assign \V151(22)  = n325 | ~n336;
  assign n338 = \V56(13)  & ~n203;
  assign n339 = ~n197 & n338;
  assign n340 = ~n192 & n339;
  assign n341 = \V56(17)  & n203;
  assign n342 = ~n197 & n341;
  assign n343 = ~n192 & n342;
  assign n344 = ~n192 & n197;
  assign n345 = ~n203 & n344;
  assign n346 = \V56(20)  & n345;
  assign n347 = \V56(28)  & n203;
  assign n348 = n197 & n347;
  assign n349 = ~n192 & n348;
  assign n350 = ~n192 & ~n349;
  assign n351 = ~n346 & n350;
  assign n352 = ~n343 & n351;
  assign \V119(27)  = n340 | ~n352;
  assign n354 = \V88(10)  & ~n203;
  assign n355 = ~n197 & n354;
  assign n356 = ~n192 & n355;
  assign n357 = \V88(14)  & n203;
  assign n358 = ~n197 & n357;
  assign n359 = ~n192 & n358;
  assign n360 = \V88(17)  & ~n203;
  assign n361 = n197 & n360;
  assign n362 = ~n192 & n361;
  assign n363 = \V88(25)  & n203;
  assign n364 = n197 & n363;
  assign n365 = ~n192 & n364;
  assign n366 = n224 & ~n365;
  assign n367 = ~n362 & n366;
  assign n368 = ~n359 & n367;
  assign \V151(25)  = n356 | ~n368;
  assign n370 = \V56(12)  & ~n203;
  assign n371 = ~n197 & n370;
  assign n372 = ~n192 & n371;
  assign n373 = \V56(16)  & n203;
  assign n374 = ~n197 & n373;
  assign n375 = ~n192 & n374;
  assign n376 = \V56(19)  & n345;
  assign n377 = \V56(27)  & n203;
  assign n378 = n197 & n377;
  assign n379 = ~n192 & n378;
  assign n380 = ~n192 & ~n379;
  assign n381 = ~n376 & n380;
  assign n382 = ~n375 & n381;
  assign \V119(26)  = n372 | ~n382;
  assign n384 = \V88(9)  & ~n203;
  assign n385 = ~n197 & n384;
  assign n386 = ~n192 & n385;
  assign n387 = \V88(13)  & n203;
  assign n388 = ~n197 & n387;
  assign n389 = ~n192 & n388;
  assign n390 = \V88(16)  & ~n203;
  assign n391 = n197 & n390;
  assign n392 = ~n192 & n391;
  assign n393 = \V88(24)  & n203;
  assign n394 = n197 & n393;
  assign n395 = ~n192 & n394;
  assign n396 = n224 & ~n395;
  assign n397 = ~n392 & n396;
  assign n398 = ~n389 & n397;
  assign \V151(24)  = n386 | ~n398;
  assign n400 = \V56(15)  & ~n203;
  assign n401 = ~n197 & n400;
  assign n402 = ~n192 & n401;
  assign n403 = \V56(19)  & n203;
  assign n404 = ~n197 & n403;
  assign n405 = ~n192 & n404;
  assign n406 = \V56(22)  & n345;
  assign n407 = \V56(30)  & n203;
  assign n408 = n197 & n407;
  assign n409 = ~n192 & n408;
  assign n410 = ~n192 & ~n409;
  assign n411 = ~n406 & n410;
  assign n412 = ~n405 & n411;
  assign \V119(29)  = n402 | ~n412;
  assign n414 = \V88(2)  & ~n203;
  assign n415 = ~n197 & n414;
  assign n416 = ~n192 & n415;
  assign n417 = \V88(6)  & n203;
  assign n418 = ~n197 & n417;
  assign n419 = ~n192 & n418;
  assign n420 = n197 & n384;
  assign n421 = ~n192 & n420;
  assign n422 = n197 & n264;
  assign n423 = ~n192 & n422;
  assign n424 = n224 & ~n423;
  assign n425 = ~n421 & n424;
  assign n426 = ~n419 & n425;
  assign \V151(17)  = n416 | ~n426;
  assign n428 = \V56(14)  & ~n203;
  assign n429 = ~n197 & n428;
  assign n430 = ~n192 & n429;
  assign n431 = \V56(18)  & n203;
  assign n432 = ~n197 & n431;
  assign n433 = ~n192 & n432;
  assign n434 = \V56(21)  & n345;
  assign n435 = \V56(29)  & n203;
  assign n436 = n197 & n435;
  assign n437 = ~n192 & n436;
  assign n438 = ~n192 & ~n437;
  assign n439 = ~n434 & n438;
  assign n440 = ~n433 & n439;
  assign \V119(28)  = n430 | ~n440;
  assign n442 = \V88(1)  & ~n203;
  assign n443 = ~n197 & n442;
  assign n444 = ~n192 & n443;
  assign n445 = \V88(5)  & n203;
  assign n446 = ~n197 & n445;
  assign n447 = ~n192 & n446;
  assign n448 = n197 & n307;
  assign n449 = ~n192 & n448;
  assign n450 = n197 & n207;
  assign n451 = ~n192 & n450;
  assign n452 = n224 & ~n451;
  assign n453 = ~n449 & n452;
  assign n454 = ~n447 & n453;
  assign \V151(16)  = n444 | ~n454;
  assign n456 = \V88(4)  & ~n203;
  assign n457 = ~n197 & n456;
  assign n458 = ~n192 & n457;
  assign n459 = \V88(8)  & n203;
  assign n460 = ~n197 & n459;
  assign n461 = ~n192 & n460;
  assign n462 = n197 & n229;
  assign n463 = ~n192 & n462;
  assign n464 = \V88(19)  & n203;
  assign n465 = n197 & n464;
  assign n466 = ~n192 & n465;
  assign n467 = n224 & ~n466;
  assign n468 = ~n463 & n467;
  assign n469 = ~n461 & n468;
  assign \V151(19)  = n458 | ~n469;
  assign n471 = \V88(3)  & ~n203;
  assign n472 = ~n197 & n471;
  assign n473 = ~n192 & n472;
  assign n474 = \V88(7)  & n203;
  assign n475 = ~n197 & n474;
  assign n476 = ~n192 & n475;
  assign n477 = n197 & n354;
  assign n478 = ~n192 & n477;
  assign n479 = n197 & n248;
  assign n480 = ~n192 & n479;
  assign n481 = n224 & ~n480;
  assign n482 = ~n478 & n481;
  assign n483 = ~n476 & n482;
  assign \V151(18)  = n473 | ~n483;
  assign n485 = \V56(7)  & ~n203;
  assign n486 = ~n197 & n485;
  assign n487 = ~n192 & n486;
  assign n488 = \V56(11)  & n203;
  assign n489 = ~n197 & n488;
  assign n490 = ~n192 & n489;
  assign n491 = \V56(14)  & n345;
  assign n492 = \V56(22)  & n203;
  assign n493 = n197 & n492;
  assign n494 = ~n192 & n493;
  assign n495 = ~n192 & ~n494;
  assign n496 = ~n491 & n495;
  assign n497 = ~n490 & n496;
  assign \V119(21)  = n487 | ~n497;
  assign n499 = \V56(6)  & ~n203;
  assign n500 = ~n197 & n499;
  assign n501 = ~n192 & n500;
  assign n502 = \V56(10)  & n203;
  assign n503 = ~n197 & n502;
  assign n504 = ~n192 & n503;
  assign n505 = \V56(13)  & n345;
  assign n506 = \V56(21)  & n203;
  assign n507 = n197 & n506;
  assign n508 = ~n192 & n507;
  assign n509 = ~n192 & ~n508;
  assign n510 = ~n505 & n509;
  assign n511 = ~n504 & n510;
  assign \V119(20)  = n501 | ~n511;
  assign n513 = \V56(9)  & ~n203;
  assign n514 = ~n197 & n513;
  assign n515 = ~n192 & n514;
  assign n516 = \V56(13)  & n203;
  assign n517 = ~n197 & n516;
  assign n518 = ~n192 & n517;
  assign n519 = \V56(16)  & n345;
  assign n520 = \V56(24)  & n203;
  assign n521 = n197 & n520;
  assign n522 = ~n192 & n521;
  assign n523 = ~n192 & ~n522;
  assign n524 = ~n519 & n523;
  assign n525 = ~n518 & n524;
  assign \V119(23)  = n515 | ~n525;
  assign n527 = \V56(28)  & ~n203;
  assign n528 = ~n197 & n527;
  assign n529 = ~n192 & n528;
  assign n530 = \V88(0)  & n203;
  assign n531 = ~n197 & n530;
  assign n532 = ~n192 & n531;
  assign n533 = n197 & n471;
  assign n534 = ~n192 & n533;
  assign n535 = n197 & n326;
  assign n536 = ~n192 & n535;
  assign n537 = n224 & ~n536;
  assign n538 = ~n534 & n537;
  assign n539 = ~n532 & n538;
  assign \V151(11)  = n529 | ~n539;
  assign n541 = \V56(8)  & ~n203;
  assign n542 = ~n197 & n541;
  assign n543 = ~n192 & n542;
  assign n544 = \V56(12)  & n203;
  assign n545 = ~n197 & n544;
  assign n546 = ~n192 & n545;
  assign n547 = \V56(15)  & n345;
  assign n548 = \V56(23)  & n203;
  assign n549 = n197 & n548;
  assign n550 = ~n192 & n549;
  assign n551 = ~n192 & ~n550;
  assign n552 = ~n547 & n551;
  assign n553 = ~n546 & n552;
  assign \V119(22)  = n543 | ~n553;
  assign n555 = \V56(27)  & ~n203;
  assign n556 = ~n197 & n555;
  assign n557 = ~n192 & n556;
  assign n558 = \V56(31)  & n203;
  assign n559 = ~n197 & n558;
  assign n560 = ~n192 & n559;
  assign n561 = n197 & n414;
  assign n562 = ~n192 & n561;
  assign n563 = n197 & n280;
  assign n564 = ~n192 & n563;
  assign n565 = n224 & ~n564;
  assign n566 = ~n562 & n565;
  assign n567 = ~n560 & n566;
  assign \V151(10)  = n557 | ~n567;
  assign n569 = \V56(11)  & ~n203;
  assign n570 = ~n197 & n569;
  assign n571 = ~n192 & n570;
  assign n572 = \V56(15)  & n203;
  assign n573 = ~n197 & n572;
  assign n574 = ~n192 & n573;
  assign n575 = \V56(18)  & n345;
  assign n576 = \V56(26)  & n203;
  assign n577 = n197 & n576;
  assign n578 = ~n192 & n577;
  assign n579 = ~n192 & ~n578;
  assign n580 = ~n575 & n579;
  assign n581 = ~n574 & n580;
  assign \V119(25)  = n571 | ~n581;
  assign n583 = \V56(20)  & ~n203;
  assign n584 = ~n197 & n583;
  assign n585 = ~n192 & n584;
  assign n586 = ~n197 & n520;
  assign n587 = ~n192 & n586;
  assign n588 = n197 & n555;
  assign n589 = ~n192 & n588;
  assign n590 = \V88(3)  & n203;
  assign n591 = n197 & n590;
  assign n592 = ~n192 & n591;
  assign n593 = n224 & ~n592;
  assign n594 = ~n589 & n593;
  assign n595 = ~n587 & n594;
  assign \V151(3)  = n585 | ~n595;
  assign n597 = \V56(30)  & ~n203;
  assign n598 = ~n197 & n597;
  assign n599 = ~n192 & n598;
  assign n600 = \V88(2)  & n203;
  assign n601 = ~n197 & n600;
  assign n602 = ~n192 & n601;
  assign n603 = n197 & n292;
  assign n604 = ~n192 & n603;
  assign n605 = n197 & n387;
  assign n606 = ~n192 & n605;
  assign n607 = n224 & ~n606;
  assign n608 = ~n604 & n607;
  assign n609 = ~n602 & n608;
  assign \V151(13)  = n599 | ~n609;
  assign n611 = \V56(10)  & ~n203;
  assign n612 = ~n197 & n611;
  assign n613 = ~n192 & n612;
  assign n614 = \V56(14)  & n203;
  assign n615 = ~n197 & n614;
  assign n616 = ~n192 & n615;
  assign n617 = \V56(17)  & n345;
  assign n618 = \V56(25)  & n203;
  assign n619 = n197 & n618;
  assign n620 = ~n192 & n619;
  assign n621 = ~n192 & ~n620;
  assign n622 = ~n617 & n621;
  assign n623 = ~n616 & n622;
  assign \V119(24)  = n613 | ~n623;
  assign n625 = \V56(19)  & ~n203;
  assign n626 = ~n197 & n625;
  assign n627 = ~n192 & n626;
  assign n628 = ~n197 & n548;
  assign n629 = ~n192 & n628;
  assign n630 = \V56(26)  & ~n203;
  assign n631 = n197 & n630;
  assign n632 = ~n192 & n631;
  assign n633 = n197 & n600;
  assign n634 = ~n192 & n633;
  assign n635 = n224 & ~n634;
  assign n636 = ~n632 & n635;
  assign n637 = ~n629 & n636;
  assign \V151(2)  = n627 | ~n637;
  assign n639 = \V56(29)  & ~n203;
  assign n640 = ~n197 & n639;
  assign n641 = ~n192 & n640;
  assign n642 = \V88(1)  & n203;
  assign n643 = ~n197 & n642;
  assign n644 = ~n192 & n643;
  assign n645 = n197 & n456;
  assign n646 = ~n192 & n645;
  assign n647 = n197 & n310;
  assign n648 = ~n192 & n647;
  assign n649 = n224 & ~n648;
  assign n650 = ~n646 & n649;
  assign n651 = ~n644 & n650;
  assign \V151(12)  = n641 | ~n651;
  assign n653 = \V56(3)  & ~n203;
  assign n654 = ~n197 & n653;
  assign n655 = ~n192 & n654;
  assign n656 = \V56(7)  & n203;
  assign n657 = ~n197 & n656;
  assign n658 = ~n192 & n657;
  assign n659 = \V56(10)  & n345;
  assign n660 = n197 & n431;
  assign n661 = ~n192 & n660;
  assign n662 = ~n192 & ~n661;
  assign n663 = ~n659 & n662;
  assign n664 = ~n658 & n663;
  assign \V119(17)  = n655 | ~n664;
  assign n666 = \V56(22)  & ~n203;
  assign n667 = ~n197 & n666;
  assign n668 = ~n192 & n667;
  assign n669 = ~n197 & n576;
  assign n670 = ~n192 & n669;
  assign n671 = n197 & n639;
  assign n672 = ~n192 & n671;
  assign n673 = n197 & n445;
  assign n674 = ~n192 & n673;
  assign n675 = n224 & ~n674;
  assign n676 = ~n672 & n675;
  assign n677 = ~n670 & n676;
  assign \V151(5)  = n668 | ~n677;
  assign n679 = \V88(0)  & ~n203;
  assign n680 = ~n197 & n679;
  assign n681 = ~n192 & n680;
  assign n682 = \V88(4)  & n203;
  assign n683 = ~n197 & n682;
  assign n684 = ~n192 & n683;
  assign n685 = n197 & n323;
  assign n686 = ~n192 & n685;
  assign n687 = n197 & n232;
  assign n688 = ~n192 & n687;
  assign n689 = n224 & ~n688;
  assign n690 = ~n686 & n689;
  assign n691 = ~n684 & n690;
  assign \V151(15)  = n681 | ~n691;
  assign n693 = \V56(2)  & ~n203;
  assign n694 = ~n197 & n693;
  assign n695 = ~n192 & n694;
  assign n696 = \V56(6)  & n203;
  assign n697 = ~n197 & n696;
  assign n698 = ~n192 & n697;
  assign n699 = \V56(9)  & n345;
  assign n700 = n197 & n341;
  assign n701 = ~n192 & n700;
  assign n702 = ~n192 & ~n701;
  assign n703 = ~n699 & n702;
  assign n704 = ~n698 & n703;
  assign \V119(16)  = n695 | ~n704;
  assign n706 = \V56(21)  & ~n203;
  assign n707 = ~n197 & n706;
  assign n708 = ~n192 & n707;
  assign n709 = ~n197 & n618;
  assign n710 = ~n192 & n709;
  assign n711 = n197 & n527;
  assign n712 = ~n192 & n711;
  assign n713 = n197 & n682;
  assign n714 = ~n192 & n713;
  assign n715 = n224 & ~n714;
  assign n716 = ~n712 & n715;
  assign n717 = ~n710 & n716;
  assign \V151(4)  = n708 | ~n717;
  assign n719 = \V56(31)  & ~n203;
  assign n720 = ~n197 & n719;
  assign n721 = ~n192 & n720;
  assign n722 = ~n197 & n590;
  assign n723 = ~n192 & n722;
  assign n724 = n197 & n277;
  assign n725 = ~n192 & n724;
  assign n726 = n197 & n357;
  assign n727 = ~n192 & n726;
  assign n728 = n224 & ~n727;
  assign n729 = ~n725 & n728;
  assign n730 = ~n723 & n729;
  assign \V151(14)  = n721 | ~n730;
  assign n732 = \V56(5)  & ~n203;
  assign n733 = ~n197 & n732;
  assign n734 = ~n192 & n733;
  assign n735 = \V56(9)  & n203;
  assign n736 = ~n197 & n735;
  assign n737 = ~n192 & n736;
  assign n738 = \V56(12)  & n345;
  assign n739 = \V56(20)  & n203;
  assign n740 = n197 & n739;
  assign n741 = ~n192 & n740;
  assign n742 = ~n192 & ~n741;
  assign n743 = ~n738 & n742;
  assign n744 = ~n737 & n743;
  assign \V119(19)  = n734 | ~n744;
  assign n746 = \V56(4)  & ~n203;
  assign n747 = ~n197 & n746;
  assign n748 = ~n192 & n747;
  assign n749 = \V56(8)  & n203;
  assign n750 = ~n197 & n749;
  assign n751 = ~n192 & n750;
  assign n752 = \V56(11)  & n345;
  assign n753 = n197 & n403;
  assign n754 = ~n192 & n753;
  assign n755 = ~n192 & ~n754;
  assign n756 = ~n752 & n755;
  assign n757 = ~n751 & n756;
  assign \V119(18)  = n748 | ~n757;
  assign n759 = \V56(18)  & ~n203;
  assign n760 = ~n197 & n759;
  assign n761 = ~n192 & n760;
  assign n762 = ~n197 & n492;
  assign n763 = ~n192 & n762;
  assign n764 = \V56(25)  & ~n203;
  assign n765 = n197 & n764;
  assign n766 = ~n192 & n765;
  assign n767 = n197 & n642;
  assign n768 = ~n192 & n767;
  assign n769 = n224 & ~n768;
  assign n770 = ~n766 & n769;
  assign n771 = ~n763 & n770;
  assign \V151(1)  = n761 | ~n771;
  assign n773 = \V56(17)  & ~n203;
  assign n774 = ~n197 & n773;
  assign n775 = ~n192 & n774;
  assign n776 = ~n197 & n506;
  assign n777 = ~n192 & n776;
  assign n778 = \V56(24)  & ~n203;
  assign n779 = n197 & n778;
  assign n780 = ~n192 & n779;
  assign n781 = n197 & n530;
  assign n782 = ~n192 & n781;
  assign n783 = n224 & ~n782;
  assign n784 = ~n780 & n783;
  assign n785 = ~n777 & n784;
  assign \V151(0)  = n775 | ~n785;
  assign n787 = \V24(11)  & ~n203;
  assign n788 = ~n197 & n787;
  assign n789 = ~n192 & n788;
  assign n790 = \V56(1)  & n203;
  assign n791 = ~n197 & n790;
  assign n792 = ~n192 & n791;
  assign n793 = \V56(4)  & n345;
  assign n794 = n197 & n544;
  assign n795 = ~n192 & n794;
  assign n796 = ~n192 & ~n795;
  assign n797 = ~n793 & n796;
  assign n798 = ~n792 & n797;
  assign \V119(11)  = n789 | ~n798;
  assign n800 = ~n197 & n778;
  assign n801 = ~n192 & n800;
  assign n802 = ~n197 & n347;
  assign n803 = ~n192 & n802;
  assign n804 = n197 & n719;
  assign n805 = ~n192 & n804;
  assign n806 = n197 & n474;
  assign n807 = ~n192 & n806;
  assign n808 = n224 & ~n807;
  assign n809 = ~n805 & n808;
  assign n810 = ~n803 & n809;
  assign \V151(7)  = n801 | ~n810;
  assign n812 = \V24(10)  & ~n203;
  assign n813 = ~n197 & n812;
  assign n814 = ~n192 & n813;
  assign n815 = \V56(3)  & n345;
  assign n816 = n197 & n488;
  assign n817 = ~n192 & n816;
  assign n818 = ~n192 & ~n817;
  assign n819 = ~n815 & n818;
  assign n820 = ~n328 & n819;
  assign \V119(10)  = n814 | ~n820;
  assign n822 = \V56(23)  & ~n203;
  assign n823 = ~n197 & n822;
  assign n824 = ~n192 & n823;
  assign n825 = ~n197 & n377;
  assign n826 = ~n192 & n825;
  assign n827 = n197 & n597;
  assign n828 = ~n192 & n827;
  assign n829 = n197 & n417;
  assign n830 = ~n192 & n829;
  assign n831 = n224 & ~n830;
  assign n832 = ~n828 & n831;
  assign n833 = ~n826 & n832;
  assign \V151(6)  = n824 | ~n833;
  assign n835 = \V24(13)  & ~n203;
  assign n836 = ~n197 & n835;
  assign n837 = ~n192 & n836;
  assign n838 = \V56(3)  & n203;
  assign n839 = ~n197 & n838;
  assign n840 = ~n192 & n839;
  assign n841 = \V56(6)  & n345;
  assign n842 = n197 & n614;
  assign n843 = ~n192 & n842;
  assign n844 = ~n192 & ~n843;
  assign n845 = ~n841 & n844;
  assign n846 = ~n840 & n845;
  assign \V119(13)  = n837 | ~n846;
  assign n848 = ~n197 & n630;
  assign n849 = ~n192 & n848;
  assign n850 = ~n197 & n407;
  assign n851 = ~n192 & n850;
  assign n852 = n197 & n442;
  assign n853 = ~n192 & n852;
  assign n854 = n197 & n295;
  assign n855 = ~n192 & n854;
  assign n856 = n224 & ~n855;
  assign n857 = ~n853 & n856;
  assign n858 = ~n851 & n857;
  assign \V151(9)  = n849 | ~n858;
  assign n860 = \V24(12)  & ~n203;
  assign n861 = ~n197 & n860;
  assign n862 = ~n192 & n861;
  assign n863 = \V56(2)  & n203;
  assign n864 = ~n197 & n863;
  assign n865 = ~n192 & n864;
  assign n866 = \V56(5)  & n345;
  assign n867 = n197 & n516;
  assign n868 = ~n192 & n867;
  assign n869 = ~n192 & ~n868;
  assign n870 = ~n866 & n869;
  assign n871 = ~n865 & n870;
  assign \V119(12)  = n862 | ~n871;
  assign n873 = ~n197 & n764;
  assign n874 = ~n192 & n873;
  assign n875 = ~n197 & n435;
  assign n876 = ~n192 & n875;
  assign n877 = n197 & n679;
  assign n878 = ~n192 & n877;
  assign n879 = n197 & n459;
  assign n880 = ~n192 & n879;
  assign n881 = n224 & ~n880;
  assign n882 = ~n878 & n881;
  assign n883 = ~n876 & n882;
  assign \V151(8)  = n874 | ~n883;
  assign n885 = \V56(1)  & ~n203;
  assign n886 = ~n197 & n885;
  assign n887 = ~n192 & n886;
  assign n888 = \V56(5)  & n203;
  assign n889 = ~n197 & n888;
  assign n890 = ~n192 & n889;
  assign n891 = \V56(8)  & n345;
  assign n892 = n197 & n373;
  assign n893 = ~n192 & n892;
  assign n894 = ~n192 & ~n893;
  assign n895 = ~n891 & n894;
  assign n896 = ~n890 & n895;
  assign \V119(15)  = n887 | ~n896;
  assign n898 = \V24(14)  & ~n203;
  assign n899 = ~n197 & n898;
  assign n900 = ~n192 & n899;
  assign n901 = \V56(4)  & n203;
  assign n902 = ~n197 & n901;
  assign n903 = ~n192 & n902;
  assign n904 = \V56(7)  & n345;
  assign n905 = n197 & n572;
  assign n906 = ~n192 & n905;
  assign n907 = ~n192 & ~n906;
  assign n908 = ~n904 & n907;
  assign n909 = ~n903 & n908;
  assign \V119(14)  = n900 | ~n909;
  assign n911 = ~n197 & n390;
  assign n912 = ~n192 & n911;
  assign n913 = ~n197 & n300;
  assign n914 = ~n192 & n913;
  assign n915 = \V88(23)  & ~n203;
  assign n916 = n197 & n915;
  assign n917 = ~n192 & n916;
  assign n918 = \V88(31)  & n203;
  assign n919 = n197 & n918;
  assign n920 = ~n192 & n919;
  assign n921 = n224 & ~n920;
  assign n922 = ~n917 & n921;
  assign n923 = ~n914 & n922;
  assign \V151(31)  = n912 | ~n923;
  assign n925 = ~n197 & n313;
  assign n926 = ~n192 & n925;
  assign n927 = ~n197 & n464;
  assign n928 = ~n192 & n927;
  assign n929 = \V88(22)  & ~n203;
  assign n930 = n197 & n929;
  assign n931 = ~n192 & n930;
  assign n932 = \V88(30)  & n203;
  assign n933 = n197 & n932;
  assign n934 = ~n192 & n933;
  assign n935 = n224 & ~n934;
  assign n936 = ~n931 & n935;
  assign n937 = ~n928 & n936;
  assign \V151(30)  = n926 | ~n937;
  assign n939 = \V56(16)  & ~n203;
  assign n940 = ~n197 & n939;
  assign n941 = ~n192 & n940;
  assign n942 = ~n197 & n739;
  assign n943 = ~n192 & n942;
  assign n944 = \V56(23)  & n345;
  assign n945 = n197 & n558;
  assign n946 = ~n192 & n945;
  assign n947 = ~n192 & ~n946;
  assign n948 = ~n944 & n947;
  assign n949 = ~n943 & n948;
  assign \V119(30)  = n941 | ~n949;
  assign n951 = \V24(3)  & ~n203;
  assign n952 = ~n197 & n951;
  assign n953 = ~n192 & n952;
  assign n954 = n197 & n901;
  assign n955 = ~n192 & n954;
  assign n956 = ~n192 & ~n955;
  assign n957 = ~n345 & n956;
  assign n958 = ~n684 & n957;
  assign \V119(3)  = n953 | ~n958;
  assign n960 = \V24(2)  & ~n203;
  assign n961 = ~n197 & n960;
  assign n962 = ~n192 & n961;
  assign n963 = n197 & n838;
  assign n964 = ~n192 & n963;
  assign n965 = ~n192 & ~n964;
  assign n966 = ~n345 & n965;
  assign n967 = ~n723 & n966;
  assign \V119(2)  = n962 | ~n967;
  assign n969 = \V24(5)  & ~n203;
  assign n970 = ~n197 & n969;
  assign n971 = ~n192 & n970;
  assign n972 = n197 & n696;
  assign n973 = ~n192 & n972;
  assign n974 = ~n192 & ~n973;
  assign n975 = ~n345 & n974;
  assign n976 = ~n419 & n975;
  assign \V119(5)  = n971 | ~n976;
  assign n978 = \V24(4)  & ~n203;
  assign n979 = ~n197 & n978;
  assign n980 = ~n192 & n979;
  assign n981 = n197 & n888;
  assign n982 = ~n192 & n981;
  assign n983 = ~n192 & ~n982;
  assign n984 = ~n345 & n983;
  assign n985 = ~n447 & n984;
  assign \V119(4)  = n980 | ~n985;
  assign n987 = \V24(1)  & ~n203;
  assign n988 = ~n197 & n987;
  assign n989 = ~n192 & n988;
  assign n990 = n197 & n863;
  assign n991 = ~n192 & n990;
  assign n992 = ~n192 & ~n991;
  assign n993 = ~n345 & n992;
  assign n994 = ~n602 & n993;
  assign \V119(1)  = n989 | ~n994;
  assign n996 = \V24(0)  & ~n203;
  assign n997 = ~n197 & n996;
  assign n998 = ~n192 & n997;
  assign n999 = n197 & n790;
  assign n1000 = ~n192 & n999;
  assign n1001 = ~n192 & ~n1000;
  assign n1002 = ~n345 & n1001;
  assign n1003 = ~n644 & n1002;
  assign \V119(0)  = n998 | ~n1003;
  assign n1005 = \V24(7)  & ~n203;
  assign n1006 = ~n197 & n1005;
  assign n1007 = ~n192 & n1006;
  assign n1008 = \V56(0)  & n345;
  assign n1009 = n197 & n749;
  assign n1010 = ~n192 & n1009;
  assign n1011 = ~n192 & ~n1010;
  assign n1012 = ~n1008 & n1011;
  assign n1013 = ~n461 & n1012;
  assign \V119(7)  = n1007 | ~n1013;
  assign n1015 = \V24(6)  & ~n203;
  assign n1016 = ~n197 & n1015;
  assign n1017 = ~n192 & n1016;
  assign n1018 = n197 & n656;
  assign n1019 = ~n192 & n1018;
  assign n1020 = ~n192 & ~n1019;
  assign n1021 = ~n345 & n1020;
  assign n1022 = ~n476 & n1021;
  assign \V119(6)  = n1017 | ~n1022;
  assign n1024 = \V24(9)  & ~n203;
  assign n1025 = ~n197 & n1024;
  assign n1026 = ~n192 & n1025;
  assign n1027 = \V56(2)  & n345;
  assign n1028 = n197 & n502;
  assign n1029 = ~n192 & n1028;
  assign n1030 = ~n192 & ~n1029;
  assign n1031 = ~n1027 & n1030;
  assign n1032 = ~n282 & n1031;
  assign \V119(9)  = n1026 | ~n1032;
  assign n1034 = \V24(8)  & ~n203;
  assign n1035 = ~n197 & n1034;
  assign n1036 = ~n192 & n1035;
  assign n1037 = \V56(1)  & n345;
  assign n1038 = n197 & n735;
  assign n1039 = ~n192 & n1038;
  assign n1040 = ~n192 & ~n1039;
  assign n1041 = ~n1037 & n1040;
  assign n1042 = ~n297 & n1041;
  assign \V119(8)  = n1036 | ~n1042;
endmodule


