// Benchmark "ksa_64" written by ABC on Sat Apr 23 20:18:05 2016

module ksa_64 ( 
    a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7, a8, b8,
    a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15, b15,
    a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22, b22,
    a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29, b29,
    a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36, b36,
    a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43, b43,
    a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50, b50,
    a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57, b57,
    a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64  );
  input  a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7,
    a8, b8, a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15,
    b15, a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22,
    b22, a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29,
    b29, a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36,
    b36, a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43,
    b43, a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50,
    b50, a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57,
    b57, a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64;
  wire n194, n195, n197, n198, n199, n200, n201, n203, n204, n205, n206,
    n207, n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n230, n231, n232, n233,
    n234, n235, n236, n237, n239, n240, n241, n242, n243, n244, n245, n246,
    n248, n249, n250, n251, n252, n253, n254, n255, n257, n258, n259, n260,
    n261, n262, n263, n264, n266, n267, n268, n269, n270, n271, n272, n273,
    n275, n276, n277, n278, n279, n280, n281, n282, n284, n285, n286, n287,
    n288, n289, n290, n291, n293, n294, n295, n296, n297, n298, n299, n300,
    n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314,
    n315, n316, n317, n318, n320, n321, n322, n323, n324, n325, n326, n327,
    n329, n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
    n342, n343, n344, n345, n347, n348, n349, n350, n351, n352, n353, n354,
    n356, n357, n358, n359, n360, n361, n362, n363, n365, n366, n367, n368,
    n369, n370, n371, n372, n374, n375, n376, n377, n378, n379, n380, n381,
    n383, n384, n385, n386, n387, n388, n389, n390, n392, n393, n394, n395,
    n396, n397, n398, n399, n401, n402, n403, n404, n405, n406, n407, n408,
    n410, n411, n412, n413, n414, n415, n416, n417, n419, n420, n421, n422,
    n423, n424, n425, n426, n428, n429, n430, n431, n432, n433, n434, n435,
    n437, n438, n439, n440, n441, n442, n443, n444, n446, n447, n448, n449,
    n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461, n462,
    n464, n465, n466, n467, n468, n469, n470, n471, n473, n474, n475, n476,
    n477, n478, n479, n480, n482, n483, n484, n485, n486, n487, n488, n489,
    n491, n492, n493, n494, n495, n496, n497, n498, n500, n501, n502, n503,
    n504, n505, n506, n507, n509, n510, n511, n512, n513, n514, n515, n516,
    n518, n519, n520, n521, n522, n523, n524, n525, n527, n528, n529, n530,
    n531, n532, n533, n534, n536, n537, n538, n539, n540, n541, n542, n543,
    n545, n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557,
    n558, n559, n560, n561, n563, n564, n565, n566, n567, n568, n569, n570,
    n572, n573, n574, n575, n576, n577, n578, n579, n581, n582, n583, n584,
    n585, n586, n587, n588, n590, n591, n592, n593, n594, n595, n596, n597,
    n599, n600, n601, n602, n603, n604, n605, n606, n608, n609, n610, n611,
    n612, n613, n614, n615, n617, n618, n619, n620, n621, n622, n623, n624,
    n626, n627, n628, n629, n630, n631, n632, n633, n635, n636, n637, n638,
    n639, n640, n641, n642, n644, n645, n646, n647, n648, n649, n650, n651,
    n653, n654, n655, n656, n657, n658, n659, n660, n662, n663, n664, n665,
    n666, n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n678,
    n680, n681, n682, n683, n684, n685, n686, n687, n689, n690, n691, n692,
    n693, n694, n695, n696, n698, n699, n700, n701, n702, n703, n704, n705,
    n707, n708, n709, n710, n711, n712, n713, n714, n716, n717, n718, n719,
    n720, n721, n722, n723, n725, n726, n727, n728, n729, n730, n731, n732,
    n734, n735, n736, n737, n738, n739, n740, n741, n743, n744, n745, n746,
    n747, n748, n749, n750, n752, n753, n754, n755, n756, n757, n758, n759,
    n761, n762;
  assign n194 = a0 & b0;
  assign n195 = ~a0 & ~b0;
  assign s0 = ~n194 & ~n195;
  assign n197 = a1 & b1;
  assign n198 = ~a1 & ~b1;
  assign n199 = ~n197 & ~n198;
  assign n200 = n194 & n199;
  assign n201 = ~n194 & ~n199;
  assign s1 = ~n200 & ~n201;
  assign n203 = ~n197 & ~n200;
  assign n204 = a2 & b2;
  assign n205 = ~a2 & ~b2;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n203 & n206;
  assign n208 = n203 & ~n206;
  assign s2 = ~n207 & ~n208;
  assign n210 = n200 & n206;
  assign n211 = ~n197 & ~n204;
  assign n212 = ~n205 & ~n211;
  assign n213 = ~n210 & ~n212;
  assign n214 = a3 & b3;
  assign n215 = ~a3 & ~b3;
  assign n216 = ~n214 & ~n215;
  assign n217 = n213 & ~n216;
  assign n218 = ~n213 & n216;
  assign s3 = ~n217 & ~n218;
  assign n220 = n207 & n216;
  assign n221 = ~n204 & ~n214;
  assign n222 = ~n215 & ~n221;
  assign n223 = ~n220 & ~n222;
  assign n224 = a4 & b4;
  assign n225 = ~a4 & ~b4;
  assign n226 = ~n224 & ~n225;
  assign n227 = n223 & ~n226;
  assign n228 = ~n223 & n226;
  assign s4 = ~n227 & ~n228;
  assign n230 = a5 & b5;
  assign n231 = ~a5 & ~b5;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n214 & ~n224;
  assign n234 = ~n218 & n233;
  assign n235 = ~n225 & ~n234;
  assign n236 = ~n232 & ~n235;
  assign n237 = n232 & n235;
  assign s5 = ~n236 & ~n237;
  assign n239 = a6 & b6;
  assign n240 = ~a6 & ~b6;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~n224 & ~n230;
  assign n243 = ~n228 & n242;
  assign n244 = ~n231 & ~n243;
  assign n245 = ~n241 & ~n244;
  assign n246 = n241 & n244;
  assign s6 = ~n245 & ~n246;
  assign n248 = a7 & b7;
  assign n249 = ~a7 & ~b7;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n230 & ~n239;
  assign n252 = ~n237 & n251;
  assign n253 = ~n240 & ~n252;
  assign n254 = ~n250 & ~n253;
  assign n255 = n250 & n253;
  assign s7 = ~n254 & ~n255;
  assign n257 = a8 & b8;
  assign n258 = ~a8 & ~b8;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~n239 & ~n248;
  assign n261 = ~n246 & n260;
  assign n262 = ~n249 & ~n261;
  assign n263 = n259 & n262;
  assign n264 = ~n259 & ~n262;
  assign s8 = ~n263 & ~n264;
  assign n266 = a9 & b9;
  assign n267 = ~a9 & ~b9;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~n248 & ~n257;
  assign n270 = ~n255 & n269;
  assign n271 = ~n258 & ~n270;
  assign n272 = ~n268 & ~n271;
  assign n273 = n268 & n271;
  assign s9 = ~n272 & ~n273;
  assign n275 = a10 & b10;
  assign n276 = ~a10 & ~b10;
  assign n277 = ~n275 & ~n276;
  assign n278 = ~n257 & ~n266;
  assign n279 = ~n263 & n278;
  assign n280 = ~n267 & ~n279;
  assign n281 = ~n277 & ~n280;
  assign n282 = n277 & n280;
  assign s10 = ~n281 & ~n282;
  assign n284 = a11 & b11;
  assign n285 = ~a11 & ~b11;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~n266 & ~n275;
  assign n288 = ~n273 & n287;
  assign n289 = ~n276 & ~n288;
  assign n290 = n286 & n289;
  assign n291 = ~n286 & ~n289;
  assign s11 = ~n290 & ~n291;
  assign n293 = a12 & b12;
  assign n294 = ~a12 & ~b12;
  assign n295 = ~n293 & ~n294;
  assign n296 = ~n275 & ~n284;
  assign n297 = ~n282 & n296;
  assign n298 = ~n285 & ~n297;
  assign n299 = n295 & n298;
  assign n300 = ~n295 & ~n298;
  assign s12 = ~n299 & ~n300;
  assign n302 = a13 & b13;
  assign n303 = ~a13 & ~b13;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~n284 & ~n293;
  assign n306 = ~n290 & n305;
  assign n307 = ~n294 & ~n306;
  assign n308 = ~n304 & ~n307;
  assign n309 = n304 & n307;
  assign s13 = ~n308 & ~n309;
  assign n311 = a14 & b14;
  assign n312 = ~a14 & ~b14;
  assign n313 = ~n311 & ~n312;
  assign n314 = ~n293 & ~n302;
  assign n315 = ~n299 & n314;
  assign n316 = ~n303 & ~n315;
  assign n317 = ~n313 & ~n316;
  assign n318 = n313 & n316;
  assign s14 = ~n317 & ~n318;
  assign n320 = a15 & b15;
  assign n321 = ~a15 & ~b15;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n302 & ~n311;
  assign n324 = ~n309 & n323;
  assign n325 = ~n312 & ~n324;
  assign n326 = n322 & n325;
  assign n327 = ~n322 & ~n325;
  assign s15 = ~n326 & ~n327;
  assign n329 = a16 & b16;
  assign n330 = ~a16 & ~b16;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n311 & ~n320;
  assign n333 = ~n318 & n332;
  assign n334 = ~n321 & ~n333;
  assign n335 = n331 & n334;
  assign n336 = ~n331 & ~n334;
  assign s16 = ~n335 & ~n336;
  assign n338 = a17 & b17;
  assign n339 = ~a17 & ~b17;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~n320 & ~n329;
  assign n342 = ~n326 & n341;
  assign n343 = ~n330 & ~n342;
  assign n344 = ~n340 & ~n343;
  assign n345 = n340 & n343;
  assign s17 = ~n344 & ~n345;
  assign n347 = a18 & b18;
  assign n348 = ~a18 & ~b18;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~n329 & ~n338;
  assign n351 = ~n335 & n350;
  assign n352 = ~n339 & ~n351;
  assign n353 = n349 & n352;
  assign n354 = ~n349 & ~n352;
  assign s18 = ~n353 & ~n354;
  assign n356 = a19 & b19;
  assign n357 = ~a19 & ~b19;
  assign n358 = ~n356 & ~n357;
  assign n359 = ~n338 & ~n347;
  assign n360 = ~n345 & n359;
  assign n361 = ~n348 & ~n360;
  assign n362 = n358 & n361;
  assign n363 = ~n358 & ~n361;
  assign s19 = ~n362 & ~n363;
  assign n365 = a20 & b20;
  assign n366 = ~a20 & ~b20;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~n347 & ~n356;
  assign n369 = ~n353 & n368;
  assign n370 = ~n357 & ~n369;
  assign n371 = ~n367 & ~n370;
  assign n372 = n367 & n370;
  assign s20 = ~n371 & ~n372;
  assign n374 = a21 & b21;
  assign n375 = ~a21 & ~b21;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n356 & ~n365;
  assign n378 = ~n362 & n377;
  assign n379 = ~n366 & ~n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = n376 & n379;
  assign s21 = ~n380 & ~n381;
  assign n383 = a22 & b22;
  assign n384 = ~a22 & ~b22;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n365 & ~n374;
  assign n387 = ~n372 & n386;
  assign n388 = ~n375 & ~n387;
  assign n389 = n385 & n388;
  assign n390 = ~n385 & ~n388;
  assign s22 = ~n389 & ~n390;
  assign n392 = a23 & b23;
  assign n393 = ~a23 & ~b23;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n374 & ~n383;
  assign n396 = ~n381 & n395;
  assign n397 = ~n384 & ~n396;
  assign n398 = ~n394 & ~n397;
  assign n399 = n394 & n397;
  assign s23 = ~n398 & ~n399;
  assign n401 = a24 & b24;
  assign n402 = ~a24 & ~b24;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n383 & ~n392;
  assign n405 = ~n389 & n404;
  assign n406 = ~n393 & ~n405;
  assign n407 = ~n403 & ~n406;
  assign n408 = n403 & n406;
  assign s24 = ~n407 & ~n408;
  assign n410 = a25 & b25;
  assign n411 = ~a25 & ~b25;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n392 & ~n401;
  assign n414 = ~n399 & n413;
  assign n415 = ~n402 & ~n414;
  assign n416 = ~n412 & ~n415;
  assign n417 = n412 & n415;
  assign s25 = ~n416 & ~n417;
  assign n419 = a26 & b26;
  assign n420 = ~a26 & ~b26;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n401 & ~n410;
  assign n423 = ~n408 & n422;
  assign n424 = ~n411 & ~n423;
  assign n425 = ~n421 & ~n424;
  assign n426 = n421 & n424;
  assign s26 = ~n425 & ~n426;
  assign n428 = a27 & b27;
  assign n429 = ~a27 & ~b27;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~n410 & ~n419;
  assign n432 = ~n417 & n431;
  assign n433 = ~n420 & ~n432;
  assign n434 = ~n430 & ~n433;
  assign n435 = n430 & n433;
  assign s27 = ~n434 & ~n435;
  assign n437 = a28 & b28;
  assign n438 = ~a28 & ~b28;
  assign n439 = ~n437 & ~n438;
  assign n440 = ~n419 & ~n428;
  assign n441 = ~n426 & n440;
  assign n442 = ~n429 & ~n441;
  assign n443 = n439 & n442;
  assign n444 = ~n439 & ~n442;
  assign s28 = ~n443 & ~n444;
  assign n446 = a29 & b29;
  assign n447 = ~a29 & ~b29;
  assign n448 = ~n446 & ~n447;
  assign n449 = ~n428 & ~n437;
  assign n450 = ~n435 & n449;
  assign n451 = ~n438 & ~n450;
  assign n452 = n448 & n451;
  assign n453 = ~n448 & ~n451;
  assign s29 = ~n452 & ~n453;
  assign n455 = a30 & b30;
  assign n456 = ~a30 & ~b30;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n437 & ~n446;
  assign n459 = ~n443 & n458;
  assign n460 = ~n447 & ~n459;
  assign n461 = ~n457 & ~n460;
  assign n462 = n457 & n460;
  assign s30 = ~n461 & ~n462;
  assign n464 = a31 & b31;
  assign n465 = ~a31 & ~b31;
  assign n466 = ~n464 & ~n465;
  assign n467 = ~n446 & ~n455;
  assign n468 = ~n452 & n467;
  assign n469 = ~n456 & ~n468;
  assign n470 = ~n466 & ~n469;
  assign n471 = n466 & n469;
  assign s31 = ~n470 & ~n471;
  assign n473 = a32 & b32;
  assign n474 = ~a32 & ~b32;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n455 & ~n464;
  assign n477 = ~n462 & n476;
  assign n478 = ~n465 & ~n477;
  assign n479 = ~n475 & ~n478;
  assign n480 = n475 & n478;
  assign s32 = ~n479 & ~n480;
  assign n482 = a33 & b33;
  assign n483 = ~a33 & ~b33;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n464 & ~n473;
  assign n486 = ~n471 & n485;
  assign n487 = ~n474 & ~n486;
  assign n488 = ~n484 & ~n487;
  assign n489 = n484 & n487;
  assign s33 = ~n488 & ~n489;
  assign n491 = a34 & b34;
  assign n492 = ~a34 & ~b34;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n473 & ~n482;
  assign n495 = ~n480 & n494;
  assign n496 = ~n483 & ~n495;
  assign n497 = n493 & n496;
  assign n498 = ~n493 & ~n496;
  assign s34 = ~n497 & ~n498;
  assign n500 = a35 & b35;
  assign n501 = ~a35 & ~b35;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~n482 & ~n491;
  assign n504 = ~n489 & n503;
  assign n505 = ~n492 & ~n504;
  assign n506 = ~n502 & ~n505;
  assign n507 = n502 & n505;
  assign s35 = ~n506 & ~n507;
  assign n509 = a36 & b36;
  assign n510 = ~a36 & ~b36;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~n491 & ~n500;
  assign n513 = ~n497 & n512;
  assign n514 = ~n501 & ~n513;
  assign n515 = ~n511 & ~n514;
  assign n516 = n511 & n514;
  assign s36 = ~n515 & ~n516;
  assign n518 = a37 & b37;
  assign n519 = ~a37 & ~b37;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n500 & ~n509;
  assign n522 = ~n507 & n521;
  assign n523 = ~n510 & ~n522;
  assign n524 = ~n520 & ~n523;
  assign n525 = n520 & n523;
  assign s37 = ~n524 & ~n525;
  assign n527 = a38 & b38;
  assign n528 = ~a38 & ~b38;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~n509 & ~n518;
  assign n531 = ~n516 & n530;
  assign n532 = ~n519 & ~n531;
  assign n533 = ~n529 & ~n532;
  assign n534 = n529 & n532;
  assign s38 = ~n533 & ~n534;
  assign n536 = a39 & b39;
  assign n537 = ~a39 & ~b39;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n518 & ~n527;
  assign n540 = ~n525 & n539;
  assign n541 = ~n528 & ~n540;
  assign n542 = ~n538 & ~n541;
  assign n543 = n538 & n541;
  assign s39 = ~n542 & ~n543;
  assign n545 = a40 & b40;
  assign n546 = ~a40 & ~b40;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n527 & ~n536;
  assign n549 = ~n534 & n548;
  assign n550 = ~n537 & ~n549;
  assign n551 = ~n547 & ~n550;
  assign n552 = n547 & n550;
  assign s40 = ~n551 & ~n552;
  assign n554 = a41 & b41;
  assign n555 = ~a41 & ~b41;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n536 & ~n545;
  assign n558 = ~n543 & n557;
  assign n559 = ~n546 & ~n558;
  assign n560 = ~n556 & ~n559;
  assign n561 = n556 & n559;
  assign s41 = ~n560 & ~n561;
  assign n563 = a42 & b42;
  assign n564 = ~a42 & ~b42;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n545 & ~n554;
  assign n567 = ~n552 & n566;
  assign n568 = ~n555 & ~n567;
  assign n569 = ~n565 & ~n568;
  assign n570 = n565 & n568;
  assign s42 = ~n569 & ~n570;
  assign n572 = a43 & b43;
  assign n573 = ~a43 & ~b43;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n554 & ~n563;
  assign n576 = ~n561 & n575;
  assign n577 = ~n564 & ~n576;
  assign n578 = ~n574 & ~n577;
  assign n579 = n574 & n577;
  assign s43 = ~n578 & ~n579;
  assign n581 = a44 & b44;
  assign n582 = ~a44 & ~b44;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n563 & ~n572;
  assign n585 = ~n570 & n584;
  assign n586 = ~n573 & ~n585;
  assign n587 = ~n583 & ~n586;
  assign n588 = n583 & n586;
  assign s44 = ~n587 & ~n588;
  assign n590 = a45 & b45;
  assign n591 = ~a45 & ~b45;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n572 & ~n581;
  assign n594 = ~n579 & n593;
  assign n595 = ~n582 & ~n594;
  assign n596 = ~n592 & ~n595;
  assign n597 = n592 & n595;
  assign s45 = ~n596 & ~n597;
  assign n599 = a46 & b46;
  assign n600 = ~a46 & ~b46;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n581 & ~n590;
  assign n603 = ~n588 & n602;
  assign n604 = ~n591 & ~n603;
  assign n605 = ~n601 & ~n604;
  assign n606 = n601 & n604;
  assign s46 = ~n605 & ~n606;
  assign n608 = a47 & b47;
  assign n609 = ~a47 & ~b47;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~n590 & ~n599;
  assign n612 = ~n597 & n611;
  assign n613 = ~n600 & ~n612;
  assign n614 = ~n610 & ~n613;
  assign n615 = n610 & n613;
  assign s47 = ~n614 & ~n615;
  assign n617 = a48 & b48;
  assign n618 = ~a48 & ~b48;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n599 & ~n608;
  assign n621 = ~n606 & n620;
  assign n622 = ~n609 & ~n621;
  assign n623 = ~n619 & ~n622;
  assign n624 = n619 & n622;
  assign s48 = ~n623 & ~n624;
  assign n626 = a49 & b49;
  assign n627 = ~a49 & ~b49;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~n608 & ~n617;
  assign n630 = ~n615 & n629;
  assign n631 = ~n618 & ~n630;
  assign n632 = ~n628 & ~n631;
  assign n633 = n628 & n631;
  assign s49 = ~n632 & ~n633;
  assign n635 = a50 & b50;
  assign n636 = ~a50 & ~b50;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n617 & ~n626;
  assign n639 = ~n624 & n638;
  assign n640 = ~n627 & ~n639;
  assign n641 = ~n637 & ~n640;
  assign n642 = n637 & n640;
  assign s50 = ~n641 & ~n642;
  assign n644 = a51 & b51;
  assign n645 = ~a51 & ~b51;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~n626 & ~n635;
  assign n648 = ~n633 & n647;
  assign n649 = ~n636 & ~n648;
  assign n650 = ~n646 & ~n649;
  assign n651 = n646 & n649;
  assign s51 = ~n650 & ~n651;
  assign n653 = a52 & b52;
  assign n654 = ~a52 & ~b52;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n635 & ~n644;
  assign n657 = ~n642 & n656;
  assign n658 = ~n645 & ~n657;
  assign n659 = ~n655 & ~n658;
  assign n660 = n655 & n658;
  assign s52 = ~n659 & ~n660;
  assign n662 = a53 & b53;
  assign n663 = ~a53 & ~b53;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n644 & ~n653;
  assign n666 = ~n651 & n665;
  assign n667 = ~n654 & ~n666;
  assign n668 = ~n664 & ~n667;
  assign n669 = n664 & n667;
  assign s53 = ~n668 & ~n669;
  assign n671 = a54 & b54;
  assign n672 = ~a54 & ~b54;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n653 & ~n662;
  assign n675 = ~n660 & n674;
  assign n676 = ~n663 & ~n675;
  assign n677 = ~n673 & ~n676;
  assign n678 = n673 & n676;
  assign s54 = ~n677 & ~n678;
  assign n680 = a55 & b55;
  assign n681 = ~a55 & ~b55;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~n662 & ~n671;
  assign n684 = ~n669 & n683;
  assign n685 = ~n672 & ~n684;
  assign n686 = ~n682 & ~n685;
  assign n687 = n682 & n685;
  assign s55 = ~n686 & ~n687;
  assign n689 = a56 & b56;
  assign n690 = ~a56 & ~b56;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~n671 & ~n680;
  assign n693 = ~n678 & n692;
  assign n694 = ~n681 & ~n693;
  assign n695 = ~n691 & ~n694;
  assign n696 = n691 & n694;
  assign s56 = ~n695 & ~n696;
  assign n698 = a57 & b57;
  assign n699 = ~a57 & ~b57;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~n680 & ~n689;
  assign n702 = ~n687 & n701;
  assign n703 = ~n690 & ~n702;
  assign n704 = n700 & n703;
  assign n705 = ~n700 & ~n703;
  assign s57 = ~n704 & ~n705;
  assign n707 = a58 & b58;
  assign n708 = ~a58 & ~b58;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n689 & ~n698;
  assign n711 = ~n696 & n710;
  assign n712 = ~n699 & ~n711;
  assign n713 = n709 & n712;
  assign n714 = ~n709 & ~n712;
  assign s58 = ~n713 & ~n714;
  assign n716 = a59 & b59;
  assign n717 = ~a59 & ~b59;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n698 & ~n707;
  assign n720 = ~n704 & n719;
  assign n721 = ~n708 & ~n720;
  assign n722 = n718 & n721;
  assign n723 = ~n718 & ~n721;
  assign s59 = ~n722 & ~n723;
  assign n725 = a60 & b60;
  assign n726 = ~a60 & ~b60;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n707 & ~n716;
  assign n729 = ~n713 & n728;
  assign n730 = ~n717 & ~n729;
  assign n731 = n727 & n730;
  assign n732 = ~n727 & ~n730;
  assign s60 = ~n731 & ~n732;
  assign n734 = a61 & b61;
  assign n735 = ~a61 & ~b61;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~n716 & ~n725;
  assign n738 = ~n722 & n737;
  assign n739 = ~n726 & ~n738;
  assign n740 = n736 & n739;
  assign n741 = ~n736 & ~n739;
  assign s61 = ~n740 & ~n741;
  assign n743 = a62 & b62;
  assign n744 = ~a62 & ~b62;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n725 & ~n734;
  assign n747 = ~n731 & n746;
  assign n748 = ~n735 & ~n747;
  assign n749 = ~n745 & ~n748;
  assign n750 = n745 & n748;
  assign s62 = ~n749 & ~n750;
  assign n752 = a63 & b63;
  assign n753 = ~a63 & ~b63;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n734 & ~n743;
  assign n756 = ~n740 & n755;
  assign n757 = ~n744 & ~n756;
  assign n758 = ~n754 & n757;
  assign n759 = n754 & ~n757;
  assign s63 = n758 | n759;
  assign n761 = ~n743 & ~n752;
  assign n762 = ~n750 & n761;
  assign s64 = ~n753 & ~n762;
endmodule


