// Benchmark "moa_12x8" written by ABC on Sat Apr 23 20:18:06 2016

module moa_12x8 ( 
    a0_0, a1_0, a2_0, a3_0, a4_0, a5_0, a6_0, a7_0, a0_1, a1_1, a2_1, a3_1,
    a4_1, a5_1, a6_1, a7_1, a0_2, a1_2, a2_2, a3_2, a4_2, a5_2, a6_2, a7_2,
    a0_3, a1_3, a2_3, a3_3, a4_3, a5_3, a6_3, a7_3, a0_4, a1_4, a2_4, a3_4,
    a4_4, a5_4, a6_4, a7_4, a0_5, a1_5, a2_5, a3_5, a4_5, a5_5, a6_5, a7_5,
    a0_6, a1_6, a2_6, a3_6, a4_6, a5_6, a6_6, a7_6, a0_7, a1_7, a2_7, a3_7,
    a4_7, a5_7, a6_7, a7_7, a0_8, a1_8, a2_8, a3_8, a4_8, a5_8, a6_8, a7_8,
    a0_9, a1_9, a2_9, a3_9, a4_9, a5_9, a6_9, a7_9, a0_10, a1_10, a2_10,
    a3_10, a4_10, a5_10, a6_10, a7_10, a0_11, a1_11, a2_11, a3_11, a4_11,
    a5_11, a6_11, a7_11,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12  );
  input  a0_0, a1_0, a2_0, a3_0, a4_0, a5_0, a6_0, a7_0, a0_1, a1_1,
    a2_1, a3_1, a4_1, a5_1, a6_1, a7_1, a0_2, a1_2, a2_2, a3_2, a4_2, a5_2,
    a6_2, a7_2, a0_3, a1_3, a2_3, a3_3, a4_3, a5_3, a6_3, a7_3, a0_4, a1_4,
    a2_4, a3_4, a4_4, a5_4, a6_4, a7_4, a0_5, a1_5, a2_5, a3_5, a4_5, a5_5,
    a6_5, a7_5, a0_6, a1_6, a2_6, a3_6, a4_6, a5_6, a6_6, a7_6, a0_7, a1_7,
    a2_7, a3_7, a4_7, a5_7, a6_7, a7_7, a0_8, a1_8, a2_8, a3_8, a4_8, a5_8,
    a6_8, a7_8, a0_9, a1_9, a2_9, a3_9, a4_9, a5_9, a6_9, a7_9, a0_10,
    a1_10, a2_10, a3_10, a4_10, a5_10, a6_10, a7_10, a0_11, a1_11, a2_11,
    a3_11, a4_11, a5_11, a6_11, a7_11;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12;
  wire n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n775, n776;
  assign n110 = a0_0 & a0_1;
  assign n111 = ~a0_0 & ~a0_1;
  assign n112 = ~n110 & ~n111;
  assign n113 = a0_2 & n112;
  assign n114 = ~a0_2 & ~n112;
  assign n115 = ~n113 & ~n114;
  assign n116 = a0_3 & a0_4;
  assign n117 = ~a0_3 & ~a0_4;
  assign n118 = ~n116 & ~n117;
  assign n119 = a0_5 & n118;
  assign n120 = ~a0_5 & ~n118;
  assign n121 = ~n119 & ~n120;
  assign n122 = n115 & n121;
  assign n123 = ~n115 & ~n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = a0_6 & a0_7;
  assign n126 = ~a0_6 & ~a0_7;
  assign n127 = ~n125 & ~n126;
  assign n128 = a0_8 & n127;
  assign n129 = ~a0_8 & ~n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = a0_9 & a0_10;
  assign n132 = ~a0_9 & ~a0_10;
  assign n133 = ~n131 & ~n132;
  assign n134 = a0_11 & n133;
  assign n135 = ~a0_11 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = n130 & n136;
  assign n138 = ~n130 & ~n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = n124 & n139;
  assign n141 = ~n124 & ~n139;
  assign s0 = ~n140 & ~n141;
  assign n143 = a1_6 & a1_7;
  assign n144 = ~a1_6 & ~a1_7;
  assign n145 = ~n143 & ~n144;
  assign n146 = a1_8 & n145;
  assign n147 = ~a1_8 & ~n145;
  assign n148 = ~n146 & ~n147;
  assign n149 = a1_9 & a1_10;
  assign n150 = ~a1_9 & ~a1_10;
  assign n151 = ~n149 & ~n150;
  assign n152 = a1_11 & n151;
  assign n153 = ~a1_11 & ~n151;
  assign n154 = ~n152 & ~n153;
  assign n155 = n148 & n154;
  assign n156 = ~n148 & ~n154;
  assign n157 = ~n155 & ~n156;
  assign n158 = a1_0 & a1_1;
  assign n159 = ~a1_0 & ~a1_1;
  assign n160 = ~n158 & ~n159;
  assign n161 = a1_2 & n160;
  assign n162 = ~a1_2 & ~n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = a1_3 & a1_4;
  assign n165 = ~a1_3 & ~a1_4;
  assign n166 = ~n164 & ~n165;
  assign n167 = a1_5 & n166;
  assign n168 = ~a1_5 & ~n166;
  assign n169 = ~n167 & ~n168;
  assign n170 = n163 & n169;
  assign n171 = ~n163 & ~n169;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~n110 & ~n113;
  assign n174 = ~n116 & ~n119;
  assign n175 = ~n173 & ~n174;
  assign n176 = n173 & n174;
  assign n177 = ~n175 & ~n176;
  assign n178 = n122 & n177;
  assign n179 = ~n122 & ~n177;
  assign n180 = ~n178 & ~n179;
  assign n181 = ~n125 & ~n128;
  assign n182 = ~n131 & ~n134;
  assign n183 = ~n181 & ~n182;
  assign n184 = n181 & n182;
  assign n185 = ~n183 & ~n184;
  assign n186 = n137 & n185;
  assign n187 = ~n137 & ~n185;
  assign n188 = ~n186 & ~n187;
  assign n189 = n180 & n188;
  assign n190 = ~n180 & ~n188;
  assign n191 = ~n189 & ~n190;
  assign n192 = n172 & n191;
  assign n193 = ~n172 & ~n191;
  assign n194 = ~n192 & ~n193;
  assign n195 = n157 & n194;
  assign n196 = ~n157 & ~n194;
  assign n197 = ~n195 & ~n196;
  assign n198 = n140 & n197;
  assign n199 = ~n140 & ~n197;
  assign s1 = ~n198 & ~n199;
  assign n201 = ~n195 & ~n198;
  assign n202 = ~n189 & ~n192;
  assign n203 = a2_6 & a2_7;
  assign n204 = ~a2_6 & ~a2_7;
  assign n205 = ~n203 & ~n204;
  assign n206 = a2_8 & n205;
  assign n207 = ~a2_8 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = a2_9 & a2_10;
  assign n210 = ~a2_9 & ~a2_10;
  assign n211 = ~n209 & ~n210;
  assign n212 = a2_11 & n211;
  assign n213 = ~a2_11 & ~n211;
  assign n214 = ~n212 & ~n213;
  assign n215 = n208 & n214;
  assign n216 = ~n208 & ~n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~n143 & ~n146;
  assign n219 = ~n149 & ~n152;
  assign n220 = ~n218 & ~n219;
  assign n221 = n218 & n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = n155 & n222;
  assign n224 = ~n155 & ~n222;
  assign n225 = ~n223 & ~n224;
  assign n226 = a2_0 & a2_1;
  assign n227 = ~a2_0 & ~a2_1;
  assign n228 = ~n226 & ~n227;
  assign n229 = a2_2 & n228;
  assign n230 = ~a2_2 & ~n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = a2_3 & a2_4;
  assign n233 = ~a2_3 & ~a2_4;
  assign n234 = ~n232 & ~n233;
  assign n235 = a2_5 & n234;
  assign n236 = ~a2_5 & ~n234;
  assign n237 = ~n235 & ~n236;
  assign n238 = n231 & n237;
  assign n239 = ~n231 & ~n237;
  assign n240 = ~n238 & ~n239;
  assign n241 = n225 & n240;
  assign n242 = ~n225 & ~n240;
  assign n243 = ~n241 & ~n242;
  assign n244 = n217 & n243;
  assign n245 = ~n217 & ~n243;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~n158 & ~n161;
  assign n248 = ~n164 & ~n167;
  assign n249 = ~n247 & ~n248;
  assign n250 = n247 & n248;
  assign n251 = ~n249 & ~n250;
  assign n252 = n170 & n251;
  assign n253 = ~n170 & ~n251;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~n175 & ~n178;
  assign n256 = ~n183 & ~n186;
  assign n257 = ~n255 & ~n256;
  assign n258 = n255 & n256;
  assign n259 = ~n257 & ~n258;
  assign n260 = n254 & n259;
  assign n261 = ~n254 & ~n259;
  assign n262 = ~n260 & ~n261;
  assign n263 = n246 & n262;
  assign n264 = ~n246 & ~n262;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n202 & n265;
  assign n267 = n202 & ~n265;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~n201 & n268;
  assign n270 = n201 & ~n268;
  assign s2 = ~n269 & ~n270;
  assign n272 = ~n266 & ~n269;
  assign n273 = a3_6 & a3_7;
  assign n274 = ~a3_6 & ~a3_7;
  assign n275 = ~n273 & ~n274;
  assign n276 = a3_8 & n275;
  assign n277 = ~a3_8 & ~n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = a3_9 & a3_10;
  assign n280 = ~a3_9 & ~a3_10;
  assign n281 = ~n279 & ~n280;
  assign n282 = a3_11 & n281;
  assign n283 = ~a3_11 & ~n281;
  assign n284 = ~n282 & ~n283;
  assign n285 = n278 & n284;
  assign n286 = ~n278 & ~n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~n203 & ~n206;
  assign n289 = ~n209 & ~n212;
  assign n290 = ~n288 & ~n289;
  assign n291 = n288 & n289;
  assign n292 = ~n290 & ~n291;
  assign n293 = n215 & n292;
  assign n294 = ~n215 & ~n292;
  assign n295 = ~n293 & ~n294;
  assign n296 = a3_0 & a3_1;
  assign n297 = ~a3_0 & ~a3_1;
  assign n298 = ~n296 & ~n297;
  assign n299 = a3_2 & n298;
  assign n300 = ~a3_2 & ~n298;
  assign n301 = ~n299 & ~n300;
  assign n302 = a3_3 & a3_4;
  assign n303 = ~a3_3 & ~a3_4;
  assign n304 = ~n302 & ~n303;
  assign n305 = a3_5 & n304;
  assign n306 = ~a3_5 & ~n304;
  assign n307 = ~n305 & ~n306;
  assign n308 = n301 & n307;
  assign n309 = ~n301 & ~n307;
  assign n310 = ~n308 & ~n309;
  assign n311 = n295 & n310;
  assign n312 = ~n295 & ~n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = n287 & n313;
  assign n315 = ~n287 & ~n313;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~n226 & ~n229;
  assign n318 = ~n232 & ~n235;
  assign n319 = ~n317 & ~n318;
  assign n320 = n317 & n318;
  assign n321 = ~n319 & ~n320;
  assign n322 = n238 & n321;
  assign n323 = ~n238 & ~n321;
  assign n324 = ~n322 & ~n323;
  assign n325 = ~n249 & ~n252;
  assign n326 = ~n220 & ~n223;
  assign n327 = ~n325 & ~n326;
  assign n328 = n325 & n326;
  assign n329 = ~n327 & ~n328;
  assign n330 = n324 & n329;
  assign n331 = ~n324 & ~n329;
  assign n332 = ~n330 & ~n331;
  assign n333 = n316 & n332;
  assign n334 = ~n316 & ~n332;
  assign n335 = ~n333 & ~n334;
  assign n336 = ~n257 & ~n260;
  assign n337 = ~n241 & ~n244;
  assign n338 = ~n336 & ~n337;
  assign n339 = n336 & n337;
  assign n340 = ~n338 & ~n339;
  assign n341 = n263 & n340;
  assign n342 = ~n263 & ~n340;
  assign n343 = ~n341 & ~n342;
  assign n344 = n335 & n343;
  assign n345 = ~n335 & ~n343;
  assign n346 = ~n344 & ~n345;
  assign n347 = ~n272 & n346;
  assign n348 = n272 & ~n346;
  assign s3 = ~n347 & ~n348;
  assign n350 = ~n344 & ~n347;
  assign n351 = a4_6 & a4_7;
  assign n352 = ~a4_6 & ~a4_7;
  assign n353 = ~n351 & ~n352;
  assign n354 = a4_8 & n353;
  assign n355 = ~a4_8 & ~n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = a4_9 & a4_10;
  assign n358 = ~a4_9 & ~a4_10;
  assign n359 = ~n357 & ~n358;
  assign n360 = a4_11 & n359;
  assign n361 = ~a4_11 & ~n359;
  assign n362 = ~n360 & ~n361;
  assign n363 = n356 & n362;
  assign n364 = ~n356 & ~n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n273 & ~n276;
  assign n367 = ~n279 & ~n282;
  assign n368 = ~n366 & ~n367;
  assign n369 = n366 & n367;
  assign n370 = ~n368 & ~n369;
  assign n371 = n285 & n370;
  assign n372 = ~n285 & ~n370;
  assign n373 = ~n371 & ~n372;
  assign n374 = a4_0 & a4_1;
  assign n375 = ~a4_0 & ~a4_1;
  assign n376 = ~n374 & ~n375;
  assign n377 = a4_2 & n376;
  assign n378 = ~a4_2 & ~n376;
  assign n379 = ~n377 & ~n378;
  assign n380 = a4_3 & a4_4;
  assign n381 = ~a4_3 & ~a4_4;
  assign n382 = ~n380 & ~n381;
  assign n383 = a4_5 & n382;
  assign n384 = ~a4_5 & ~n382;
  assign n385 = ~n383 & ~n384;
  assign n386 = n379 & n385;
  assign n387 = ~n379 & ~n385;
  assign n388 = ~n386 & ~n387;
  assign n389 = n373 & n388;
  assign n390 = ~n373 & ~n388;
  assign n391 = ~n389 & ~n390;
  assign n392 = n365 & n391;
  assign n393 = ~n365 & ~n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n296 & ~n299;
  assign n396 = ~n302 & ~n305;
  assign n397 = ~n395 & ~n396;
  assign n398 = n395 & n396;
  assign n399 = ~n397 & ~n398;
  assign n400 = n308 & n399;
  assign n401 = ~n308 & ~n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n319 & ~n322;
  assign n404 = ~n290 & ~n293;
  assign n405 = ~n403 & ~n404;
  assign n406 = n403 & n404;
  assign n407 = ~n405 & ~n406;
  assign n408 = n402 & n407;
  assign n409 = ~n402 & ~n407;
  assign n410 = ~n408 & ~n409;
  assign n411 = n394 & n410;
  assign n412 = ~n394 & ~n410;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n338 & ~n341;
  assign n415 = ~n327 & ~n330;
  assign n416 = ~n311 & ~n314;
  assign n417 = ~n415 & ~n416;
  assign n418 = n415 & n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = n333 & n419;
  assign n421 = ~n333 & ~n419;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~n414 & n422;
  assign n424 = n414 & ~n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = n413 & n425;
  assign n427 = ~n413 & ~n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n350 & n428;
  assign n430 = n350 & ~n428;
  assign s4 = ~n429 & ~n430;
  assign n432 = ~n423 & ~n426;
  assign n433 = a5_6 & a5_7;
  assign n434 = ~a5_6 & ~a5_7;
  assign n435 = ~n433 & ~n434;
  assign n436 = a5_8 & n435;
  assign n437 = ~a5_8 & ~n435;
  assign n438 = ~n436 & ~n437;
  assign n439 = a5_9 & a5_10;
  assign n440 = ~a5_9 & ~a5_10;
  assign n441 = ~n439 & ~n440;
  assign n442 = a5_11 & n441;
  assign n443 = ~a5_11 & ~n441;
  assign n444 = ~n442 & ~n443;
  assign n445 = n438 & n444;
  assign n446 = ~n438 & ~n444;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n351 & ~n354;
  assign n449 = ~n357 & ~n360;
  assign n450 = ~n448 & ~n449;
  assign n451 = n448 & n449;
  assign n452 = ~n450 & ~n451;
  assign n453 = n363 & n452;
  assign n454 = ~n363 & ~n452;
  assign n455 = ~n453 & ~n454;
  assign n456 = a5_0 & a5_1;
  assign n457 = ~a5_0 & ~a5_1;
  assign n458 = ~n456 & ~n457;
  assign n459 = a5_2 & n458;
  assign n460 = ~a5_2 & ~n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = a5_3 & a5_4;
  assign n463 = ~a5_3 & ~a5_4;
  assign n464 = ~n462 & ~n463;
  assign n465 = a5_5 & n464;
  assign n466 = ~a5_5 & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = n461 & n467;
  assign n469 = ~n461 & ~n467;
  assign n470 = ~n468 & ~n469;
  assign n471 = n455 & n470;
  assign n472 = ~n455 & ~n470;
  assign n473 = ~n471 & ~n472;
  assign n474 = n447 & n473;
  assign n475 = ~n447 & ~n473;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n374 & ~n377;
  assign n478 = ~n380 & ~n383;
  assign n479 = ~n477 & ~n478;
  assign n480 = n477 & n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = n386 & n481;
  assign n483 = ~n386 & ~n481;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n397 & ~n400;
  assign n486 = ~n368 & ~n371;
  assign n487 = ~n485 & ~n486;
  assign n488 = n485 & n486;
  assign n489 = ~n487 & ~n488;
  assign n490 = n484 & n489;
  assign n491 = ~n484 & ~n489;
  assign n492 = ~n490 & ~n491;
  assign n493 = n476 & n492;
  assign n494 = ~n476 & ~n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n417 & ~n420;
  assign n497 = ~n405 & ~n408;
  assign n498 = ~n389 & ~n392;
  assign n499 = ~n497 & ~n498;
  assign n500 = n497 & n498;
  assign n501 = ~n499 & ~n500;
  assign n502 = n411 & n501;
  assign n503 = ~n411 & ~n501;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n496 & n504;
  assign n506 = n496 & ~n504;
  assign n507 = ~n505 & ~n506;
  assign n508 = n495 & n507;
  assign n509 = ~n495 & ~n507;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n432 & n510;
  assign n512 = n432 & ~n510;
  assign n513 = ~n511 & ~n512;
  assign n514 = n429 & n513;
  assign n515 = ~n429 & ~n513;
  assign s5 = ~n514 & ~n515;
  assign n517 = ~n511 & ~n514;
  assign n518 = ~n505 & ~n508;
  assign n519 = a6_6 & a6_7;
  assign n520 = ~a6_6 & ~a6_7;
  assign n521 = ~n519 & ~n520;
  assign n522 = a6_8 & n521;
  assign n523 = ~a6_8 & ~n521;
  assign n524 = ~n522 & ~n523;
  assign n525 = a6_9 & a6_10;
  assign n526 = ~a6_9 & ~a6_10;
  assign n527 = ~n525 & ~n526;
  assign n528 = a6_11 & n527;
  assign n529 = ~a6_11 & ~n527;
  assign n530 = ~n528 & ~n529;
  assign n531 = n524 & n530;
  assign n532 = ~n524 & ~n530;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n433 & ~n436;
  assign n535 = ~n439 & ~n442;
  assign n536 = ~n534 & ~n535;
  assign n537 = n534 & n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = n445 & n538;
  assign n540 = ~n445 & ~n538;
  assign n541 = ~n539 & ~n540;
  assign n542 = a6_0 & a6_1;
  assign n543 = ~a6_0 & ~a6_1;
  assign n544 = ~n542 & ~n543;
  assign n545 = a6_2 & n544;
  assign n546 = ~a6_2 & ~n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = a6_3 & a6_4;
  assign n549 = ~a6_3 & ~a6_4;
  assign n550 = ~n548 & ~n549;
  assign n551 = a6_5 & n550;
  assign n552 = ~a6_5 & ~n550;
  assign n553 = ~n551 & ~n552;
  assign n554 = n547 & n553;
  assign n555 = ~n547 & ~n553;
  assign n556 = ~n554 & ~n555;
  assign n557 = n541 & n556;
  assign n558 = ~n541 & ~n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = n533 & n559;
  assign n561 = ~n533 & ~n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n456 & ~n459;
  assign n564 = ~n462 & ~n465;
  assign n565 = ~n563 & ~n564;
  assign n566 = n563 & n564;
  assign n567 = ~n565 & ~n566;
  assign n568 = n468 & n567;
  assign n569 = ~n468 & ~n567;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n479 & ~n482;
  assign n572 = ~n450 & ~n453;
  assign n573 = ~n571 & ~n572;
  assign n574 = n571 & n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = n570 & n575;
  assign n577 = ~n570 & ~n575;
  assign n578 = ~n576 & ~n577;
  assign n579 = n562 & n578;
  assign n580 = ~n562 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n499 & ~n502;
  assign n583 = ~n487 & ~n490;
  assign n584 = ~n471 & ~n474;
  assign n585 = ~n583 & ~n584;
  assign n586 = n583 & n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = n493 & n587;
  assign n589 = ~n493 & ~n587;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n582 & n590;
  assign n592 = n582 & ~n590;
  assign n593 = ~n591 & ~n592;
  assign n594 = n581 & n593;
  assign n595 = ~n581 & ~n593;
  assign n596 = ~n594 & ~n595;
  assign n597 = ~n518 & n596;
  assign n598 = n518 & ~n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n517 & n599;
  assign n601 = n517 & ~n599;
  assign s6 = ~n600 & ~n601;
  assign n603 = ~n597 & ~n600;
  assign n604 = ~n591 & ~n594;
  assign n605 = a7_6 & a7_7;
  assign n606 = ~a7_6 & ~a7_7;
  assign n607 = ~n605 & ~n606;
  assign n608 = a7_8 & n607;
  assign n609 = ~a7_8 & ~n607;
  assign n610 = ~n608 & ~n609;
  assign n611 = a7_9 & a7_10;
  assign n612 = ~a7_9 & ~a7_10;
  assign n613 = ~n611 & ~n612;
  assign n614 = a7_11 & n613;
  assign n615 = ~a7_11 & ~n613;
  assign n616 = ~n614 & ~n615;
  assign n617 = n610 & n616;
  assign n618 = ~n610 & ~n616;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n519 & ~n522;
  assign n621 = ~n525 & ~n528;
  assign n622 = ~n620 & ~n621;
  assign n623 = n620 & n621;
  assign n624 = ~n622 & ~n623;
  assign n625 = n531 & n624;
  assign n626 = ~n531 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = a7_0 & a7_1;
  assign n629 = ~a7_0 & ~a7_1;
  assign n630 = ~n628 & ~n629;
  assign n631 = a7_2 & n630;
  assign n632 = ~a7_2 & ~n630;
  assign n633 = ~n631 & ~n632;
  assign n634 = a7_3 & a7_4;
  assign n635 = ~a7_3 & ~a7_4;
  assign n636 = ~n634 & ~n635;
  assign n637 = a7_5 & n636;
  assign n638 = ~a7_5 & ~n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = n633 & n639;
  assign n641 = ~n633 & ~n639;
  assign n642 = ~n640 & ~n641;
  assign n643 = n627 & n642;
  assign n644 = ~n627 & ~n642;
  assign n645 = ~n643 & ~n644;
  assign n646 = n619 & n645;
  assign n647 = ~n619 & ~n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n542 & ~n545;
  assign n650 = ~n548 & ~n551;
  assign n651 = ~n649 & ~n650;
  assign n652 = n649 & n650;
  assign n653 = ~n651 & ~n652;
  assign n654 = n554 & n653;
  assign n655 = ~n554 & ~n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n565 & ~n568;
  assign n658 = ~n536 & ~n539;
  assign n659 = ~n657 & ~n658;
  assign n660 = n657 & n658;
  assign n661 = ~n659 & ~n660;
  assign n662 = n656 & n661;
  assign n663 = ~n656 & ~n661;
  assign n664 = ~n662 & ~n663;
  assign n665 = n648 & n664;
  assign n666 = ~n648 & ~n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n585 & ~n588;
  assign n669 = ~n573 & ~n576;
  assign n670 = ~n557 & ~n560;
  assign n671 = ~n669 & ~n670;
  assign n672 = n669 & n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = n579 & n673;
  assign n675 = ~n579 & ~n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n668 & n676;
  assign n678 = n668 & ~n676;
  assign n679 = ~n677 & ~n678;
  assign n680 = n667 & n679;
  assign n681 = ~n667 & ~n679;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~n604 & n682;
  assign n684 = n604 & ~n682;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n603 & n685;
  assign n687 = n603 & ~n685;
  assign s7 = ~n686 & ~n687;
  assign n689 = ~n683 & ~n686;
  assign n690 = ~n677 & ~n680;
  assign n691 = ~n605 & ~n608;
  assign n692 = ~n611 & ~n614;
  assign n693 = ~n691 & ~n692;
  assign n694 = n691 & n692;
  assign n695 = ~n693 & ~n694;
  assign n696 = n617 & n695;
  assign n697 = ~n617 & ~n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n628 & ~n631;
  assign n700 = ~n634 & ~n637;
  assign n701 = ~n699 & ~n700;
  assign n702 = n699 & n700;
  assign n703 = ~n701 & ~n702;
  assign n704 = n640 & n703;
  assign n705 = ~n640 & ~n703;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n651 & ~n654;
  assign n708 = ~n622 & ~n625;
  assign n709 = ~n707 & ~n708;
  assign n710 = n707 & n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = n706 & n711;
  assign n713 = ~n706 & ~n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = n698 & n714;
  assign n716 = ~n698 & ~n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~n671 & ~n674;
  assign n719 = ~n659 & ~n662;
  assign n720 = ~n643 & ~n646;
  assign n721 = ~n719 & ~n720;
  assign n722 = n719 & n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = n665 & n723;
  assign n725 = ~n665 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n718 & n726;
  assign n728 = n718 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = n717 & n729;
  assign n731 = ~n717 & ~n729;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n690 & n732;
  assign n734 = n690 & ~n732;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~n689 & n735;
  assign n737 = n689 & ~n735;
  assign s8 = ~n736 & ~n737;
  assign n739 = ~n733 & ~n736;
  assign n740 = ~n727 & ~n730;
  assign n741 = ~n701 & ~n704;
  assign n742 = ~n693 & ~n696;
  assign n743 = ~n741 & ~n742;
  assign n744 = n741 & n742;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n721 & ~n724;
  assign n747 = ~n709 & ~n712;
  assign n748 = n715 & ~n747;
  assign n749 = ~n715 & n747;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~n746 & n750;
  assign n752 = n746 & ~n750;
  assign n753 = ~n751 & ~n752;
  assign n754 = n745 & n753;
  assign n755 = ~n745 & ~n753;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n740 & n756;
  assign n758 = n740 & ~n756;
  assign n759 = ~n757 & ~n758;
  assign n760 = ~n739 & n759;
  assign n761 = n739 & ~n759;
  assign s9 = ~n760 & ~n761;
  assign n763 = ~n757 & ~n760;
  assign n764 = ~n751 & ~n754;
  assign n765 = n743 & n748;
  assign n766 = ~n743 & ~n748;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n764 & n767;
  assign n769 = n764 & ~n767;
  assign n770 = ~n768 & ~n769;
  assign n771 = ~n763 & n770;
  assign n772 = n763 & ~n770;
  assign s10 = ~n771 & ~n772;
  assign s12 = n765 & n771;
  assign n775 = ~n765 & ~n768;
  assign n776 = ~n771 & n775;
  assign s11 = ~s12 & ~n776;
endmodule


