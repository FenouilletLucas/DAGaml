// Benchmark "frg2" written by ABC on Tue May 16 16:07:49 2017

module frg2 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4, c0, c1, c2, c3, c4, d0,
    d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2, f3, f4, g0, g1, g2, g3,
    g4, h0, h1, h2, h3, h4, i0, i1, i2, i3, i4, j0, j1, j2, j3, j4, k0, k1,
    k2, k3, k4, l0, l1, l2, l3, l4, m0, m1, m2, m3, m4, n0, n1, n2, n3, n4,
    o0, o1, o2, o3, p0, p1, p2, p3, q0, q1, q2, q3, r1, r2, r3, s0, s1, s2,
    s3, t0, t1, t2, t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2, w3, x0,
    x1, x2, x3, y0, y1, y2, y3, z0, z1, z2, z3,
    a5, a6, a7, a8, a9, b5, b6, b7, b8, b9, c5, c6, c7, c8, c9, d5, d6, d7,
    d8, d9, e5, e6, e7, e8, e9, f5, f6, f7, f8, f9, g5, g6, g7, g8, g9, h5,
    h6, h7, h8, h9, i5, i6, i7, i8, i9, j5, j6, j7, j8, j9, k5, k6, k7, k8,
    k9, l5, l6, l7, l8, l9, m5, m6, m7, m8, m9, n5, n6, n7, n8, n9, o4, o5,
    o6, o7, o8, o9, p4, p5, p6, p7, p8, p9, q4, q5, q6, q7, q8, q9, r4, r5,
    r6, r7, r8, r9, s4, s5, s6, s7, s8, s9, t4, t5, t6, t7, t8, t9, u4, u5,
    u6, u7, u8, u9, v4, v5, v6, v7, v8, v9, w4, w5, w6, w7, w8, w9, x4, x5,
    x6, x7, x8, y4, y5, y6, y7, y8, z4, z5, z6, z7, z8  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4, c0, c1, c2, c3,
    c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2, f3, f4, g0, g1,
    g2, g3, g4, h0, h1, h2, h3, h4, i0, i1, i2, i3, i4, j0, j1, j2, j3, j4,
    k0, k1, k2, k3, k4, l0, l1, l2, l3, l4, m0, m1, m2, m3, m4, n0, n1, n2,
    n3, n4, o0, o1, o2, o3, p0, p1, p2, p3, q0, q1, q2, q3, r1, r2, r3, s0,
    s1, s2, s3, t0, t1, t2, t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2,
    w3, x0, x1, x2, x3, y0, y1, y2, y3, z0, z1, z2, z3;
  output a5, a6, a7, a8, a9, b5, b6, b7, b8, b9, c5, c6, c7, c8, c9, d5, d6,
    d7, d8, d9, e5, e6, e7, e8, e9, f5, f6, f7, f8, f9, g5, g6, g7, g8, g9,
    h5, h6, h7, h8, h9, i5, i6, i7, i8, i9, j5, j6, j7, j8, j9, k5, k6, k7,
    k8, k9, l5, l6, l7, l8, l9, m5, m6, m7, m8, m9, n5, n6, n7, n8, n9, o4,
    o5, o6, o7, o8, o9, p4, p5, p6, p7, p8, p9, q4, q5, q6, q7, q8, q9, r4,
    r5, r6, r7, r8, r9, s4, s5, s6, s7, s8, s9, t4, t5, t6, t7, t8, t9, u4,
    u5, u6, u7, u8, u9, v4, v5, v6, v7, v8, v9, w4, w5, w6, w7, w8, w9, x4,
    x5, x6, x7, x8, y4, y5, y6, y7, y8, z4, z5, z6, z7, z8;
  wire n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n294,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n436, n437, n438, n439, n440, n441, n442,
    n443, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n502, n503, n504, n505, n506,
    n507, n508, n510, n511, n512, n513, n514, n515, n516, n517, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n567, n568, n569, n570, n571,
    n572, n573, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n624,
    n625, n626, n627, n628, n629, n630, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n681, n682, n683, n684, n685, n686, n687, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n853, n854, n855,
    n856, n857, n858, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1225, n1227, n1228, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1278, n1280, n1281, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1354, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1466, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1559, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1810, n1811, n1812, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1854,
    n1855, n1856, n1857, n1858, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148;
  assign n283 = ~k0 & ~l0;
  assign n284 = ~j3 & n283;
  assign n285 = k0 & l0;
  assign n286 = ~j3 & n285;
  assign n287 = m0 & ~n286;
  assign n288 = ~n284 & n287;
  assign n289 = n283 & n288;
  assign n290 = n285 & n288;
  assign n291 = r3 & n288;
  assign n292 = ~n290 & ~n291;
  assign a5 = n289 | ~n292;
  assign n294 = ~k4 & m1;
  assign a6 = ~k1 | ~n294;
  assign n296 = ~a4 & z3;
  assign n297 = ~x3 & y3;
  assign n298 = n296 & n297;
  assign n299 = ~b4 & ~c4;
  assign n300 = n298 & n299;
  assign n301 = l4 & ~n300;
  assign n302 = ~i1 & ~j1;
  assign n303 = ~h1 & n302;
  assign n304 = ~k1 & ~l1;
  assign n305 = n303 & n304;
  assign n306 = o0 & ~n305;
  assign n307 = ~q0 & n306;
  assign n308 = n0 & o0;
  assign n309 = ~q0 & n308;
  assign n310 = f0 & o0;
  assign n311 = ~q0 & n310;
  assign n312 = ~n309 & ~n311;
  assign n313 = ~n307 & n312;
  assign n314 = ~r1 & ~n305;
  assign n315 = ~n301 & n314;
  assign n316 = ~n313 & ~n315;
  assign n317 = ~n0 & n305;
  assign n318 = l4 & ~s1;
  assign n319 = n301 & n317;
  assign n320 = n316 & n319;
  assign n321 = n301 & ~n318;
  assign n322 = n316 & n321;
  assign n323 = n300 & n301;
  assign n324 = n316 & n323;
  assign n325 = ~n0 & n317;
  assign n326 = n316 & n325;
  assign n327 = ~n0 & ~n318;
  assign n328 = n316 & n327;
  assign n329 = ~n0 & n300;
  assign n330 = n316 & n329;
  assign n331 = r1 & n317;
  assign n332 = n316 & n331;
  assign n333 = r1 & ~n318;
  assign n334 = n316 & n333;
  assign n335 = r1 & n300;
  assign n336 = n316 & n335;
  assign n337 = ~n334 & ~n336;
  assign n338 = ~n332 & n337;
  assign n339 = ~n330 & n338;
  assign n340 = ~n328 & n339;
  assign n341 = ~n326 & n340;
  assign n342 = ~n324 & n341;
  assign n343 = ~n322 & n342;
  assign a7 = n320 | ~n343;
  assign n345 = ~m0 & n317;
  assign n346 = l4 & ~s2;
  assign n347 = k0 & ~l0;
  assign n348 = p & n347;
  assign n349 = h & l0;
  assign n350 = h & ~k0;
  assign n351 = ~n349 & ~n350;
  assign n352 = ~n348 & n351;
  assign n353 = ~m0 & ~n0;
  assign n354 = n305 & n353;
  assign n355 = ~r2 & ~n301;
  assign n356 = ~n354 & n355;
  assign n357 = ~n300 & n346;
  assign n358 = ~n345 & n357;
  assign n359 = n345 & n352;
  assign n360 = ~n356 & ~n359;
  assign n361 = ~n358 & n360;
  assign n362 = o0 & ~q0;
  assign a8 = n361 & n362;
  assign n364 = ~j1 & ~k1;
  assign n365 = ~l1 & n364;
  assign n366 = ~k1 & z0;
  assign n367 = ~l1 & n366;
  assign n368 = a1 & ~j1;
  assign n369 = ~l1 & n368;
  assign n370 = a1 & z0;
  assign n371 = ~l1 & n370;
  assign n372 = b1 & n364;
  assign n373 = b1 & n366;
  assign n374 = b1 & n368;
  assign n375 = b1 & n370;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n373 & n376;
  assign n378 = ~n372 & n377;
  assign n379 = ~n371 & n378;
  assign n380 = ~n369 & n379;
  assign n381 = ~n367 & n380;
  assign n382 = ~n365 & n381;
  assign n383 = i1 & ~y0;
  assign n384 = h1 & ~x0;
  assign n385 = ~n382 & ~n384;
  assign n386 = ~n383 & n385;
  assign n387 = j1 & k1;
  assign n388 = ~n305 & ~n386;
  assign n389 = ~n387 & n388;
  assign n390 = f4 & ~g4;
  assign n391 = e4 & n390;
  assign n392 = ~h4 & n391;
  assign n393 = ~j1 & ~n392;
  assign n394 = n389 & n393;
  assign n395 = ~l1 & ~n392;
  assign n396 = n389 & n395;
  assign n397 = ~n394 & ~n396;
  assign n398 = k1 & l1;
  assign n399 = k4 & ~n397;
  assign n400 = ~n398 & n399;
  assign n401 = ~j1 & n304;
  assign n402 = n302 & n304;
  assign n403 = n401 & n402;
  assign n404 = n400 & n403;
  assign n405 = ~h1 & n401;
  assign n406 = n400 & n405;
  assign n407 = ~h1 & ~i1;
  assign n408 = n400 & n407;
  assign n409 = ~i1 & n402;
  assign n410 = n400 & n409;
  assign n411 = ~n408 & ~n410;
  assign n412 = ~n406 & n411;
  assign n413 = ~n404 & n412;
  assign n414 = ~q0 & r3;
  assign n415 = j1 & l1;
  assign n416 = ~n387 & ~n415;
  assign n417 = ~n398 & n416;
  assign n418 = ~n401 & n417;
  assign n419 = h1 & n417;
  assign n420 = i1 & n417;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n418 & n421;
  assign n423 = i1 & ~n401;
  assign n424 = h1 & ~n402;
  assign n425 = ~n422 & ~n424;
  assign n426 = ~n423 & n425;
  assign n427 = k4 & s3;
  assign n428 = ~n392 & n427;
  assign n429 = ~q0 & ~n386;
  assign n430 = o0 & n429;
  assign n431 = n428 & n430;
  assign n432 = n426 & n431;
  assign n433 = o0 & n414;
  assign n434 = n413 & n433;
  assign a9 = n432 | n434;
  assign n436 = ~k3 & n283;
  assign n437 = ~k3 & n285;
  assign n438 = m0 & ~n437;
  assign n439 = ~n436 & n438;
  assign n440 = n283 & n439;
  assign n441 = n285 & n439;
  assign n442 = s3 & n439;
  assign n443 = ~n441 & ~n442;
  assign b5 = n440 | ~n443;
  assign b6 = ~l1 | ~n294;
  assign n446 = e0 & o0;
  assign n447 = ~q0 & n446;
  assign n448 = ~n309 & ~n447;
  assign n449 = ~n307 & n448;
  assign n450 = ~s1 & ~n305;
  assign n451 = ~n301 & n450;
  assign n452 = ~n449 & ~n451;
  assign n453 = l4 & ~t1;
  assign n454 = n319 & n452;
  assign n455 = n301 & ~n453;
  assign n456 = n452 & n455;
  assign n457 = n323 & n452;
  assign n458 = n325 & n452;
  assign n459 = ~n0 & ~n453;
  assign n460 = n452 & n459;
  assign n461 = n329 & n452;
  assign n462 = s1 & n317;
  assign n463 = n452 & n462;
  assign n464 = s1 & ~n453;
  assign n465 = n452 & n464;
  assign n466 = s1 & n300;
  assign n467 = n452 & n466;
  assign n468 = ~n465 & ~n467;
  assign n469 = ~n463 & n468;
  assign n470 = ~n461 & n469;
  assign n471 = ~n460 & n470;
  assign n472 = ~n458 & n471;
  assign n473 = ~n457 & n472;
  assign n474 = ~n456 & n473;
  assign b7 = n454 | ~n474;
  assign n476 = ~k0 & l0;
  assign n477 = n305 & ~n476;
  assign n478 = ~n347 & n477;
  assign n479 = n353 & n478;
  assign n480 = ~n347 & ~n476;
  assign n481 = ~l4 & s2;
  assign n482 = ~n479 & n481;
  assign n483 = i & n345;
  assign n484 = n480 & n483;
  assign n485 = ~n482 & ~n484;
  assign n486 = l4 & t2;
  assign n487 = n283 & n305;
  assign n488 = n285 & n305;
  assign n489 = ~n487 & ~n488;
  assign n490 = n353 & ~n489;
  assign n491 = ~n300 & ~n486;
  assign n492 = n485 & n491;
  assign n493 = ~s2 & ~n486;
  assign n494 = n485 & n493;
  assign n495 = ~s2 & n300;
  assign n496 = n485 & n495;
  assign n497 = n485 & n490;
  assign n498 = ~n496 & ~n497;
  assign n499 = ~n494 & n498;
  assign n500 = ~n492 & n499;
  assign b8 = n362 & n500;
  assign n502 = ~q0 & s3;
  assign n503 = k4 & t3;
  assign n504 = ~n392 & n503;
  assign n505 = n430 & n504;
  assign n506 = n426 & n505;
  assign n507 = o0 & n502;
  assign n508 = n413 & n507;
  assign b9 = n506 | n508;
  assign n510 = ~l3 & n283;
  assign n511 = ~l3 & n285;
  assign n512 = m0 & ~n511;
  assign n513 = ~n510 & n512;
  assign n514 = n283 & n513;
  assign n515 = n285 & n513;
  assign n516 = t3 & n513;
  assign n517 = ~n515 & ~n516;
  assign c5 = n514 | ~n517;
  assign c6 = ~h1 | ~l4;
  assign n520 = d0 & o0;
  assign n521 = ~q0 & n520;
  assign n522 = ~n309 & ~n521;
  assign n523 = ~n307 & n522;
  assign n524 = ~t1 & ~n305;
  assign n525 = ~n301 & n524;
  assign n526 = ~n523 & ~n525;
  assign n527 = l4 & ~u1;
  assign n528 = n319 & n526;
  assign n529 = n301 & ~n527;
  assign n530 = n526 & n529;
  assign n531 = n323 & n526;
  assign n532 = n325 & n526;
  assign n533 = ~n0 & ~n527;
  assign n534 = n526 & n533;
  assign n535 = n329 & n526;
  assign n536 = t1 & n317;
  assign n537 = n526 & n536;
  assign n538 = t1 & ~n527;
  assign n539 = n526 & n538;
  assign n540 = t1 & n300;
  assign n541 = n526 & n540;
  assign n542 = ~n539 & ~n541;
  assign n543 = ~n537 & n542;
  assign n544 = ~n535 & n543;
  assign n545 = ~n534 & n544;
  assign n546 = ~n532 & n545;
  assign n547 = ~n531 & n546;
  assign n548 = ~n530 & n547;
  assign c7 = n528 | ~n548;
  assign n550 = ~l4 & t2;
  assign n551 = ~n479 & n550;
  assign n552 = j & n345;
  assign n553 = n480 & n552;
  assign n554 = ~n551 & ~n553;
  assign n555 = l4 & u2;
  assign n556 = ~n300 & ~n555;
  assign n557 = n554 & n556;
  assign n558 = ~t2 & ~n555;
  assign n559 = n554 & n558;
  assign n560 = ~t2 & n300;
  assign n561 = n554 & n560;
  assign n562 = n490 & n554;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~n559 & n563;
  assign n565 = ~n557 & n564;
  assign c8 = n362 & n565;
  assign n567 = ~q0 & t3;
  assign n568 = k4 & u3;
  assign n569 = ~n392 & n568;
  assign n570 = n430 & n569;
  assign n571 = n426 & n570;
  assign n572 = o0 & n567;
  assign n573 = n413 & n572;
  assign c9 = n571 | n573;
  assign d5 = m0 & m3;
  assign d6 = ~i1 | ~l4;
  assign n577 = m0 & o0;
  assign n578 = ~q0 & n577;
  assign n579 = ~n309 & ~n578;
  assign n580 = ~n307 & n579;
  assign n581 = ~u1 & ~n305;
  assign n582 = ~n301 & n581;
  assign n583 = ~n580 & ~n582;
  assign n584 = l4 & ~v1;
  assign n585 = n319 & n583;
  assign n586 = n301 & ~n584;
  assign n587 = n583 & n586;
  assign n588 = n323 & n583;
  assign n589 = n325 & n583;
  assign n590 = ~n0 & ~n584;
  assign n591 = n583 & n590;
  assign n592 = n329 & n583;
  assign n593 = u1 & n317;
  assign n594 = n583 & n593;
  assign n595 = u1 & ~n584;
  assign n596 = n583 & n595;
  assign n597 = u1 & n300;
  assign n598 = n583 & n597;
  assign n599 = ~n596 & ~n598;
  assign n600 = ~n594 & n599;
  assign n601 = ~n592 & n600;
  assign n602 = ~n591 & n601;
  assign n603 = ~n589 & n602;
  assign n604 = ~n588 & n603;
  assign n605 = ~n587 & n604;
  assign d7 = n585 | ~n605;
  assign n607 = ~l4 & u2;
  assign n608 = ~n479 & n607;
  assign n609 = k & n345;
  assign n610 = n480 & n609;
  assign n611 = ~n608 & ~n610;
  assign n612 = l4 & v2;
  assign n613 = ~n300 & ~n612;
  assign n614 = n611 & n613;
  assign n615 = ~u2 & ~n612;
  assign n616 = n611 & n615;
  assign n617 = ~u2 & n300;
  assign n618 = n611 & n617;
  assign n619 = n490 & n611;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~n616 & n620;
  assign n622 = ~n614 & n621;
  assign d8 = n362 & n622;
  assign n624 = ~q0 & u3;
  assign n625 = k4 & v3;
  assign n626 = ~n392 & n625;
  assign n627 = n430 & n626;
  assign n628 = n426 & n627;
  assign n629 = o0 & n624;
  assign n630 = n413 & n629;
  assign d9 = n628 | n630;
  assign e5 = m0 & n3;
  assign e6 = ~j1 | ~l4;
  assign n634 = k0 & o0;
  assign n635 = ~q0 & n634;
  assign n636 = ~n309 & ~n635;
  assign n637 = ~n307 & n636;
  assign n638 = ~v1 & ~n305;
  assign n639 = ~n301 & n638;
  assign n640 = ~n637 & ~n639;
  assign n641 = l4 & ~w1;
  assign n642 = n319 & n640;
  assign n643 = n301 & ~n641;
  assign n644 = n640 & n643;
  assign n645 = n323 & n640;
  assign n646 = n325 & n640;
  assign n647 = ~n0 & ~n641;
  assign n648 = n640 & n647;
  assign n649 = n329 & n640;
  assign n650 = v1 & n317;
  assign n651 = n640 & n650;
  assign n652 = v1 & ~n641;
  assign n653 = n640 & n652;
  assign n654 = v1 & n300;
  assign n655 = n640 & n654;
  assign n656 = ~n653 & ~n655;
  assign n657 = ~n651 & n656;
  assign n658 = ~n649 & n657;
  assign n659 = ~n648 & n658;
  assign n660 = ~n646 & n659;
  assign n661 = ~n645 & n660;
  assign n662 = ~n644 & n661;
  assign e7 = n642 | ~n662;
  assign n664 = ~l4 & v2;
  assign n665 = ~n479 & n664;
  assign n666 = l & n345;
  assign n667 = n480 & n666;
  assign n668 = ~n665 & ~n667;
  assign n669 = l4 & w2;
  assign n670 = ~n300 & ~n669;
  assign n671 = n668 & n670;
  assign n672 = ~v2 & ~n669;
  assign n673 = n668 & n672;
  assign n674 = ~v2 & n300;
  assign n675 = n668 & n674;
  assign n676 = n490 & n668;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n673 & n677;
  assign n679 = ~n671 & n678;
  assign e8 = n362 & n679;
  assign n681 = ~q0 & v3;
  assign n682 = k4 & w3;
  assign n683 = ~n392 & n682;
  assign n684 = n430 & n683;
  assign n685 = n426 & n684;
  assign n686 = o0 & n681;
  assign n687 = n413 & n686;
  assign e9 = n685 | n687;
  assign f5 = m0 & o3;
  assign f6 = ~k1 | ~l4;
  assign n691 = l0 & o0;
  assign n692 = ~q0 & n691;
  assign n693 = ~n309 & ~n692;
  assign n694 = ~n307 & n693;
  assign n695 = ~w1 & ~n305;
  assign n696 = ~n301 & n695;
  assign n697 = ~n694 & ~n696;
  assign n698 = l4 & ~x1;
  assign n699 = n319 & n697;
  assign n700 = n301 & ~n698;
  assign n701 = n697 & n700;
  assign n702 = n323 & n697;
  assign n703 = n325 & n697;
  assign n704 = ~n0 & ~n698;
  assign n705 = n697 & n704;
  assign n706 = n329 & n697;
  assign n707 = w1 & n317;
  assign n708 = n697 & n707;
  assign n709 = w1 & ~n698;
  assign n710 = n697 & n709;
  assign n711 = w1 & n300;
  assign n712 = n697 & n711;
  assign n713 = ~n710 & ~n712;
  assign n714 = ~n708 & n713;
  assign n715 = ~n706 & n714;
  assign n716 = ~n705 & n715;
  assign n717 = ~n703 & n716;
  assign n718 = ~n702 & n717;
  assign n719 = ~n701 & n718;
  assign f7 = n699 | ~n719;
  assign n721 = ~l4 & w2;
  assign n722 = ~n479 & n721;
  assign n723 = m & n345;
  assign n724 = n480 & n723;
  assign n725 = ~n722 & ~n724;
  assign n726 = l4 & x2;
  assign n727 = ~n300 & ~n726;
  assign n728 = n725 & n727;
  assign n729 = ~w2 & ~n726;
  assign n730 = n725 & n729;
  assign n731 = ~w2 & n300;
  assign n732 = n725 & n731;
  assign n733 = n490 & n725;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n730 & n734;
  assign n736 = ~n728 & n735;
  assign f8 = n362 & n736;
  assign n738 = j1 & ~n304;
  assign n739 = n401 & n407;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~k1 & ~n386;
  assign n742 = n740 & n741;
  assign n743 = ~l1 & ~n386;
  assign n744 = n740 & n743;
  assign n745 = ~n742 & ~n744;
  assign n746 = k4 & ~n392;
  assign n747 = ~n745 & n746;
  assign n748 = n403 & n747;
  assign n749 = n405 & n747;
  assign n750 = n407 & n747;
  assign n751 = n409 & n747;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n749 & n752;
  assign n754 = ~n748 & n753;
  assign n755 = ~q0 & w3;
  assign n756 = ~j1 & k1;
  assign n757 = v0 & n756;
  assign n758 = ~l1 & n757;
  assign n759 = ~k1 & l1;
  assign n760 = ~n304 & ~n759;
  assign n761 = ~n758 & n760;
  assign n762 = ~j1 & ~n759;
  assign n763 = ~n758 & n762;
  assign n764 = ~u0 & ~n759;
  assign n765 = ~n758 & n764;
  assign n766 = n738 & ~n758;
  assign n767 = ~w0 & ~n304;
  assign n768 = ~n758 & n767;
  assign n769 = ~j1 & ~w0;
  assign n770 = ~n758 & n769;
  assign n771 = ~u0 & ~w0;
  assign n772 = ~n758 & n771;
  assign n773 = j1 & ~u0;
  assign n774 = ~n758 & n773;
  assign n775 = ~n772 & ~n774;
  assign n776 = ~n770 & n775;
  assign n777 = ~n768 & n776;
  assign n778 = ~n766 & n777;
  assign n779 = ~n765 & n778;
  assign n780 = ~n763 & n779;
  assign n781 = ~n761 & n780;
  assign n782 = i1 & n401;
  assign n783 = t0 & n782;
  assign n784 = ~i1 & n781;
  assign n785 = ~n783 & ~n784;
  assign n786 = h1 & ~i1;
  assign n787 = ~n401 & n785;
  assign n788 = n785 & ~n786;
  assign n789 = ~s0 & n785;
  assign n790 = h1 & ~n401;
  assign n791 = h1 & ~n786;
  assign n792 = h1 & ~s0;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n790 & n793;
  assign n795 = ~n789 & n794;
  assign n796 = ~n788 & n795;
  assign n797 = ~n787 & n796;
  assign n798 = ~n386 & n746;
  assign n799 = n362 & n798;
  assign n800 = n797 & n799;
  assign n801 = o0 & n755;
  assign n802 = n754 & n801;
  assign f9 = n800 | n802;
  assign g5 = m0 & p3;
  assign g6 = ~l1 | ~l4;
  assign n806 = q & o0;
  assign n807 = ~q0 & n806;
  assign n808 = ~n309 & ~n807;
  assign n809 = ~n307 & n808;
  assign n810 = ~x1 & ~n305;
  assign n811 = ~n301 & n810;
  assign n812 = ~n809 & ~n811;
  assign n813 = l4 & ~y1;
  assign n814 = n319 & n812;
  assign n815 = n301 & ~n813;
  assign n816 = n812 & n815;
  assign n817 = n323 & n812;
  assign n818 = n325 & n812;
  assign n819 = ~n0 & ~n813;
  assign n820 = n812 & n819;
  assign n821 = n329 & n812;
  assign n822 = x1 & n317;
  assign n823 = n812 & n822;
  assign n824 = x1 & ~n813;
  assign n825 = n812 & n824;
  assign n826 = x1 & n300;
  assign n827 = n812 & n826;
  assign n828 = ~n825 & ~n827;
  assign n829 = ~n823 & n828;
  assign n830 = ~n821 & n829;
  assign n831 = ~n820 & n830;
  assign n832 = ~n818 & n831;
  assign n833 = ~n817 & n832;
  assign n834 = ~n816 & n833;
  assign g7 = n814 | ~n834;
  assign n836 = ~l4 & x2;
  assign n837 = ~n479 & n836;
  assign n838 = n & n345;
  assign n839 = n480 & n838;
  assign n840 = ~n837 & ~n839;
  assign n841 = l4 & y2;
  assign n842 = ~n300 & ~n841;
  assign n843 = n840 & n842;
  assign n844 = ~x2 & ~n841;
  assign n845 = n840 & n844;
  assign n846 = ~x2 & n300;
  assign n847 = n840 & n846;
  assign n848 = n490 & n840;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~n845 & n849;
  assign n851 = ~n843 & n850;
  assign g8 = n362 & n851;
  assign n853 = ~n307 & ~n309;
  assign n854 = l4 & x3;
  assign n855 = ~n300 & n854;
  assign n856 = ~n853 & ~n855;
  assign n857 = n301 & n856;
  assign n858 = x3 & n856;
  assign g9 = n857 | n858;
  assign h5 = m0 & q3;
  assign n861 = r & o0;
  assign n862 = ~q0 & n861;
  assign n863 = ~n309 & ~n862;
  assign n864 = ~n307 & n863;
  assign n865 = ~y1 & ~n305;
  assign n866 = ~n301 & n865;
  assign n867 = ~n864 & ~n866;
  assign n868 = l4 & ~z1;
  assign n869 = n319 & n867;
  assign n870 = n301 & ~n868;
  assign n871 = n867 & n870;
  assign n872 = n323 & n867;
  assign n873 = n325 & n867;
  assign n874 = ~n0 & ~n868;
  assign n875 = n867 & n874;
  assign n876 = n329 & n867;
  assign n877 = y1 & n317;
  assign n878 = n867 & n877;
  assign n879 = y1 & ~n868;
  assign n880 = n867 & n879;
  assign n881 = y1 & n300;
  assign n882 = n867 & n881;
  assign n883 = ~n880 & ~n882;
  assign n884 = ~n878 & n883;
  assign n885 = ~n876 & n884;
  assign n886 = ~n875 & n885;
  assign n887 = ~n873 & n886;
  assign n888 = ~n872 & n887;
  assign n889 = ~n871 & n888;
  assign h7 = n869 | ~n889;
  assign n891 = ~l4 & y2;
  assign n892 = ~n479 & n891;
  assign n893 = o & n345;
  assign n894 = n480 & n893;
  assign n895 = ~n892 & ~n894;
  assign n896 = l4 & z2;
  assign n897 = ~n300 & ~n896;
  assign n898 = n895 & n897;
  assign n899 = ~y2 & ~n896;
  assign n900 = n895 & n899;
  assign n901 = ~y2 & n300;
  assign n902 = n895 & n901;
  assign n903 = n490 & n895;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n900 & n904;
  assign n906 = ~n898 & n905;
  assign h8 = n362 & n906;
  assign n908 = l4 & ~x3;
  assign n909 = ~n300 & n908;
  assign n910 = ~x3 & ~y3;
  assign n911 = ~n300 & n910;
  assign n912 = l4 & n911;
  assign n913 = ~q0 & ~n305;
  assign n914 = ~n912 & n913;
  assign n915 = n0 & ~q0;
  assign n916 = ~n912 & n915;
  assign n917 = ~n914 & ~n916;
  assign n918 = o0 & ~n917;
  assign n919 = y3 & ~n909;
  assign h9 = ~n918 | n919;
  assign i5 = m0 & r3;
  assign n922 = s & o0;
  assign n923 = ~q0 & n922;
  assign n924 = ~n309 & ~n923;
  assign n925 = ~n307 & n924;
  assign n926 = ~z1 & ~n305;
  assign n927 = ~n301 & n926;
  assign n928 = ~n925 & ~n927;
  assign n929 = ~a2 & l4;
  assign n930 = n319 & n928;
  assign n931 = n301 & ~n929;
  assign n932 = n928 & n931;
  assign n933 = n323 & n928;
  assign n934 = n325 & n928;
  assign n935 = ~n0 & ~n929;
  assign n936 = n928 & n935;
  assign n937 = n329 & n928;
  assign n938 = z1 & n317;
  assign n939 = n928 & n938;
  assign n940 = z1 & ~n929;
  assign n941 = n928 & n940;
  assign n942 = z1 & n300;
  assign n943 = n928 & n942;
  assign n944 = ~n941 & ~n943;
  assign n945 = ~n939 & n944;
  assign n946 = ~n937 & n945;
  assign n947 = ~n936 & n946;
  assign n948 = ~n934 & n947;
  assign n949 = ~n933 & n948;
  assign n950 = ~n932 & n949;
  assign i7 = n930 | ~n950;
  assign n952 = n345 & n480;
  assign n953 = ~n301 & ~n952;
  assign n954 = ~q0 & z2;
  assign n955 = ~q0 & n305;
  assign n956 = o0 & n955;
  assign n957 = p & n353;
  assign n958 = n956 & n957;
  assign n959 = n480 & n958;
  assign n960 = o0 & n954;
  assign n961 = n953 & n960;
  assign i8 = n959 | n961;
  assign n963 = l4 & y3;
  assign n964 = ~x3 & ~n300;
  assign n965 = n963 & n964;
  assign n966 = n297 & ~n300;
  assign n967 = l4 & ~z3;
  assign n968 = n966 & n967;
  assign n969 = n913 & ~n968;
  assign n970 = n915 & ~n968;
  assign n971 = ~n969 & ~n970;
  assign n972 = o0 & ~n971;
  assign n973 = z3 & ~n965;
  assign i9 = ~n972 | n973;
  assign j5 = m0 & s3;
  assign n976 = t & o0;
  assign n977 = ~q0 & n976;
  assign n978 = ~n309 & ~n977;
  assign n979 = ~n307 & n978;
  assign n980 = ~a2 & ~n305;
  assign n981 = ~n301 & n980;
  assign n982 = ~n979 & ~n981;
  assign n983 = ~b2 & l4;
  assign n984 = n319 & n982;
  assign n985 = n301 & ~n983;
  assign n986 = n982 & n985;
  assign n987 = n323 & n982;
  assign n988 = n325 & n982;
  assign n989 = ~n0 & ~n983;
  assign n990 = n982 & n989;
  assign n991 = n329 & n982;
  assign n992 = a2 & n317;
  assign n993 = n982 & n992;
  assign n994 = a2 & ~n983;
  assign n995 = n982 & n994;
  assign n996 = a2 & n300;
  assign n997 = n982 & n996;
  assign n998 = ~n995 & ~n997;
  assign n999 = ~n993 & n998;
  assign n1000 = ~n991 & n999;
  assign n1001 = ~n990 & n1000;
  assign n1002 = ~n988 & n1001;
  assign n1003 = ~n987 & n1002;
  assign n1004 = ~n986 & n1003;
  assign j7 = n984 | ~n1004;
  assign n1006 = a3 & ~q0;
  assign n1007 = b3 & k4;
  assign n1008 = ~n392 & n1007;
  assign n1009 = n430 & n1008;
  assign n1010 = n426 & n1009;
  assign n1011 = o0 & n1006;
  assign n1012 = n413 & n1011;
  assign j8 = n1010 | n1012;
  assign n1014 = l4 & z3;
  assign n1015 = y3 & n1014;
  assign n1016 = ~n305 & n964;
  assign n1017 = n1015 & n1016;
  assign n1018 = n0 & n305;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n305 & n480;
  assign n1021 = n1019 & n1020;
  assign n1022 = a4 & n480;
  assign n1023 = n1019 & n1022;
  assign n1024 = a4 & ~n305;
  assign n1025 = n1019 & n1024;
  assign n1026 = a4 & m0;
  assign n1027 = n1019 & n1026;
  assign n1028 = m0 & n305;
  assign n1029 = n1019 & n1028;
  assign n1030 = ~n1027 & ~n1029;
  assign n1031 = ~n1025 & n1030;
  assign n1032 = ~n1023 & n1031;
  assign n1033 = ~n1021 & n1032;
  assign n1034 = n964 & n1015;
  assign n1035 = ~a4 & l4;
  assign n1036 = z3 & n1035;
  assign n1037 = n317 & n1034;
  assign n1038 = n1033 & n1037;
  assign n1039 = n1034 & ~n1036;
  assign n1040 = n1033 & n1039;
  assign n1041 = ~n966 & n1034;
  assign n1042 = n1033 & n1041;
  assign n1043 = n325 & n1033;
  assign n1044 = ~n0 & ~n1036;
  assign n1045 = n1033 & n1044;
  assign n1046 = ~n0 & ~n966;
  assign n1047 = n1033 & n1046;
  assign n1048 = ~a4 & n317;
  assign n1049 = n1033 & n1048;
  assign n1050 = ~a4 & ~n1036;
  assign n1051 = n1033 & n1050;
  assign n1052 = ~a4 & ~n966;
  assign n1053 = n1033 & n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~n1049 & n1054;
  assign n1056 = ~n1047 & n1055;
  assign n1057 = ~n1045 & n1056;
  assign n1058 = ~n1043 & n1057;
  assign n1059 = ~n1042 & n1058;
  assign n1060 = ~n1040 & n1059;
  assign n1061 = ~n1038 & n1060;
  assign j9 = n362 & n1061;
  assign k5 = m0 & t3;
  assign n1064 = u & o0;
  assign n1065 = ~q0 & n1064;
  assign n1066 = ~n309 & ~n1065;
  assign n1067 = ~n307 & n1066;
  assign n1068 = ~b2 & ~n305;
  assign n1069 = ~n301 & n1068;
  assign n1070 = ~n1067 & ~n1069;
  assign n1071 = ~c2 & l4;
  assign n1072 = n319 & n1070;
  assign n1073 = n301 & ~n1071;
  assign n1074 = n1070 & n1073;
  assign n1075 = n323 & n1070;
  assign n1076 = n325 & n1070;
  assign n1077 = ~n0 & ~n1071;
  assign n1078 = n1070 & n1077;
  assign n1079 = n329 & n1070;
  assign n1080 = b2 & n317;
  assign n1081 = n1070 & n1080;
  assign n1082 = b2 & ~n1071;
  assign n1083 = n1070 & n1082;
  assign n1084 = b2 & n300;
  assign n1085 = n1070 & n1084;
  assign n1086 = ~n1083 & ~n1085;
  assign n1087 = ~n1081 & n1086;
  assign n1088 = ~n1079 & n1087;
  assign n1089 = ~n1078 & n1088;
  assign n1090 = ~n1076 & n1089;
  assign n1091 = ~n1075 & n1090;
  assign n1092 = ~n1074 & n1091;
  assign k7 = n1072 | ~n1092;
  assign n1094 = b3 & ~q0;
  assign n1095 = c3 & k4;
  assign n1096 = ~n392 & n1095;
  assign n1097 = n430 & n1096;
  assign n1098 = n426 & n1097;
  assign n1099 = o0 & n1094;
  assign n1100 = n413 & n1099;
  assign k8 = n1098 | n1100;
  assign n1102 = n966 & n1036;
  assign n1103 = ~n317 & ~n1102;
  assign n1104 = b4 & ~q0;
  assign n1105 = ~q0 & n964;
  assign n1106 = ~b4 & l4;
  assign n1107 = ~a4 & n1106;
  assign n1108 = y3 & z3;
  assign n1109 = o0 & n1108;
  assign n1110 = n1107 & n1109;
  assign n1111 = ~n0 & o0;
  assign n1112 = m0 & n1111;
  assign n1113 = n955 & n1112;
  assign n1114 = n1105 & n1110;
  assign n1115 = ~n317 & n1114;
  assign n1116 = ~n1113 & ~n1115;
  assign n1117 = o0 & n1104;
  assign n1118 = n1103 & n1117;
  assign k9 = ~n1116 | n1118;
  assign l5 = g1 & ~j4;
  assign n1121 = v & o0;
  assign n1122 = ~q0 & n1121;
  assign n1123 = ~n309 & ~n1122;
  assign n1124 = ~n307 & n1123;
  assign n1125 = ~c2 & ~n305;
  assign n1126 = ~n301 & n1125;
  assign n1127 = ~n1124 & ~n1126;
  assign n1128 = ~d2 & l4;
  assign n1129 = n319 & n1127;
  assign n1130 = n301 & ~n1128;
  assign n1131 = n1127 & n1130;
  assign n1132 = n323 & n1127;
  assign n1133 = n325 & n1127;
  assign n1134 = ~n0 & ~n1128;
  assign n1135 = n1127 & n1134;
  assign n1136 = n329 & n1127;
  assign n1137 = c2 & n317;
  assign n1138 = n1127 & n1137;
  assign n1139 = c2 & ~n1128;
  assign n1140 = n1127 & n1139;
  assign n1141 = c2 & n300;
  assign n1142 = n1127 & n1141;
  assign n1143 = ~n1140 & ~n1142;
  assign n1144 = ~n1138 & n1143;
  assign n1145 = ~n1136 & n1144;
  assign n1146 = ~n1135 & n1145;
  assign n1147 = ~n1133 & n1146;
  assign n1148 = ~n1132 & n1147;
  assign n1149 = ~n1131 & n1148;
  assign l7 = n1129 | ~n1149;
  assign n1151 = c3 & ~q0;
  assign n1152 = d3 & k4;
  assign n1153 = ~n392 & n1152;
  assign n1154 = n430 & n1153;
  assign n1155 = n426 & n1154;
  assign n1156 = o0 & n1151;
  assign n1157 = n413 & n1156;
  assign l8 = n1155 | n1157;
  assign n1159 = ~x3 & n1108;
  assign n1160 = ~n300 & n1159;
  assign n1161 = n1107 & n1160;
  assign n1162 = ~n317 & ~n1161;
  assign n1163 = c4 & ~q0;
  assign n1164 = ~c4 & l4;
  assign n1165 = ~b4 & n1164;
  assign n1166 = y3 & n296;
  assign n1167 = o0 & n1166;
  assign n1168 = n1165 & n1167;
  assign n1169 = ~m0 & n1111;
  assign n1170 = n955 & n1169;
  assign n1171 = n1105 & n1168;
  assign n1172 = ~n317 & n1171;
  assign n1173 = ~n1170 & ~n1172;
  assign n1174 = o0 & n1163;
  assign n1175 = n1162 & n1174;
  assign l9 = ~n1173 | n1175;
  assign n1177 = w & o0;
  assign n1178 = ~q0 & n1177;
  assign n1179 = ~n309 & ~n1178;
  assign n1180 = ~n307 & n1179;
  assign n1181 = ~d2 & ~n305;
  assign n1182 = ~n301 & n1181;
  assign n1183 = ~n1180 & ~n1182;
  assign n1184 = ~e2 & l4;
  assign n1185 = n319 & n1183;
  assign n1186 = n301 & ~n1184;
  assign n1187 = n1183 & n1186;
  assign n1188 = n323 & n1183;
  assign n1189 = n325 & n1183;
  assign n1190 = ~n0 & ~n1184;
  assign n1191 = n1183 & n1190;
  assign n1192 = n329 & n1183;
  assign n1193 = d2 & n317;
  assign n1194 = n1183 & n1193;
  assign n1195 = d2 & ~n1184;
  assign n1196 = n1183 & n1195;
  assign n1197 = d2 & n300;
  assign n1198 = n1183 & n1197;
  assign n1199 = ~n1196 & ~n1198;
  assign n1200 = ~n1194 & n1199;
  assign n1201 = ~n1192 & n1200;
  assign n1202 = ~n1191 & n1201;
  assign n1203 = ~n1189 & n1202;
  assign n1204 = ~n1188 & n1203;
  assign n1205 = ~n1187 & n1204;
  assign m7 = n1185 | ~n1205;
  assign n1207 = d3 & ~q0;
  assign n1208 = e3 & k4;
  assign n1209 = ~n392 & n1208;
  assign n1210 = n430 & n1209;
  assign n1211 = n426 & n1210;
  assign n1212 = o0 & n1207;
  assign n1213 = n413 & n1212;
  assign m8 = n1211 | n1213;
  assign n1215 = d4 & k4;
  assign n1216 = ~n386 & ~n392;
  assign n1217 = n1215 & n1216;
  assign n1218 = ~d4 & ~n798;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = ~g1 & ~q0;
  assign n1221 = n955 & n1111;
  assign n1222 = o0 & n1220;
  assign n1223 = n1219 & n1222;
  assign m9 = n1221 | n1223;
  assign n1225 = h1 & ~k4;
  assign n5 = n0 | ~n1225;
  assign n1227 = f1 & i4;
  assign n1228 = ~f1 & ~i4;
  assign n6 = n1227 | n1228;
  assign n1230 = x & o0;
  assign n1231 = ~q0 & n1230;
  assign n1232 = ~n309 & ~n1231;
  assign n1233 = ~n307 & n1232;
  assign n1234 = ~e2 & ~n305;
  assign n1235 = ~n301 & n1234;
  assign n1236 = ~n1233 & ~n1235;
  assign n1237 = ~f2 & l4;
  assign n1238 = n319 & n1236;
  assign n1239 = n301 & ~n1237;
  assign n1240 = n1236 & n1239;
  assign n1241 = n323 & n1236;
  assign n1242 = n325 & n1236;
  assign n1243 = ~n0 & ~n1237;
  assign n1244 = n1236 & n1243;
  assign n1245 = n329 & n1236;
  assign n1246 = e2 & n317;
  assign n1247 = n1236 & n1246;
  assign n1248 = e2 & ~n1237;
  assign n1249 = n1236 & n1248;
  assign n1250 = e2 & n300;
  assign n1251 = n1236 & n1250;
  assign n1252 = ~n1249 & ~n1251;
  assign n1253 = ~n1247 & n1252;
  assign n1254 = ~n1245 & n1253;
  assign n1255 = ~n1244 & n1254;
  assign n1256 = ~n1242 & n1255;
  assign n1257 = ~n1241 & n1256;
  assign n1258 = ~n1240 & n1257;
  assign n7 = n1238 | ~n1258;
  assign n1260 = e3 & ~q0;
  assign n1261 = f3 & k4;
  assign n1262 = ~n392 & n1261;
  assign n1263 = n430 & n1262;
  assign n1264 = n426 & n1263;
  assign n1265 = o0 & n1260;
  assign n1266 = n413 & n1265;
  assign n8 = n1264 | n1266;
  assign n1268 = ~d4 & k4;
  assign n1269 = n1216 & n1268;
  assign n1270 = ~e4 & k4;
  assign n1271 = ~d4 & n1270;
  assign n1272 = n1216 & n1271;
  assign n1273 = ~n317 & ~n1272;
  assign n1274 = n1220 & n1273;
  assign n1275 = o0 & n1274;
  assign n1276 = e4 & ~n1269;
  assign n9 = ~n1275 | n1276;
  assign n1278 = i1 & ~k4;
  assign o5 = n0 | ~n1278;
  assign n1280 = x3 & y3;
  assign n1281 = n296 & n1280;
  assign o6 = n299 & n1281;
  assign n1283 = y & o0;
  assign n1284 = ~q0 & n1283;
  assign n1285 = ~n309 & ~n1284;
  assign n1286 = ~n307 & n1285;
  assign n1287 = ~f2 & ~n305;
  assign n1288 = ~n301 & n1287;
  assign n1289 = ~n1286 & ~n1288;
  assign n1290 = ~g2 & l4;
  assign n1291 = n319 & n1289;
  assign n1292 = n301 & ~n1290;
  assign n1293 = n1289 & n1292;
  assign n1294 = n323 & n1289;
  assign n1295 = n325 & n1289;
  assign n1296 = ~n0 & ~n1290;
  assign n1297 = n1289 & n1296;
  assign n1298 = n329 & n1289;
  assign n1299 = f2 & n317;
  assign n1300 = n1289 & n1299;
  assign n1301 = f2 & ~n1290;
  assign n1302 = n1289 & n1301;
  assign n1303 = f2 & n300;
  assign n1304 = n1289 & n1303;
  assign n1305 = ~n1302 & ~n1304;
  assign n1306 = ~n1300 & n1305;
  assign n1307 = ~n1298 & n1306;
  assign n1308 = ~n1297 & n1307;
  assign n1309 = ~n1295 & n1308;
  assign n1310 = ~n1294 & n1309;
  assign n1311 = ~n1293 & n1310;
  assign o7 = n1291 | ~n1311;
  assign n1313 = f3 & ~q0;
  assign n1314 = g3 & k4;
  assign n1315 = ~n392 & n1314;
  assign n1316 = n430 & n1315;
  assign n1317 = n426 & n1316;
  assign n1318 = o0 & n1313;
  assign n1319 = n413 & n1318;
  assign o8 = n1317 | n1319;
  assign n1321 = e4 & k4;
  assign n1322 = ~d4 & n1321;
  assign n1323 = n1216 & n1322;
  assign n1324 = ~f4 & k4;
  assign n1325 = e4 & n1324;
  assign n1326 = ~d4 & ~n392;
  assign n1327 = ~n386 & n1326;
  assign n1328 = n1325 & n1327;
  assign n1329 = ~n317 & ~n1328;
  assign n1330 = n1220 & n1329;
  assign n1331 = o0 & n1330;
  assign n1332 = f4 & ~n1323;
  assign o9 = ~n1331 | n1332;
  assign n1334 = ~m0 & ~t3;
  assign n1335 = ~d3 & ~l3;
  assign n1336 = ~d3 & l0;
  assign n1337 = ~l0 & ~l3;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1335 & n1338;
  assign n1340 = ~d3 & ~l0;
  assign n1341 = l0 & ~l3;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = ~n1335 & n1342;
  assign n1344 = n1339 & n1343;
  assign n1345 = ~n1334 & n1344;
  assign n1346 = k0 & n1339;
  assign n1347 = ~n1334 & n1346;
  assign n1348 = ~m0 & ~n1334;
  assign n1349 = ~k0 & n1343;
  assign n1350 = ~n1334 & n1349;
  assign n1351 = ~n1348 & ~n1350;
  assign n1352 = ~n1347 & n1351;
  assign p4 = n1345 | ~n1352;
  assign n1354 = j1 & ~k4;
  assign p5 = n0 | ~n1354;
  assign n1356 = ~g4 & ~h4;
  assign n1357 = e4 & f4;
  assign n1358 = n1356 & n1357;
  assign n1359 = d4 & ~g1;
  assign n1360 = n1357 & n1359;
  assign n1361 = n1356 & n1360;
  assign n1362 = ~b1 & l1;
  assign n1363 = ~n1361 & n1362;
  assign n1364 = n1358 & ~n1361;
  assign n1365 = ~n4 & ~n1361;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1363 & n1366;
  assign n1368 = n370 & n1367;
  assign n1369 = n368 & n1367;
  assign n1370 = n366 & n1367;
  assign n1371 = n364 & n1367;
  assign n1372 = n1358 & n1367;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1370 & n1373;
  assign n1375 = ~n1369 & n1374;
  assign n1376 = ~n1368 & n1375;
  assign n1377 = n383 & ~n1358;
  assign n1378 = n384 & ~n1358;
  assign n1379 = ~n1376 & ~n1378;
  assign n1380 = ~n1377 & n1379;
  assign n1381 = ~q0 & n1380;
  assign p6 = o0 & n1381;
  assign n1383 = z & o0;
  assign n1384 = ~q0 & n1383;
  assign n1385 = ~n309 & ~n1384;
  assign n1386 = ~n307 & n1385;
  assign n1387 = ~g2 & ~n305;
  assign n1388 = ~n301 & n1387;
  assign n1389 = ~n1386 & ~n1388;
  assign n1390 = ~h2 & l4;
  assign n1391 = n319 & n1389;
  assign n1392 = n301 & ~n1390;
  assign n1393 = n1389 & n1392;
  assign n1394 = n323 & n1389;
  assign n1395 = n325 & n1389;
  assign n1396 = ~n0 & ~n1390;
  assign n1397 = n1389 & n1396;
  assign n1398 = n329 & n1389;
  assign n1399 = g2 & n317;
  assign n1400 = n1389 & n1399;
  assign n1401 = g2 & ~n1390;
  assign n1402 = n1389 & n1401;
  assign n1403 = g2 & n300;
  assign n1404 = n1389 & n1403;
  assign n1405 = ~n1402 & ~n1404;
  assign n1406 = ~n1400 & n1405;
  assign n1407 = ~n1398 & n1406;
  assign n1408 = ~n1397 & n1407;
  assign n1409 = ~n1395 & n1408;
  assign n1410 = ~n1394 & n1409;
  assign n1411 = ~n1393 & n1410;
  assign p7 = n1391 | ~n1411;
  assign n1413 = g3 & ~q0;
  assign n1414 = h3 & k4;
  assign n1415 = ~n392 & n1414;
  assign n1416 = n430 & n1415;
  assign n1417 = n426 & n1416;
  assign n1418 = o0 & n1413;
  assign n1419 = n413 & n1418;
  assign p8 = n1417 | n1419;
  assign n1421 = f4 & k4;
  assign n1422 = e4 & n1421;
  assign n1423 = n1327 & n1422;
  assign n1424 = ~n317 & ~n1423;
  assign n1425 = ~g1 & g4;
  assign n1426 = ~q0 & n1425;
  assign n1427 = ~q0 & n1216;
  assign n1428 = ~g4 & k4;
  assign n1429 = f4 & n1428;
  assign n1430 = ~d4 & e4;
  assign n1431 = ~g1 & n1430;
  assign n1432 = o0 & n1431;
  assign n1433 = n1429 & n1432;
  assign n1434 = m0 & n347;
  assign n1435 = m0 & n476;
  assign n1436 = ~n0 & ~n1435;
  assign n1437 = ~n1434 & n1436;
  assign n1438 = o0 & n1437;
  assign n1439 = n955 & n1438;
  assign n1440 = n1427 & n1433;
  assign n1441 = ~n317 & n1440;
  assign n1442 = ~n1439 & ~n1441;
  assign n1443 = o0 & n1426;
  assign n1444 = n1424 & n1443;
  assign p9 = ~n1442 | n1444;
  assign n1446 = ~m0 & ~s3;
  assign n1447 = ~c3 & ~k3;
  assign n1448 = ~c3 & l0;
  assign n1449 = ~k3 & ~l0;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = ~n1447 & n1450;
  assign n1452 = ~c3 & ~l0;
  assign n1453 = ~k3 & l0;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1447 & n1454;
  assign n1456 = n1451 & n1455;
  assign n1457 = ~n1446 & n1456;
  assign n1458 = k0 & n1451;
  assign n1459 = ~n1446 & n1458;
  assign n1460 = ~m0 & ~n1446;
  assign n1461 = ~k0 & n1455;
  assign n1462 = ~n1446 & n1461;
  assign n1463 = ~n1460 & ~n1462;
  assign n1464 = ~n1459 & n1463;
  assign q4 = n1457 | ~n1464;
  assign n1466 = k1 & ~k4;
  assign q5 = n0 | ~n1466;
  assign n1468 = c1 & e1;
  assign n1469 = d1 & e1;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n317 & n1470;
  assign n1472 = ~g1 & h1;
  assign n1473 = ~q0 & n1472;
  assign n1474 = ~e1 & n305;
  assign n1475 = ~d1 & n1474;
  assign n1476 = ~c1 & ~q0;
  assign n1477 = o0 & n1476;
  assign n1478 = ~n0 & n1477;
  assign n1479 = n1475 & n1478;
  assign n1480 = o0 & n1473;
  assign n1481 = ~n1471 & n1480;
  assign q6 = n1479 | n1481;
  assign n1483 = a0 & o0;
  assign n1484 = ~q0 & n1483;
  assign n1485 = ~n309 & ~n1484;
  assign n1486 = ~n307 & n1485;
  assign n1487 = ~h2 & ~n305;
  assign n1488 = ~n301 & n1487;
  assign n1489 = ~n1486 & ~n1488;
  assign n1490 = ~i2 & l4;
  assign n1491 = n319 & n1489;
  assign n1492 = n301 & ~n1490;
  assign n1493 = n1489 & n1492;
  assign n1494 = n323 & n1489;
  assign n1495 = n325 & n1489;
  assign n1496 = ~n0 & ~n1490;
  assign n1497 = n1489 & n1496;
  assign n1498 = n329 & n1489;
  assign n1499 = h2 & n317;
  assign n1500 = n1489 & n1499;
  assign n1501 = h2 & ~n1490;
  assign n1502 = n1489 & n1501;
  assign n1503 = h2 & n300;
  assign n1504 = n1489 & n1503;
  assign n1505 = ~n1502 & ~n1504;
  assign n1506 = ~n1500 & n1505;
  assign n1507 = ~n1498 & n1506;
  assign n1508 = ~n1497 & n1507;
  assign n1509 = ~n1495 & n1508;
  assign n1510 = ~n1494 & n1509;
  assign n1511 = ~n1493 & n1510;
  assign q7 = n1491 | ~n1511;
  assign n1513 = h3 & ~q0;
  assign n1514 = i3 & k4;
  assign n1515 = ~n392 & n1514;
  assign n1516 = n430 & n1515;
  assign n1517 = n426 & n1516;
  assign n1518 = o0 & n1513;
  assign n1519 = n413 & n1518;
  assign q8 = n1517 | n1519;
  assign n1521 = ~n392 & n1430;
  assign n1522 = ~n386 & n1521;
  assign n1523 = n1429 & n1522;
  assign n1524 = ~n317 & ~n1523;
  assign n1525 = ~g1 & h4;
  assign n1526 = ~q0 & n1525;
  assign n1527 = ~h4 & k4;
  assign n1528 = ~g4 & n1527;
  assign n1529 = ~d4 & n1357;
  assign n1530 = ~g1 & ~n392;
  assign n1531 = n1529 & n1530;
  assign n1532 = n1528 & n1531;
  assign n1533 = n430 & n1532;
  assign n1534 = ~n317 & n1533;
  assign n1535 = ~n1113 & ~n1534;
  assign n1536 = o0 & n1526;
  assign n1537 = n1524 & n1536;
  assign q9 = ~n1535 | n1537;
  assign n1539 = ~m0 & ~r3;
  assign n1540 = ~b3 & ~j3;
  assign n1541 = ~b3 & l0;
  assign n1542 = ~j3 & ~l0;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1540 & n1543;
  assign n1545 = ~b3 & ~l0;
  assign n1546 = ~j3 & l0;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1540 & n1547;
  assign n1549 = n1544 & n1548;
  assign n1550 = ~n1539 & n1549;
  assign n1551 = k0 & n1544;
  assign n1552 = ~n1539 & n1551;
  assign n1553 = ~m0 & ~n1539;
  assign n1554 = ~k0 & n1548;
  assign n1555 = ~n1539 & n1554;
  assign n1556 = ~n1553 & ~n1555;
  assign n1557 = ~n1552 & n1556;
  assign r4 = n1550 | ~n1557;
  assign n1559 = ~k4 & l1;
  assign r5 = n0 | ~n1559;
  assign n1561 = ~e1 & ~n0;
  assign n1562 = n305 & n1561;
  assign n1563 = ~i1 & ~n1562;
  assign n1564 = n362 & ~n1563;
  assign n1565 = ~n0 & n1474;
  assign n1566 = d1 & ~e1;
  assign n1567 = ~c1 & ~d1;
  assign n1568 = ~c1 & ~e1;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = ~n1566 & n1569;
  assign n1571 = n1565 & n1570;
  assign n1572 = n1564 & n1571;
  assign n1573 = n0 & n1565;
  assign n1574 = n1564 & n1573;
  assign n1575 = ~n305 & n1565;
  assign n1576 = n1564 & n1575;
  assign n1577 = ~g1 & n1570;
  assign n1578 = n1564 & n1577;
  assign n1579 = ~g1 & ~n305;
  assign n1580 = n1564 & n1579;
  assign n1581 = ~g1 & n0;
  assign n1582 = n1564 & n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584 = ~n1578 & n1583;
  assign n1585 = ~n1576 & n1584;
  assign n1586 = ~n1574 & n1585;
  assign r6 = n1572 | ~n1586;
  assign n1588 = b0 & o0;
  assign n1589 = ~q0 & n1588;
  assign n1590 = ~n309 & ~n1589;
  assign n1591 = ~n307 & n1590;
  assign n1592 = ~i2 & ~n305;
  assign n1593 = ~n301 & n1592;
  assign n1594 = ~n1591 & ~n1593;
  assign n1595 = ~j2 & l4;
  assign n1596 = n319 & n1594;
  assign n1597 = n301 & ~n1595;
  assign n1598 = n1594 & n1597;
  assign n1599 = n323 & n1594;
  assign n1600 = n325 & n1594;
  assign n1601 = ~n0 & ~n1595;
  assign n1602 = n1594 & n1601;
  assign n1603 = n329 & n1594;
  assign n1604 = i2 & n317;
  assign n1605 = n1594 & n1604;
  assign n1606 = i2 & ~n1595;
  assign n1607 = n1594 & n1606;
  assign n1608 = i2 & n300;
  assign n1609 = n1594 & n1608;
  assign n1610 = ~n1607 & ~n1609;
  assign n1611 = ~n1605 & n1610;
  assign n1612 = ~n1603 & n1611;
  assign n1613 = ~n1602 & n1612;
  assign n1614 = ~n1600 & n1613;
  assign n1615 = ~n1599 & n1614;
  assign n1616 = ~n1598 & n1615;
  assign r7 = n1596 | ~n1616;
  assign n1618 = i3 & ~q0;
  assign n1619 = j3 & k4;
  assign n1620 = ~n392 & n1619;
  assign n1621 = n430 & n1620;
  assign n1622 = n426 & n1621;
  assign n1623 = o0 & n1618;
  assign n1624 = n413 & n1623;
  assign r8 = n1622 | n1624;
  assign n1626 = ~q0 & ~n300;
  assign n1627 = o0 & n1626;
  assign n1628 = i4 & n1;
  assign n1629 = n1627 & ~n1628;
  assign n1630 = i4 & l4;
  assign n1631 = n1629 & n1630;
  assign n1632 = l4 & n1;
  assign n1633 = n1629 & n1632;
  assign r9 = n1631 | n1633;
  assign n1635 = ~m0 & ~q3;
  assign n1636 = ~a3 & ~i3;
  assign n1637 = ~a3 & l0;
  assign n1638 = ~i3 & ~l0;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = ~n1636 & n1639;
  assign n1641 = ~a3 & ~l0;
  assign n1642 = ~i3 & l0;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1636 & n1643;
  assign n1645 = n1640 & n1644;
  assign n1646 = ~n1635 & n1645;
  assign n1647 = k0 & n1640;
  assign n1648 = ~n1635 & n1647;
  assign n1649 = ~m0 & ~n1635;
  assign n1650 = ~k0 & n1644;
  assign n1651 = ~n1635 & n1650;
  assign n1652 = ~n1649 & ~n1651;
  assign n1653 = ~n1648 & n1652;
  assign s4 = n1646 | ~n1653;
  assign n1655 = ~a4 & n299;
  assign n1656 = n1108 & n1655;
  assign n1657 = f1 & ~i4;
  assign n1658 = ~f1 & i4;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = n1656 & n1659;
  assign n1661 = ~n1655 & n1656;
  assign n1662 = ~n1108 & n1656;
  assign n1663 = n1 & n1659;
  assign n1664 = n1 & ~n1655;
  assign n1665 = n1 & ~n1108;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1663 & n1666;
  assign n1668 = ~n1662 & n1667;
  assign n1669 = ~n1661 & n1668;
  assign s5 = n1660 | ~n1669;
  assign n1671 = ~j1 & ~n1562;
  assign n1672 = n362 & ~n1671;
  assign n1673 = ~d1 & ~e1;
  assign n1674 = c1 & ~e1;
  assign n1675 = ~n1567 & ~n1674;
  assign n1676 = ~n1673 & n1675;
  assign n1677 = n1565 & n1676;
  assign n1678 = n1672 & n1677;
  assign n1679 = n1573 & n1672;
  assign n1680 = n1575 & n1672;
  assign n1681 = ~g1 & n1676;
  assign n1682 = n1672 & n1681;
  assign n1683 = n1579 & n1672;
  assign n1684 = n1581 & n1672;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1682 & n1685;
  assign n1687 = ~n1680 & n1686;
  assign n1688 = ~n1679 & n1687;
  assign s6 = n1678 | ~n1688;
  assign n1690 = c0 & o0;
  assign n1691 = ~q0 & n1690;
  assign n1692 = ~n309 & ~n1691;
  assign n1693 = ~n307 & n1692;
  assign n1694 = ~j2 & ~n305;
  assign n1695 = ~n301 & n1694;
  assign n1696 = ~n1693 & ~n1695;
  assign n1697 = ~k2 & l4;
  assign n1698 = n319 & n1696;
  assign n1699 = n301 & ~n1697;
  assign n1700 = n1696 & n1699;
  assign n1701 = n323 & n1696;
  assign n1702 = n325 & n1696;
  assign n1703 = ~n0 & ~n1697;
  assign n1704 = n1696 & n1703;
  assign n1705 = n329 & n1696;
  assign n1706 = j2 & n317;
  assign n1707 = n1696 & n1706;
  assign n1708 = j2 & ~n1697;
  assign n1709 = n1696 & n1708;
  assign n1710 = j2 & n300;
  assign n1711 = n1696 & n1710;
  assign n1712 = ~n1709 & ~n1711;
  assign n1713 = ~n1707 & n1712;
  assign n1714 = ~n1705 & n1713;
  assign n1715 = ~n1704 & n1714;
  assign n1716 = ~n1702 & n1715;
  assign n1717 = ~n1701 & n1716;
  assign n1718 = ~n1700 & n1717;
  assign s7 = n1698 | ~n1718;
  assign n1720 = j3 & ~q0;
  assign n1721 = k3 & k4;
  assign n1722 = ~n392 & n1721;
  assign n1723 = n430 & n1722;
  assign n1724 = n426 & n1723;
  assign n1725 = o0 & n1720;
  assign n1726 = n413 & n1725;
  assign s8 = n1724 | n1726;
  assign n1728 = ~i1 & n304;
  assign n1729 = ~j1 & t0;
  assign n1730 = n304 & n1729;
  assign n1731 = n304 & ~n392;
  assign n1732 = ~n393 & ~n1731;
  assign n1733 = ~n386 & ~n1732;
  assign n1734 = ~n398 & n1733;
  assign n1735 = k4 & n4;
  assign n1736 = n1734 & n1735;
  assign n1737 = ~h1 & ~u0;
  assign n1738 = n1728 & n1737;
  assign n1739 = i1 & ~n1730;
  assign n1740 = n1736 & ~n1739;
  assign n1741 = ~n1738 & n1740;
  assign n1742 = ~i1 & s0;
  assign n1743 = n401 & n1742;
  assign n1744 = ~k1 & ~w0;
  assign n1745 = ~l1 & ~v0;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n304 & n1746;
  assign n1748 = n1743 & n1747;
  assign n1749 = n1741 & n1748;
  assign n1750 = ~n302 & n1743;
  assign n1751 = n1741 & n1750;
  assign n1752 = h1 & n1743;
  assign n1753 = n1741 & n1752;
  assign n1754 = ~h1 & ~n302;
  assign n1755 = n1741 & n1754;
  assign n1756 = ~h1 & n1747;
  assign n1757 = n1741 & n1756;
  assign n1758 = ~n1755 & ~n1757;
  assign n1759 = ~n1753 & n1758;
  assign n1760 = ~n1751 & n1759;
  assign n1761 = ~n1749 & n1760;
  assign n1762 = ~g1 & j4;
  assign n1763 = ~q0 & n1762;
  assign n1764 = ~n386 & n1530;
  assign n1765 = ~j4 & n1735;
  assign n1766 = n362 & n1765;
  assign n1767 = n1764 & n1766;
  assign n1768 = n797 & n1767;
  assign n1769 = o0 & n1763;
  assign n1770 = n1761 & n1769;
  assign s9 = n1768 | n1770;
  assign n1772 = ~k1 & ~n1562;
  assign n1773 = n362 & ~n1772;
  assign n1774 = n1569 & ~n1673;
  assign n1775 = n1565 & n1774;
  assign n1776 = n1773 & n1775;
  assign n1777 = n1573 & n1773;
  assign n1778 = n1575 & n1773;
  assign n1779 = ~g1 & n1774;
  assign n1780 = n1773 & n1779;
  assign n1781 = n1579 & n1773;
  assign n1782 = n1581 & n1773;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1780 & n1783;
  assign n1785 = ~n1778 & n1784;
  assign n1786 = ~n1777 & n1785;
  assign t6 = n1776 | ~n1786;
  assign n1788 = ~l2 & l4;
  assign n1789 = i & n347;
  assign n1790 = a & l0;
  assign n1791 = a & ~k0;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1789 & n1792;
  assign n1794 = ~k2 & ~n301;
  assign n1795 = ~n354 & n1794;
  assign n1796 = ~n300 & n1788;
  assign n1797 = ~n345 & n1796;
  assign n1798 = n345 & n1793;
  assign n1799 = ~n1795 & ~n1798;
  assign n1800 = ~n1797 & n1799;
  assign t7 = n362 & n1800;
  assign n1802 = k3 & ~q0;
  assign n1803 = k4 & l3;
  assign n1804 = ~n392 & n1803;
  assign n1805 = n430 & n1804;
  assign n1806 = n426 & n1805;
  assign n1807 = o0 & n1802;
  assign n1808 = n413 & n1807;
  assign t8 = n1806 | n1808;
  assign n1810 = m1 & ~q0;
  assign n1811 = o0 & n1810;
  assign n1812 = n1166 & n1811;
  assign t9 = n299 & n1812;
  assign n1814 = n362 & ~n1562;
  assign n1815 = ~d1 & n305;
  assign n1816 = ~c1 & ~n0;
  assign n1817 = n1815 & n1816;
  assign n1818 = ~g1 & l1;
  assign n1819 = n1814 & n1818;
  assign n1820 = n1814 & n1817;
  assign u6 = n1819 | n1820;
  assign n1822 = l4 & ~m2;
  assign n1823 = j & n347;
  assign n1824 = b & l0;
  assign n1825 = b & ~k0;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1823 & n1826;
  assign n1828 = ~l2 & ~n301;
  assign n1829 = ~n354 & n1828;
  assign n1830 = ~n300 & n1822;
  assign n1831 = ~n345 & n1830;
  assign n1832 = n345 & n1827;
  assign n1833 = ~n1829 & ~n1832;
  assign n1834 = ~n1831 & n1833;
  assign u7 = n362 & n1834;
  assign n1836 = l3 & ~q0;
  assign n1837 = k4 & m3;
  assign n1838 = ~n392 & n1837;
  assign n1839 = n430 & n1838;
  assign n1840 = n426 & n1839;
  assign n1841 = o0 & n1836;
  assign n1842 = n413 & n1841;
  assign u8 = n1840 | n1842;
  assign u9 = m1 & n1627;
  assign n1845 = ~e3 & n283;
  assign n1846 = ~e3 & n285;
  assign n1847 = m0 & ~n1846;
  assign n1848 = ~n1845 & n1847;
  assign n1849 = n283 & n1848;
  assign n1850 = n285 & n1848;
  assign n1851 = m3 & n1848;
  assign n1852 = ~n1850 & ~n1851;
  assign v4 = n1849 | ~n1852;
  assign n1854 = m1 & n1380;
  assign n1855 = n362 & ~n1854;
  assign n1856 = ~n0 & p0;
  assign n1857 = n1855 & n1856;
  assign n1858 = m1 & n1855;
  assign v6 = n1857 | n1858;
  assign n1860 = l4 & ~n2;
  assign n1861 = k & n347;
  assign n1862 = c & l0;
  assign n1863 = c & ~k0;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = ~n1861 & n1864;
  assign n1866 = ~m2 & ~n301;
  assign n1867 = ~n354 & n1866;
  assign n1868 = ~n300 & n1860;
  assign n1869 = ~n345 & n1868;
  assign n1870 = n345 & n1865;
  assign n1871 = ~n1867 & ~n1870;
  assign n1872 = ~n1869 & n1871;
  assign v7 = n362 & n1872;
  assign n1874 = m3 & ~q0;
  assign n1875 = k4 & n3;
  assign n1876 = ~n392 & n1875;
  assign n1877 = n430 & n1876;
  assign n1878 = n426 & n1877;
  assign n1879 = o0 & n1874;
  assign n1880 = n413 & n1879;
  assign v8 = n1878 | n1880;
  assign n1882 = ~a1 & k1;
  assign n1883 = ~n392 & ~n1882;
  assign n1884 = ~n1362 & n1883;
  assign n1885 = y0 & z0;
  assign n1886 = n1884 & n1885;
  assign n1887 = ~i1 & z0;
  assign n1888 = n1884 & n1887;
  assign n1889 = ~j1 & y0;
  assign n1890 = n1884 & n1889;
  assign n1891 = n302 & n1884;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = ~n1888 & n1892;
  assign n1894 = ~n1886 & n1893;
  assign n1895 = n4 & ~n1894;
  assign n1896 = ~n384 & n1895;
  assign n1897 = n386 & ~n1896;
  assign n1898 = n362 & ~n1897;
  assign n1899 = n1896 & n1898;
  assign n1900 = n1380 & n1898;
  assign v9 = n1899 | n1900;
  assign n1902 = ~f3 & n283;
  assign n1903 = ~f3 & n285;
  assign n1904 = m0 & ~n1903;
  assign n1905 = ~n1902 & n1904;
  assign n1906 = n283 & n1905;
  assign n1907 = n285 & n1905;
  assign n1908 = n3 & n1905;
  assign n1909 = ~n1907 & ~n1908;
  assign w4 = n1906 | ~n1909;
  assign n1911 = j0 & o0;
  assign n1912 = ~q0 & n1911;
  assign n1913 = ~n309 & ~n1912;
  assign n1914 = ~n307 & n1913;
  assign n1915 = ~n1 & ~n305;
  assign n1916 = ~n301 & n1915;
  assign n1917 = ~n1914 & ~n1916;
  assign n1918 = l4 & ~o1;
  assign n1919 = n319 & n1917;
  assign n1920 = n301 & ~n1918;
  assign n1921 = n1917 & n1920;
  assign n1922 = n323 & n1917;
  assign n1923 = n325 & n1917;
  assign n1924 = ~n0 & ~n1918;
  assign n1925 = n1917 & n1924;
  assign n1926 = n329 & n1917;
  assign n1927 = n1 & n317;
  assign n1928 = n1917 & n1927;
  assign n1929 = n1 & ~n1918;
  assign n1930 = n1917 & n1929;
  assign n1931 = n1 & n300;
  assign n1932 = n1917 & n1931;
  assign n1933 = ~n1930 & ~n1932;
  assign n1934 = ~n1928 & n1933;
  assign n1935 = ~n1926 & n1934;
  assign n1936 = ~n1925 & n1935;
  assign n1937 = ~n1923 & n1936;
  assign n1938 = ~n1922 & n1937;
  assign n1939 = ~n1921 & n1938;
  assign w6 = n1919 | ~n1939;
  assign n1941 = l4 & ~o2;
  assign n1942 = l & n347;
  assign n1943 = d & l0;
  assign n1944 = d & ~k0;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = ~n1942 & n1945;
  assign n1947 = ~n2 & ~n301;
  assign n1948 = ~n354 & n1947;
  assign n1949 = ~n300 & n1941;
  assign n1950 = ~n345 & n1949;
  assign n1951 = n345 & n1946;
  assign n1952 = ~n1948 & ~n1951;
  assign n1953 = ~n1950 & n1952;
  assign w7 = n362 & n1953;
  assign n1955 = n3 & ~q0;
  assign n1956 = k4 & o3;
  assign n1957 = ~n392 & n1956;
  assign n1958 = n430 & n1957;
  assign n1959 = n426 & n1958;
  assign n1960 = o0 & n1955;
  assign n1961 = n413 & n1960;
  assign w8 = n1959 | n1961;
  assign w9 = k4 & n430;
  assign n1964 = ~g3 & n283;
  assign n1965 = ~g3 & n285;
  assign n1966 = m0 & ~n1965;
  assign n1967 = ~n1964 & n1966;
  assign n1968 = n283 & n1967;
  assign n1969 = n285 & n1967;
  assign n1970 = o3 & n1967;
  assign n1971 = ~n1969 & ~n1970;
  assign x4 = n1968 | ~n1971;
  assign x5 = ~h1 | ~n294;
  assign n1974 = i0 & o0;
  assign n1975 = ~q0 & n1974;
  assign n1976 = ~n309 & ~n1975;
  assign n1977 = ~n307 & n1976;
  assign n1978 = ~o1 & ~n305;
  assign n1979 = ~n301 & n1978;
  assign n1980 = ~n1977 & ~n1979;
  assign n1981 = l4 & ~p1;
  assign n1982 = n319 & n1980;
  assign n1983 = n301 & ~n1981;
  assign n1984 = n1980 & n1983;
  assign n1985 = n323 & n1980;
  assign n1986 = n325 & n1980;
  assign n1987 = ~n0 & ~n1981;
  assign n1988 = n1980 & n1987;
  assign n1989 = n329 & n1980;
  assign n1990 = o1 & n317;
  assign n1991 = n1980 & n1990;
  assign n1992 = o1 & ~n1981;
  assign n1993 = n1980 & n1992;
  assign n1994 = o1 & n300;
  assign n1995 = n1980 & n1994;
  assign n1996 = ~n1993 & ~n1995;
  assign n1997 = ~n1991 & n1996;
  assign n1998 = ~n1989 & n1997;
  assign n1999 = ~n1988 & n1998;
  assign n2000 = ~n1986 & n1999;
  assign n2001 = ~n1985 & n2000;
  assign n2002 = ~n1984 & n2001;
  assign x6 = n1982 | ~n2002;
  assign n2004 = l4 & ~p2;
  assign n2005 = m & n347;
  assign n2006 = e & l0;
  assign n2007 = e & ~k0;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~n2005 & n2008;
  assign n2010 = ~o2 & ~n301;
  assign n2011 = ~n354 & n2010;
  assign n2012 = ~n300 & n2004;
  assign n2013 = ~n345 & n2012;
  assign n2014 = n345 & n2009;
  assign n2015 = ~n2011 & ~n2014;
  assign n2016 = ~n2013 & n2015;
  assign x7 = n362 & n2016;
  assign n2018 = o3 & ~q0;
  assign n2019 = k4 & p3;
  assign n2020 = ~n392 & n2019;
  assign n2021 = n430 & n2020;
  assign n2022 = n426 & n2021;
  assign n2023 = o0 & n2018;
  assign n2024 = n413 & n2023;
  assign x8 = n2022 | n2024;
  assign n2026 = ~h3 & n283;
  assign n2027 = ~h3 & n285;
  assign n2028 = m0 & ~n2027;
  assign n2029 = ~n2026 & n2028;
  assign n2030 = n283 & n2029;
  assign n2031 = n285 & n2029;
  assign n2032 = p3 & n2029;
  assign n2033 = ~n2031 & ~n2032;
  assign y4 = n2030 | ~n2033;
  assign y5 = ~i1 | ~n294;
  assign n2036 = h0 & o0;
  assign n2037 = ~q0 & n2036;
  assign n2038 = ~n309 & ~n2037;
  assign n2039 = ~n307 & n2038;
  assign n2040 = ~p1 & ~n305;
  assign n2041 = ~n301 & n2040;
  assign n2042 = ~n2039 & ~n2041;
  assign n2043 = l4 & ~q1;
  assign n2044 = n319 & n2042;
  assign n2045 = n301 & ~n2043;
  assign n2046 = n2042 & n2045;
  assign n2047 = n323 & n2042;
  assign n2048 = n325 & n2042;
  assign n2049 = ~n0 & ~n2043;
  assign n2050 = n2042 & n2049;
  assign n2051 = n329 & n2042;
  assign n2052 = p1 & n317;
  assign n2053 = n2042 & n2052;
  assign n2054 = p1 & ~n2043;
  assign n2055 = n2042 & n2054;
  assign n2056 = p1 & n300;
  assign n2057 = n2042 & n2056;
  assign n2058 = ~n2055 & ~n2057;
  assign n2059 = ~n2053 & n2058;
  assign n2060 = ~n2051 & n2059;
  assign n2061 = ~n2050 & n2060;
  assign n2062 = ~n2048 & n2061;
  assign n2063 = ~n2047 & n2062;
  assign n2064 = ~n2046 & n2063;
  assign y6 = n2044 | ~n2064;
  assign n2066 = l4 & ~q2;
  assign n2067 = n & n347;
  assign n2068 = f & l0;
  assign n2069 = f & ~k0;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2067 & n2070;
  assign n2072 = ~p2 & ~n301;
  assign n2073 = ~n354 & n2072;
  assign n2074 = ~n300 & n2066;
  assign n2075 = ~n345 & n2074;
  assign n2076 = n345 & n2071;
  assign n2077 = ~n2073 & ~n2076;
  assign n2078 = ~n2075 & n2077;
  assign y7 = n362 & n2078;
  assign n2080 = p3 & ~q0;
  assign n2081 = k4 & q3;
  assign n2082 = ~n392 & n2081;
  assign n2083 = n430 & n2082;
  assign n2084 = n426 & n2083;
  assign n2085 = o0 & n2080;
  assign n2086 = n413 & n2085;
  assign y8 = n2084 | n2086;
  assign n2088 = ~i3 & n283;
  assign n2089 = ~i3 & n285;
  assign n2090 = m0 & ~n2089;
  assign n2091 = ~n2088 & n2090;
  assign n2092 = n283 & n2091;
  assign n2093 = n285 & n2091;
  assign n2094 = q3 & n2091;
  assign n2095 = ~n2093 & ~n2094;
  assign z4 = n2092 | ~n2095;
  assign z5 = ~j1 | ~n294;
  assign n2098 = g0 & o0;
  assign n2099 = ~q0 & n2098;
  assign n2100 = ~n309 & ~n2099;
  assign n2101 = ~n307 & n2100;
  assign n2102 = ~q1 & ~n305;
  assign n2103 = ~n301 & n2102;
  assign n2104 = ~n2101 & ~n2103;
  assign n2105 = l4 & ~r1;
  assign n2106 = n319 & n2104;
  assign n2107 = n301 & ~n2105;
  assign n2108 = n2104 & n2107;
  assign n2109 = n323 & n2104;
  assign n2110 = n325 & n2104;
  assign n2111 = ~n0 & ~n2105;
  assign n2112 = n2104 & n2111;
  assign n2113 = n329 & n2104;
  assign n2114 = q1 & n317;
  assign n2115 = n2104 & n2114;
  assign n2116 = q1 & ~n2105;
  assign n2117 = n2104 & n2116;
  assign n2118 = q1 & n300;
  assign n2119 = n2104 & n2118;
  assign n2120 = ~n2117 & ~n2119;
  assign n2121 = ~n2115 & n2120;
  assign n2122 = ~n2113 & n2121;
  assign n2123 = ~n2112 & n2122;
  assign n2124 = ~n2110 & n2123;
  assign n2125 = ~n2109 & n2124;
  assign n2126 = ~n2108 & n2125;
  assign z6 = n2106 | ~n2126;
  assign n2128 = l4 & ~r2;
  assign n2129 = o & n347;
  assign n2130 = g & l0;
  assign n2131 = g & ~k0;
  assign n2132 = ~n2130 & ~n2131;
  assign n2133 = ~n2129 & n2132;
  assign n2134 = ~q2 & ~n301;
  assign n2135 = ~n354 & n2134;
  assign n2136 = ~n300 & n2128;
  assign n2137 = ~n345 & n2136;
  assign n2138 = n345 & n2133;
  assign n2139 = ~n2135 & ~n2138;
  assign n2140 = ~n2137 & n2139;
  assign z7 = n362 & n2140;
  assign n2142 = ~q0 & q3;
  assign n2143 = k4 & r3;
  assign n2144 = ~n392 & n2143;
  assign n2145 = n430 & n2144;
  assign n2146 = n426 & n2145;
  assign n2147 = o0 & n2142;
  assign n2148 = n413 & n2147;
  assign z8 = n2146 | n2148;
  assign h6 = ~h1;
  assign i6 = ~i1;
  assign j6 = ~j1;
  assign k6 = ~k1;
  assign l6 = ~l1;
  assign o4 = ~g1;
  assign m5 = m4;
  assign m6 = k4;
  assign t4 = u3;
  assign t5 = s5;
  assign u4 = v3;
  assign u5 = s5;
  assign v5 = s5;
  assign w5 = s5;
endmodule


