// Benchmark "rot" written by ABC on Tue May 16 16:07:52 2017

module rot ( 
    z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r,
    s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4, c0, c1,
    c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2, f3, g0,
    g1, g2, g3, h0, h1, h2, h3, i0, i1, i2, i3, j0, j1, j2, j3, k0, k1, k2,
    k3, l0, l1, l2, l3, m0, m1, m2, m3, n0, n1, n2, n3, o0, o1, o2, o3, p0,
    p1, p2, p3, q0, q1, q2, q3, r0, r1, r2, r3, s0, s1, s2, s3, t0, t1, t2,
    t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2, w3, x0, x1, x2, x3, y0,
    y1, y2, y3,
    z4, z5, z6, z7, a5, a6, a7, a8, b5, b6, b7, b8, c5, c6, c7, c8, d5, d6,
    d7, d8, e5, e6, e7, e8, f4, f5, f6, f7, f8, g4, g5, g6, g7, g8, h4, h5,
    h6, h7, h8, i4, i5, i6, i7, j4, j5, j6, j7, k4, k5, k6, k7, l4, l5, l6,
    l7, m4, m5, m6, m7, n4, n5, n6, n7, o4, o5, o6, o7, p4, p5, p6, p7, q4,
    q5, q6, q7, r4, r5, r6, r7, s4, s5, s6, s7, t4, t5, t6, t7, u4, u5, u6,
    u7, v4, v5, v6, v7, w4, w5, w6, w7, x4, x5, x6, x7, y4, y5, y6, y7  );
  input  z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p,
    q, r, s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4,
    c0, c1, c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2,
    f3, g0, g1, g2, g3, h0, h1, h2, h3, i0, i1, i2, i3, j0, j1, j2, j3, k0,
    k1, k2, k3, l0, l1, l2, l3, m0, m1, m2, m3, n0, n1, n2, n3, o0, o1, o2,
    o3, p0, p1, p2, p3, q0, q1, q2, q3, r0, r1, r2, r3, s0, s1, s2, s3, t0,
    t1, t2, t3, u0, u1, u2, u3, v0, v1, v2, v3, w0, w1, w2, w3, x0, x1, x2,
    x3, y0, y1, y2, y3;
  output z4, z5, z6, z7, a5, a6, a7, a8, b5, b6, b7, b8, c5, c6, c7, c8, d5,
    d6, d7, d8, e5, e6, e7, e8, f4, f5, f6, f7, f8, g4, g5, g6, g7, g8, h4,
    h5, h6, h7, h8, i4, i5, i6, i7, j4, j5, j6, j7, k4, k5, k6, k7, l4, l5,
    l6, l7, m4, m5, m6, m7, n4, n5, n6, n7, o4, o5, o6, o7, p4, p5, p6, p7,
    q4, q5, q6, q7, r4, r5, r6, r7, s4, s5, s6, s7, t4, t5, t6, t7, u4, u5,
    u6, u7, v4, v5, v6, v7, w4, w5, w6, w7, x4, x5, x6, x7, y4, y5, y6, y7;
  wire n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n290, n291,
    n294, n295, n297, n298, n299, n300, n301, n303, n305, n306, n308, n309,
    n310, n311, n313, n314, n316, n317, n318, n319, n320, n322, n323, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n374,
    n376, n377, n378, n379, n380, n381, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n425, n426,
    n428, n430, n431, n432, n435, n436, n437, n438, n440, n441, n443, n444,
    n446, n448, n449, n451, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n479, n481, n482, n483, n484, n485, n487, n488, n489,
    n490, n491, n493, n494, n496, n497, n498, n499, n500, n501, n502, n504,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n544, n545, n546, n547, n548, n549, n551, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n568, n569, n571, n572, n573,
    n574, n575, n576, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n715, n717, n718, n719, n720, n721, n722,
    n724, n725, n726, n728, n729, n730, n734, n735, n736, n737, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n766, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n849, n850, n851,
    n852, n853, n854, n855, n856, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1002, n1003, n1004, n1005, n1006, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1056, n1057, n1058, n1059, n1060,
    n1061, n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1149, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1160, n1161, n1162, n1163, n1164, n1166,
    n1167, n1168, n1170, n1171, n1172, n1174, n1175, n1176, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1212, n1213, n1214, n1215, n1216, n1218, n1219, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1275, n1276, n1277,
    n1278, n1279, n1280, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1292, n1293, n1294, n1296, n1297, n1298, n1299, n1301, n1303;
  assign z4 = b4 & v0;
  assign n244 = ~h0 & t0;
  assign n245 = n3 & n244;
  assign n246 = ~m & ~d0;
  assign n247 = ~w2 & n246;
  assign n248 = x2 & n247;
  assign n249 = ~h0 & n248;
  assign n250 = u2 & n249;
  assign n251 = ~s0 & n250;
  assign n252 = ~k & d0;
  assign n253 = ~w2 & n252;
  assign n254 = x2 & n253;
  assign n255 = ~h0 & n254;
  assign n256 = u2 & n255;
  assign n257 = ~s0 & n256;
  assign n258 = ~u & n248;
  assign n259 = u2 & n258;
  assign n260 = s0 & n259;
  assign n261 = ~u & n254;
  assign n262 = u2 & n261;
  assign n263 = s0 & n262;
  assign n264 = ~h & u3;
  assign n265 = ~h0 & n264;
  assign n266 = u2 & n265;
  assign n267 = ~s0 & n266;
  assign n268 = ~u & n264;
  assign n269 = u2 & n268;
  assign n270 = s0 & n269;
  assign n271 = ~i & u3;
  assign n272 = ~l & ~d0;
  assign n273 = ~j & d0;
  assign n274 = g & ~n273;
  assign n275 = ~n272 & n274;
  assign n276 = ~n271 & n275;
  assign n277 = ~n270 & n276;
  assign n278 = ~n267 & n277;
  assign n279 = ~n263 & n278;
  assign n280 = ~n260 & n279;
  assign n281 = ~n257 & n280;
  assign n282 = ~n251 & n281;
  assign n283 = m2 & x1;
  assign n284 = y1 & n283;
  assign n285 = w2 & n282;
  assign n286 = w2 & ~x2;
  assign n287 = x2 & ~n284;
  assign n288 = ~n286 & ~n287;
  assign d8 = n285 | ~n288;
  assign n290 = ~i2 & ~k2;
  assign n291 = ~d8 & n290;
  assign z5 = n245 | ~n291;
  assign z6 = ~z0 & ~y0;
  assign n294 = m & d0;
  assign n295 = k & ~d0;
  assign z7 = n294 | n295;
  assign n297 = ~x & e0;
  assign n298 = y & n297;
  assign n299 = x & n0;
  assign n300 = ~y & n0;
  assign n301 = ~n299 & ~n300;
  assign a6 = n298 | ~n301;
  assign n303 = ~n282 & n284;
  assign a8 = c4 | n303;
  assign n305 = ~c1 & d1;
  assign n306 = c1 & ~d1;
  assign b5 = n305 | n306;
  assign n308 = m2 & q2;
  assign n309 = m1 & m2;
  assign n310 = m2 & r0;
  assign n311 = ~n309 & ~n310;
  assign b6 = n308 | ~n311;
  assign n313 = ~w2 & x2;
  assign n314 = n284 & n313;
  assign b8 = n282 & n314;
  assign n316 = c1 & d1;
  assign n317 = ~e1 & n316;
  assign n318 = ~d1 & e1;
  assign n319 = ~c1 & e1;
  assign n320 = ~n318 & ~n319;
  assign c5 = n317 | ~n320;
  assign n322 = w1 & x1;
  assign n323 = ~y1 & n322;
  assign c6 = m2 & n323;
  assign n325 = ~f2 & ~g2;
  assign n326 = h2 & n325;
  assign n327 = f2 & ~g2;
  assign n328 = ~h2 & n327;
  assign n329 = ~n326 & ~n328;
  assign n330 = ~p1 & r1;
  assign n331 = ~s1 & n330;
  assign n332 = l2 & n331;
  assign n333 = o2 & n332;
  assign n334 = ~n329 & n333;
  assign n335 = h2 & n334;
  assign n336 = ~p1 & ~r1;
  assign n337 = s1 & n336;
  assign n338 = l2 & n337;
  assign n339 = o2 & n338;
  assign n340 = ~n329 & n339;
  assign n341 = h2 & n340;
  assign n342 = f2 & n334;
  assign n343 = f2 & n340;
  assign n344 = z1 & n331;
  assign n345 = o2 & n344;
  assign n346 = h2 & n345;
  assign n347 = z1 & n337;
  assign n348 = o2 & n347;
  assign n349 = h2 & n348;
  assign n350 = f2 & n345;
  assign n351 = f2 & n348;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~n349 & n352;
  assign n354 = ~n346 & n353;
  assign n355 = ~n343 & n354;
  assign n356 = ~n342 & n355;
  assign n357 = ~n341 & n356;
  assign n358 = ~n335 & n357;
  assign n359 = q & l2;
  assign n360 = p2 & n359;
  assign n361 = q2 & n360;
  assign n362 = n358 & ~n361;
  assign n363 = o1 & n362;
  assign n364 = ~y3 & n363;
  assign n365 = ~s1 & ~n361;
  assign n366 = o1 & n365;
  assign n367 = ~y3 & n366;
  assign n368 = m1 & ~n361;
  assign n369 = n358 & n368;
  assign n370 = ~s1 & n368;
  assign n371 = ~n369 & ~n370;
  assign n372 = ~n367 & n371;
  assign c7 = n364 | ~n372;
  assign n374 = w2 & ~n284;
  assign c8 = ~a4 | n374;
  assign n376 = n & ~p;
  assign n377 = q & n376;
  assign n378 = ~c1 & ~d1;
  assign n379 = ~e1 & n378;
  assign n380 = l2 & n379;
  assign n381 = l2 & ~n377;
  assign d5 = n380 | n381;
  assign n383 = o1 & n369;
  assign n384 = ~y3 & n383;
  assign n385 = o1 & n370;
  assign n386 = ~y3 & n385;
  assign n387 = q2 & ~n361;
  assign n388 = o1 & n387;
  assign n389 = ~y3 & n388;
  assign n390 = p2 & ~n361;
  assign n391 = o1 & n390;
  assign n392 = ~y3 & n391;
  assign n393 = ~l2 & ~n361;
  assign n394 = o1 & n393;
  assign n395 = ~y3 & n394;
  assign n396 = ~q & ~n361;
  assign n397 = o1 & n396;
  assign n398 = ~y3 & n397;
  assign n399 = i1 & m1;
  assign n400 = ~n361 & n399;
  assign n401 = n358 & n400;
  assign n402 = ~s1 & n400;
  assign n403 = i1 & q2;
  assign n404 = ~n361 & n403;
  assign n405 = i1 & p2;
  assign n406 = ~n361 & n405;
  assign n407 = i1 & ~l2;
  assign n408 = ~n361 & n407;
  assign n409 = ~q & i1;
  assign n410 = ~n361 & n409;
  assign n411 = ~n408 & ~n410;
  assign n412 = ~n406 & n411;
  assign n413 = ~n404 & n412;
  assign n414 = ~n402 & n413;
  assign n415 = ~n401 & n414;
  assign n416 = ~n398 & n415;
  assign n417 = ~n395 & n416;
  assign n418 = ~n392 & n417;
  assign n419 = ~n389 & n418;
  assign n420 = ~n386 & n419;
  assign d7 = n384 | ~n420;
  assign n422 = ~d1 & ~e1;
  assign n423 = l2 & n422;
  assign e5 = n381 | n423;
  assign n425 = ~p2 & q2;
  assign n426 = p2 & ~q2;
  assign e6 = n425 | n426;
  assign n428 = e4 & i1;
  assign i7 = y3 & n428;
  assign n430 = z3 & i7;
  assign n431 = l3 & n430;
  assign n432 = s & n430;
  assign e7 = n431 | n432;
  assign e8 = ~w0 & ~x0;
  assign n435 = x & j1;
  assign n436 = ~y & n435;
  assign n437 = y & e0;
  assign n438 = ~n297 & ~n437;
  assign f4 = n436 | ~n438;
  assign n440 = ~c1 & ~e1;
  assign n441 = l2 & n440;
  assign f5 = n381 | n441;
  assign n443 = m2 & p2;
  assign n444 = ~n310 & ~n443;
  assign f6 = n308 | ~n444;
  assign n446 = ~n309 & ~n443;
  assign f7 = n308 | ~n446;
  assign n448 = k1 & y1;
  assign n449 = p0 & ~y1;
  assign g4 = n448 | n449;
  assign n451 = ~e1 & l2;
  assign g5 = n381 | n451;
  assign n453 = r0 & x1;
  assign n454 = ~y1 & n453;
  assign n455 = m2 & n454;
  assign n456 = ~q2 & n455;
  assign n457 = ~p2 & n455;
  assign n458 = ~n456 & ~n457;
  assign n459 = p & ~m2;
  assign n460 = p2 & n459;
  assign n461 = q2 & n460;
  assign n462 = n458 & ~n461;
  assign n463 = v3 & n462;
  assign n464 = ~p0 & ~n462;
  assign g6 = n463 | n464;
  assign n466 = ~x1 & y1;
  assign n467 = m2 & n466;
  assign n468 = q & ~m2;
  assign n469 = p2 & n468;
  assign n470 = q2 & n469;
  assign n471 = ~q2 & n467;
  assign n472 = ~p2 & n467;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~n470 & n473;
  assign n475 = q3 & n474;
  assign n476 = ~k1 & ~n474;
  assign g7 = n475 | n476;
  assign h4 = v2 | d8;
  assign n479 = l2 & n378;
  assign h5 = n381 | n479;
  assign n481 = p0 & ~n462;
  assign n482 = ~q0 & n481;
  assign n483 = w3 & n462;
  assign n484 = q0 & n464;
  assign n485 = ~n483 & ~n484;
  assign h6 = n482 | ~n485;
  assign n487 = k1 & ~n474;
  assign n488 = ~l1 & n487;
  assign n489 = r3 & n474;
  assign n490 = l1 & n476;
  assign n491 = ~n489 & ~n490;
  assign h7 = n488 | ~n491;
  assign n493 = ~w2 & d8;
  assign n494 = ~w2 & ~x2;
  assign h8 = n493 | n494;
  assign n496 = ~g0 & h0;
  assign n497 = u2 & n496;
  assign n498 = ~s0 & n497;
  assign n499 = ~t & u;
  assign n500 = u2 & n499;
  assign n501 = s0 & n500;
  assign n502 = ~d8 & ~n501;
  assign i4 = n498 | ~n502;
  assign n504 = ~d1 & l2;
  assign i5 = n381 | n504;
  assign n506 = ~y0 & e8;
  assign n507 = ~z0 & n506;
  assign n508 = u1 & n507;
  assign n509 = w0 & ~x0;
  assign n510 = y0 & n509;
  assign n511 = ~z0 & n510;
  assign n512 = u1 & n511;
  assign n513 = ~w0 & x0;
  assign n514 = ~y0 & n513;
  assign n515 = z0 & n514;
  assign n516 = u1 & n515;
  assign n517 = w0 & x0;
  assign n518 = y0 & n517;
  assign n519 = z0 & n518;
  assign n520 = u1 & n519;
  assign n521 = ~n516 & ~n520;
  assign n522 = ~n512 & n521;
  assign n523 = ~n508 & n522;
  assign n524 = ~z0 & n514;
  assign n525 = y0 & e8;
  assign n526 = ~z0 & n525;
  assign n527 = z0 & w0;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~n524 & n528;
  assign n530 = j2 & ~n523;
  assign n531 = j2 & ~n529;
  assign n532 = ~n530 & ~n531;
  assign n533 = k0 & l0;
  assign n534 = m0 & n533;
  assign n535 = n532 & n534;
  assign n536 = ~n3 & ~o3;
  assign n537 = ~t3 & n536;
  assign n538 = a2 & ~n537;
  assign n539 = j0 & n535;
  assign n540 = n535 & n538;
  assign n541 = ~n245 & n540;
  assign n542 = ~n539 & ~n541;
  assign i6 = l3 & ~n542;
  assign n544 = h0 & u2;
  assign n545 = ~s0 & n544;
  assign n546 = c2 & d8;
  assign n547 = u & u2;
  assign n548 = s0 & n547;
  assign n549 = ~n546 & ~n548;
  assign j4 = n545 | ~n549;
  assign n551 = ~c1 & l2;
  assign j5 = n381 | n551;
  assign n553 = r1 & ~n358;
  assign n554 = t0 & n496;
  assign n555 = ~l3 & n554;
  assign n556 = ~q2 & r0;
  assign n557 = ~n553 & n556;
  assign n558 = ~p2 & r0;
  assign n559 = ~n553 & n558;
  assign n560 = ~l2 & r0;
  assign n561 = ~n553 & n560;
  assign n562 = ~n555 & ~n561;
  assign n563 = ~n559 & n562;
  assign j6 = n557 | ~n563;
  assign j7 = ~m1 & ~d8;
  assign k6 = ~k2 & ~m0;
  assign k7 = i1 | n467;
  assign n568 = n & c1;
  assign n569 = d1 & n568;
  assign l5 = e1 & n569;
  assign n571 = ~k2 & m2;
  assign n572 = ~i3 & n571;
  assign n573 = h3 & n571;
  assign n574 = ~k2 & p2;
  assign n575 = ~k6 & ~n574;
  assign n576 = ~n573 & n575;
  assign l6 = n572 | ~n576;
  assign n578 = ~n358 & ~j4;
  assign n579 = a & f0;
  assign n580 = ~n578 & ~n579;
  assign n581 = r2 & n580;
  assign n582 = b2 & v1;
  assign n583 = ~d8 & n582;
  assign n584 = f3 & ~n583;
  assign n585 = ~h3 & i3;
  assign n586 = m3 & n585;
  assign n587 = ~n583 & n586;
  assign n588 = ~n584 & ~n587;
  assign n589 = h3 & ~i3;
  assign n590 = m3 & n589;
  assign n591 = ~n583 & n590;
  assign n592 = e3 & ~n583;
  assign n593 = ~n591 & ~n592;
  assign n594 = n588 & n593;
  assign n595 = g3 & ~n583;
  assign n596 = ~n553 & n595;
  assign n597 = ~n594 & n596;
  assign n598 = n1 & d8;
  assign n599 = ~b2 & n1;
  assign n600 = n1 & ~s1;
  assign n601 = n1 & r1;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n599 & n602;
  assign n604 = ~n598 & n603;
  assign n605 = s0 & d8;
  assign n606 = ~b2 & s0;
  assign n607 = s0 & s1;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n605 & n608;
  assign n610 = y2 & ~d8;
  assign n611 = ~n553 & n610;
  assign n612 = ~n594 & n611;
  assign n613 = n597 & n612;
  assign n614 = ~z3 & n613;
  assign n615 = u2 & ~d8;
  assign n616 = ~z3 & n615;
  assign n617 = ~s & n616;
  assign n618 = ~l3 & n617;
  assign n619 = v2 & ~n604;
  assign n620 = ~d8 & n619;
  assign n621 = ~z3 & n620;
  assign n622 = u2 & ~n609;
  assign n623 = ~d8 & n622;
  assign n624 = ~z3 & n623;
  assign n625 = v2 & ~y3;
  assign n626 = ~d8 & n625;
  assign n627 = ~z3 & n626;
  assign n628 = w2 & n284;
  assign n629 = n282 & n628;
  assign n630 = ~n286 & ~n629;
  assign n631 = ~n627 & n630;
  assign n632 = ~n624 & n631;
  assign n633 = ~n621 & n632;
  assign n634 = ~n618 & n633;
  assign n635 = ~n614 & n634;
  assign n636 = ~n581 & ~n635;
  assign n637 = u2 & n636;
  assign n638 = s & ~l3;
  assign n639 = ~n597 & ~n638;
  assign l7 = n637 | ~n639;
  assign n641 = ~f & ~r1;
  assign n642 = s1 & n641;
  assign n643 = ~e & ~r1;
  assign n644 = s1 & n643;
  assign n645 = ~d & ~r1;
  assign n646 = s1 & n645;
  assign n647 = ~f & b1;
  assign n648 = ~d & b1;
  assign n649 = ~e & b1;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n647 & n650;
  assign n652 = ~n646 & n651;
  assign n653 = ~n644 & n652;
  assign m5 = n642 | ~n653;
  assign n655 = ~z2 & ~a3;
  assign n656 = b3 & ~c3;
  assign n657 = ~n553 & n656;
  assign n658 = n655 & n657;
  assign n659 = o0 & n658;
  assign n660 = l2 & n659;
  assign n661 = ~a3 & b3;
  assign n662 = ~c3 & n661;
  assign n663 = n655 & n662;
  assign n664 = o0 & n663;
  assign n665 = l2 & n664;
  assign n666 = z2 & b3;
  assign n667 = ~c3 & n666;
  assign n668 = n655 & n667;
  assign n669 = o0 & n668;
  assign n670 = l2 & n669;
  assign n671 = d3 & ~n553;
  assign n672 = n655 & n671;
  assign n673 = o0 & n672;
  assign n674 = l2 & n673;
  assign n675 = ~a3 & d3;
  assign n676 = n655 & n675;
  assign n677 = o0 & n676;
  assign n678 = l2 & n677;
  assign n679 = z2 & d3;
  assign n680 = n655 & n679;
  assign n681 = o0 & n680;
  assign n682 = l2 & n681;
  assign n683 = ~b3 & ~c3;
  assign n684 = ~d3 & n683;
  assign n685 = ~n553 & n684;
  assign n686 = n655 & n685;
  assign n687 = ~a3 & ~b3;
  assign n688 = ~c3 & n687;
  assign n689 = ~d3 & n688;
  assign n690 = n655 & n689;
  assign n691 = z2 & ~b3;
  assign n692 = ~c3 & n691;
  assign n693 = ~d3 & n692;
  assign n694 = n655 & n693;
  assign n695 = ~n690 & ~n694;
  assign n696 = ~n686 & n695;
  assign n697 = ~n682 & n696;
  assign n698 = ~n678 & n697;
  assign n699 = ~n674 & n698;
  assign n700 = ~n670 & n699;
  assign n701 = ~n665 & n700;
  assign n702 = ~n660 & n701;
  assign n703 = m3 & ~n553;
  assign n704 = n702 & n703;
  assign n705 = n655 & n704;
  assign n706 = h3 & i3;
  assign n707 = n702 & n706;
  assign n708 = n655 & n707;
  assign n709 = ~n705 & ~n708;
  assign n710 = n244 & n702;
  assign n711 = n655 & n710;
  assign n712 = h3 & ~n709;
  assign n713 = ~n555 & ~n711;
  assign m6 = n712 | ~n713;
  assign n715 = ~n537 & n604;
  assign m7 = ~n597 & n715;
  assign n717 = e1 & n316;
  assign n718 = n467 & n717;
  assign n719 = ~w1 & n284;
  assign n720 = ~n & n467;
  assign n721 = n458 & ~n720;
  assign n722 = ~n719 & n721;
  assign n4 = n718 | ~n722;
  assign n724 = ~f2 & g2;
  assign n725 = h2 & n724;
  assign n726 = ~l2 & n725;
  assign n5 = a | n726;
  assign n728 = n589 & n709;
  assign n729 = i3 & ~n709;
  assign n730 = ~n711 & ~n729;
  assign n6 = n728 | ~n730;
  assign n7 = n597 & n604;
  assign o4 = w1 & n284;
  assign n734 = ~g2 & h2;
  assign n735 = ~l2 & n734;
  assign n736 = h2 & ~l2;
  assign n737 = f2 & n736;
  assign o5 = n735 | n737;
  assign n739 = ~n585 & ~n589;
  assign n740 = n703 & ~n739;
  assign n741 = ~n655 & n740;
  assign n742 = ~n702 & n740;
  assign n743 = ~n655 & n706;
  assign n744 = ~n702 & n706;
  assign n745 = ~n655 & n711;
  assign n746 = ~n702 & n711;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n744 & n747;
  assign n749 = ~n743 & n748;
  assign n750 = ~n742 & n749;
  assign n751 = ~n741 & n750;
  assign n752 = z2 & n739;
  assign n753 = n702 & n752;
  assign n754 = z2 & n751;
  assign n755 = n702 & n754;
  assign n756 = ~h0 & ~n751;
  assign n757 = ~s0 & n756;
  assign n758 = z2 & ~n751;
  assign n759 = n739 & n758;
  assign n760 = ~u & ~n751;
  assign n761 = s0 & n760;
  assign n762 = ~n759 & ~n761;
  assign n763 = ~n757 & n762;
  assign n764 = ~n755 & n763;
  assign o6 = n753 | ~n764;
  assign n766 = n537 & ~n597;
  assign o7 = ~n604 | n766;
  assign n768 = ~a & ~t2;
  assign n769 = n581 & n768;
  assign n770 = ~g2 & n769;
  assign n771 = ~h2 & n770;
  assign n772 = l2 & n771;
  assign n773 = ~a & t1;
  assign n774 = n581 & n773;
  assign n775 = ~g2 & n774;
  assign n776 = ~h2 & n775;
  assign n777 = l2 & n776;
  assign n778 = ~n635 & n768;
  assign n779 = ~g2 & n778;
  assign n780 = ~h2 & n779;
  assign n781 = l2 & n780;
  assign n782 = ~n635 & n773;
  assign n783 = ~g2 & n782;
  assign n784 = ~h2 & n783;
  assign n785 = l2 & n784;
  assign n786 = ~f2 & n769;
  assign n787 = ~g2 & n786;
  assign n788 = l2 & n787;
  assign n789 = ~f2 & n774;
  assign n790 = ~g2 & n789;
  assign n791 = l2 & n790;
  assign n792 = ~f2 & n778;
  assign n793 = ~g2 & n792;
  assign n794 = l2 & n793;
  assign n795 = ~f2 & n782;
  assign n796 = ~g2 & n795;
  assign n797 = l2 & n796;
  assign n798 = z1 & n769;
  assign n799 = ~l2 & n798;
  assign n800 = z1 & n774;
  assign n801 = ~l2 & n800;
  assign n802 = z1 & n778;
  assign n803 = ~l2 & n802;
  assign n804 = z1 & n782;
  assign n805 = ~l2 & n804;
  assign n806 = ~h2 & n786;
  assign n807 = ~h2 & n789;
  assign n808 = ~h2 & n792;
  assign n809 = ~h2 & n795;
  assign n810 = ~h2 & n798;
  assign n811 = ~h2 & n800;
  assign n812 = ~h2 & n802;
  assign n813 = ~h2 & n804;
  assign n814 = ~g2 & n798;
  assign n815 = ~g2 & n800;
  assign n816 = ~g2 & n802;
  assign n817 = ~g2 & n804;
  assign n818 = ~f2 & n798;
  assign n819 = ~f2 & n800;
  assign n820 = ~f2 & n802;
  assign n821 = ~f2 & n804;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~n819 & n822;
  assign n824 = ~n818 & n823;
  assign n825 = ~n817 & n824;
  assign n826 = ~n816 & n825;
  assign n827 = ~n815 & n826;
  assign n828 = ~n814 & n827;
  assign n829 = ~n813 & n828;
  assign n830 = ~n812 & n829;
  assign n831 = ~n811 & n830;
  assign n832 = ~n810 & n831;
  assign n833 = ~n809 & n832;
  assign n834 = ~n808 & n833;
  assign n835 = ~n807 & n834;
  assign n836 = ~n806 & n835;
  assign n837 = ~n805 & n836;
  assign n838 = ~n803 & n837;
  assign n839 = ~n801 & n838;
  assign n840 = ~n799 & n839;
  assign n841 = ~n797 & n840;
  assign n842 = ~n794 & n841;
  assign n843 = ~n791 & n842;
  assign n844 = ~n788 & n843;
  assign n845 = ~n785 & n844;
  assign n846 = ~n781 & n845;
  assign n847 = ~n777 & n846;
  assign p4 = n772 | ~n847;
  assign n849 = g2 & l2;
  assign n850 = g2 & ~h2;
  assign n851 = f2 & l2;
  assign n852 = ~h2 & ~l2;
  assign n853 = f2 & ~h2;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~n851 & n854;
  assign n856 = ~n850 & n855;
  assign p5 = n849 | ~n856;
  assign n858 = a3 & h0;
  assign n859 = ~n553 & n858;
  assign n860 = ~s0 & n859;
  assign n861 = n702 & n860;
  assign n862 = z2 & h0;
  assign n863 = a3 & n862;
  assign n864 = ~s0 & n863;
  assign n865 = n702 & n864;
  assign n866 = u & a3;
  assign n867 = ~n553 & n866;
  assign n868 = s0 & n867;
  assign n869 = n702 & n868;
  assign n870 = z2 & u;
  assign n871 = a3 & n870;
  assign n872 = s0 & n871;
  assign n873 = n702 & n872;
  assign n874 = ~n751 & n858;
  assign n875 = ~n553 & n874;
  assign n876 = ~s0 & n875;
  assign n877 = ~n751 & n863;
  assign n878 = ~s0 & n877;
  assign n879 = ~n751 & n866;
  assign n880 = ~n553 & n879;
  assign n881 = s0 & n880;
  assign n882 = ~n751 & n871;
  assign n883 = s0 & n882;
  assign n884 = a3 & n751;
  assign n885 = ~n553 & n884;
  assign n886 = n702 & n885;
  assign n887 = z2 & a3;
  assign n888 = n751 & n887;
  assign n889 = n702 & n888;
  assign n890 = ~h0 & i0;
  assign n891 = ~n751 & n890;
  assign n892 = ~s0 & n891;
  assign n893 = ~n739 & ~n751;
  assign n894 = ~u & v;
  assign n895 = ~n751 & n894;
  assign n896 = s0 & n895;
  assign n897 = ~n893 & ~n896;
  assign n898 = ~n892 & n897;
  assign n899 = ~n889 & n898;
  assign n900 = ~n886 & n899;
  assign n901 = ~n883 & n900;
  assign n902 = ~n881 & n901;
  assign n903 = ~n878 & n902;
  assign n904 = ~n876 & n903;
  assign n905 = ~n873 & n904;
  assign n906 = ~n869 & n905;
  assign n907 = ~n865 & n906;
  assign p6 = n861 | ~n907;
  assign n909 = n428 & n604;
  assign n910 = ~d8 & n909;
  assign n911 = ~n597 & n910;
  assign n912 = y3 & n911;
  assign n913 = n609 & n912;
  assign n914 = a4 & n913;
  assign n915 = l3 & n914;
  assign n916 = ~n542 & n604;
  assign n917 = ~d8 & n916;
  assign n918 = ~n597 & n917;
  assign n919 = y3 & n918;
  assign n920 = n609 & n919;
  assign n921 = a4 & n920;
  assign n922 = l3 & n921;
  assign n923 = s & n914;
  assign n924 = s & n921;
  assign n925 = ~d8 & n428;
  assign n926 = ~n597 & n925;
  assign n927 = ~v2 & n926;
  assign n928 = n609 & n927;
  assign n929 = a4 & n928;
  assign n930 = l3 & n929;
  assign n931 = ~d8 & ~n542;
  assign n932 = ~n597 & n931;
  assign n933 = ~v2 & n932;
  assign n934 = n609 & n933;
  assign n935 = a4 & n934;
  assign n936 = l3 & n935;
  assign n937 = s & n929;
  assign n938 = s & n935;
  assign n939 = ~u2 & n911;
  assign n940 = y3 & n939;
  assign n941 = a4 & n940;
  assign n942 = ~u2 & n918;
  assign n943 = y3 & n942;
  assign n944 = a4 & n943;
  assign n945 = ~d8 & n604;
  assign n946 = n597 & n945;
  assign n947 = y3 & n946;
  assign n948 = n594 & n947;
  assign n949 = a4 & n948;
  assign n950 = n553 & n947;
  assign n951 = a4 & n950;
  assign n952 = ~y2 & n946;
  assign n953 = y3 & n952;
  assign n954 = a4 & n953;
  assign n955 = ~u2 & n926;
  assign n956 = ~v2 & n955;
  assign n957 = a4 & n956;
  assign n958 = ~u2 & n932;
  assign n959 = ~v2 & n958;
  assign n960 = a4 & n959;
  assign n961 = ~d8 & n597;
  assign n962 = ~v2 & n961;
  assign n963 = n594 & n962;
  assign n964 = a4 & n963;
  assign n965 = n553 & n962;
  assign n966 = a4 & n965;
  assign n967 = ~y2 & n962;
  assign n968 = a4 & n967;
  assign n969 = ~n581 & n961;
  assign n970 = a4 & n969;
  assign n971 = ~d8 & ~n604;
  assign n972 = ~n581 & n971;
  assign n973 = a4 & n972;
  assign n974 = ~n581 & n925;
  assign n975 = a4 & n974;
  assign n976 = ~n581 & n931;
  assign n977 = a4 & n976;
  assign n978 = ~v2 & n971;
  assign n979 = a4 & n978;
  assign n980 = ~n977 & ~n979;
  assign n981 = ~n975 & n980;
  assign n982 = ~n973 & n981;
  assign n983 = ~n970 & n982;
  assign n984 = ~n968 & n983;
  assign n985 = ~n966 & n984;
  assign n986 = ~n964 & n985;
  assign n987 = ~n960 & n986;
  assign n988 = ~n957 & n987;
  assign n989 = ~n954 & n988;
  assign n990 = ~n951 & n989;
  assign n991 = ~n949 & n990;
  assign n992 = ~n944 & n991;
  assign n993 = ~n941 & n992;
  assign n994 = ~n938 & n993;
  assign n995 = ~n937 & n994;
  assign n996 = ~n936 & n995;
  assign n997 = ~n930 & n996;
  assign n998 = ~n924 & n997;
  assign n999 = ~n923 & n998;
  assign n1000 = ~n922 & n999;
  assign p7 = n915 | ~n1000;
  assign n1002 = ~a & t2;
  assign n1003 = ~t1 & n1002;
  assign n1004 = ~f2 & n1003;
  assign n1005 = ~h2 & n1004;
  assign n1006 = a1 & t2;
  assign q4 = n1005 | n1006;
  assign n1008 = g0 & t0;
  assign n1009 = ~l2 & n1008;
  assign n1010 = ~n523 & n1009;
  assign n1011 = o & ~p;
  assign n1012 = ~q & n1011;
  assign n1013 = ~h0 & ~l3;
  assign n1014 = n538 & n1013;
  assign n1015 = t0 & n1014;
  assign n1016 = n655 & n1015;
  assign n1017 = ~l3 & n538;
  assign n1018 = t0 & n1017;
  assign n1019 = n581 & n1018;
  assign n1020 = ~u2 & n1018;
  assign n1021 = z3 & ~h0;
  assign n1022 = ~s0 & n1021;
  assign n1023 = ~h0 & d8;
  assign n1024 = ~s0 & n1023;
  assign n1025 = z3 & ~u;
  assign n1026 = s0 & n1025;
  assign n1027 = ~u & d8;
  assign n1028 = s0 & n1027;
  assign n1029 = n538 & n1010;
  assign n1030 = n709 & ~n739;
  assign n1031 = n529 & ~n532;
  assign n1032 = ~n532 & ~n1012;
  assign n1033 = ~l2 & ~n532;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1031 & n1034;
  assign n1036 = ~n1030 & n1035;
  assign n1037 = ~n1029 & n1036;
  assign n1038 = ~n1028 & n1037;
  assign n1039 = ~n1026 & n1038;
  assign n1040 = ~n1024 & n1039;
  assign n1041 = ~n1022 & n1040;
  assign n1042 = ~n1020 & n1041;
  assign n1043 = ~n1019 & n1042;
  assign n1044 = ~n1016 & n1043;
  assign n1045 = n245 & n538;
  assign n1046 = j0 & n245;
  assign n1047 = ~n535 & n538;
  assign n1048 = j0 & ~n535;
  assign n1049 = n538 & ~n1044;
  assign n1050 = j0 & ~n1044;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = ~n1048 & n1051;
  assign n1053 = ~n1047 & n1052;
  assign n1054 = ~n1046 & n1053;
  assign q5 = n1045 | ~n1054;
  assign n1056 = c3 & o0;
  assign n1057 = b3 & o0;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = b3 & n1058;
  assign n1060 = n702 & n1059;
  assign n1061 = z2 & ~n702;
  assign q6 = n1060 | n1061;
  assign n1063 = d4 & ~s1;
  assign n1064 = ~s1 & n303;
  assign n1065 = ~s1 & d8;
  assign n1066 = ~n1064 & ~n1065;
  assign q7 = n1063 | ~n1066;
  assign n1068 = h2 & n329;
  assign n1069 = ~q1 & n1068;
  assign n1070 = ~r1 & n1069;
  assign n1071 = ~s1 & n1070;
  assign n1072 = ~g2 & n1071;
  assign n1073 = ~o & n1072;
  assign n1074 = ~p & n1073;
  assign n1075 = ~q & n1074;
  assign n1076 = a & h2;
  assign n1077 = ~q1 & n1076;
  assign n1078 = ~r1 & n1077;
  assign n1079 = ~s1 & n1078;
  assign n1080 = ~g2 & n1079;
  assign n1081 = ~o & n1080;
  assign n1082 = ~p & n1081;
  assign n1083 = ~q & n1082;
  assign n1084 = ~f1 & n1068;
  assign n1085 = ~g1 & n1084;
  assign n1086 = ~h1 & n1085;
  assign n1087 = g2 & n1086;
  assign n1088 = ~o & n1087;
  assign n1089 = ~p & n1088;
  assign n1090 = ~q & n1089;
  assign n1091 = ~f1 & n1076;
  assign n1092 = ~g1 & n1091;
  assign n1093 = ~h1 & n1092;
  assign n1094 = g2 & n1093;
  assign n1095 = ~o & n1094;
  assign n1096 = ~p & n1095;
  assign n1097 = ~q & n1096;
  assign n1098 = a & ~h2;
  assign n1099 = ~f1 & n1098;
  assign n1100 = ~g1 & n1099;
  assign n1101 = ~h1 & n1100;
  assign n1102 = ~q1 & n1101;
  assign n1103 = ~r1 & n1102;
  assign n1104 = ~s1 & n1103;
  assign n1105 = g2 & n1104;
  assign n1106 = ~q1 & n1098;
  assign n1107 = ~r1 & n1106;
  assign n1108 = ~s1 & n1107;
  assign n1109 = ~g2 & n1108;
  assign n1110 = o0 & n329;
  assign n1111 = ~q1 & n1110;
  assign n1112 = ~r1 & n1111;
  assign n1113 = ~s1 & n1112;
  assign n1114 = ~g2 & n1113;
  assign n1115 = a & o0;
  assign n1116 = ~q1 & n1115;
  assign n1117 = ~r1 & n1116;
  assign n1118 = ~s1 & n1117;
  assign n1119 = ~g2 & n1118;
  assign n1120 = ~f1 & n1110;
  assign n1121 = ~g1 & n1120;
  assign n1122 = ~h1 & n1121;
  assign n1123 = g2 & n1122;
  assign n1124 = ~f1 & n1115;
  assign n1125 = ~g1 & n1124;
  assign n1126 = ~h1 & n1125;
  assign n1127 = g2 & n1126;
  assign n1128 = a & ~l2;
  assign n1129 = ~h2 & n1128;
  assign n1130 = ~q1 & n1129;
  assign n1131 = ~r1 & n1130;
  assign n1132 = ~s1 & n1131;
  assign n1133 = ~o & n736;
  assign n1134 = ~p & n1133;
  assign n1135 = ~q & n1134;
  assign n1136 = ~l2 & o0;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~n1132 & n1137;
  assign n1139 = ~n1127 & n1138;
  assign n1140 = ~n1123 & n1139;
  assign n1141 = ~n1119 & n1140;
  assign n1142 = ~n1114 & n1141;
  assign n1143 = ~n1109 & n1142;
  assign n1144 = ~n1105 & n1143;
  assign n1145 = ~n1097 & n1144;
  assign n1146 = ~n1090 & n1145;
  assign n1147 = ~n1083 & n1146;
  assign r4 = n1075 | ~n1147;
  assign n1149 = ~n555 & n1044;
  assign r5 = ~n542 & n1149;
  assign n1151 = c3 & n1058;
  assign n1152 = n702 & n1151;
  assign n1153 = ~n553 & n1152;
  assign n1154 = b3 & c3;
  assign n1155 = n1058 & n1154;
  assign n1156 = n702 & n1155;
  assign n1157 = a3 & ~n702;
  assign n1158 = ~n1156 & ~n1157;
  assign r6 = n1153 | ~n1158;
  assign n1160 = ~r1 & s1;
  assign n1161 = d4 & n1160;
  assign n1162 = n303 & n1160;
  assign n1163 = d8 & n1160;
  assign n1164 = ~n1162 & ~n1163;
  assign r7 = n1161 | ~n1164;
  assign n1166 = ~a & f0;
  assign n1167 = ~a & j4;
  assign n1168 = ~n358 & n1167;
  assign s4 = n1166 | n1168;
  assign n1170 = j2 & n529;
  assign n1171 = n523 & n1170;
  assign n1172 = ~o3 & n538;
  assign s5 = n1171 | n1172;
  assign n1174 = d3 & n702;
  assign n1175 = ~o0 & n1174;
  assign n1176 = c3 & ~n1058;
  assign s6 = n1175 | n1176;
  assign n1178 = a & d;
  assign n1179 = e & n1178;
  assign n1180 = f & n1179;
  assign n1181 = a & ~n;
  assign n1182 = a & ~s1;
  assign n1183 = a & r1;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1181 & n1184;
  assign n1186 = ~n1180 & n1185;
  assign n1187 = o2 & ~n1186;
  assign n1188 = n2 & ~n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = i0 & n636;
  assign n1191 = ~i4 & n1190;
  assign n1192 = ~s0 & n1191;
  assign n1193 = v & n636;
  assign n1194 = ~i4 & n1193;
  assign n1195 = s0 & n1194;
  assign n1196 = n2 & ~n636;
  assign n1197 = n1189 & n1196;
  assign n1198 = ~n2 & ~n636;
  assign n1199 = ~n1189 & n1198;
  assign n1200 = y2 & n636;
  assign n1201 = ~n594 & n1200;
  assign n1202 = i4 & n636;
  assign n1203 = ~h4 & n1202;
  assign n1204 = ~i4 & n636;
  assign n1205 = h4 & n1204;
  assign n1206 = ~n1203 & ~n1205;
  assign n1207 = ~n1201 & n1206;
  assign n1208 = ~n1199 & n1207;
  assign n1209 = ~n1197 & n1208;
  assign n1210 = ~n1195 & n1209;
  assign t4 = n1192 | ~n1210;
  assign n1212 = k0 & ~n655;
  assign n1213 = h0 & k0;
  assign n1214 = k0 & ~n538;
  assign n1215 = ~l2 & ~n1214;
  assign n1216 = ~n1213 & n1215;
  assign t5 = n1212 | ~n1216;
  assign n1218 = ~k2 & l2;
  assign n1219 = n1012 & n1218;
  assign t6 = n1171 | n1219;
  assign n1221 = ~o2 & n1198;
  assign n1222 = ~n1189 & n1221;
  assign n1223 = ~n593 & n1200;
  assign n1224 = ~n588 & n1223;
  assign n1225 = o2 & ~n636;
  assign n1226 = n1189 & n1225;
  assign n1227 = o2 & n1196;
  assign n1228 = n1206 & ~n1227;
  assign n1229 = ~n1226 & n1228;
  assign n1230 = ~n1224 & n1229;
  assign u4 = n1222 | ~n1230;
  assign n1232 = l0 & u2;
  assign n1233 = ~n581 & n1232;
  assign n1234 = l2 & ~n329;
  assign n1235 = l0 & ~n538;
  assign n1236 = l0 & ~s0;
  assign n1237 = ~z1 & ~n1236;
  assign n1238 = ~n1235 & n1237;
  assign n1239 = ~n1234 & n1238;
  assign u5 = n1233 | ~n1239;
  assign u6 = n523 & n1008;
  assign n1242 = n580 & ~n635;
  assign n1243 = o2 & n1242;
  assign n1244 = o2 & n581;
  assign n1245 = n2 & n1242;
  assign n1246 = n2 & n581;
  assign n1247 = ~n635 & n1186;
  assign n1248 = n580 & n1247;
  assign n1249 = r2 & n1186;
  assign n1250 = n580 & n1249;
  assign n1251 = ~n1248 & ~n1250;
  assign n1252 = ~n1246 & n1251;
  assign n1253 = ~n1245 & n1252;
  assign n1254 = ~n1244 & n1253;
  assign v4 = n1243 | ~n1254;
  assign n1256 = ~o & ~n555;
  assign n1257 = p & n1256;
  assign n1258 = ~q & n1257;
  assign n1259 = l2 & n1258;
  assign n1260 = ~i3 & n1259;
  assign n1261 = h3 & n1259;
  assign n1262 = p & ~n555;
  assign n1263 = ~q & n1262;
  assign n1264 = l2 & n1263;
  assign n1265 = p2 & n1264;
  assign n1266 = ~w1 & ~n555;
  assign n1267 = x1 & n1266;
  assign n1268 = ~y1 & n1267;
  assign n1269 = m2 & n1268;
  assign n1270 = m0 & ~n555;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~n1265 & n1271;
  assign n1273 = ~n1261 & n1272;
  assign v5 = n1260 | ~n1273;
  assign n1275 = b & ~n636;
  assign n1276 = n1186 & n1275;
  assign n1277 = ~b & ~n636;
  assign n1278 = ~n1186 & n1277;
  assign n1279 = d2 & n636;
  assign n1280 = ~n1278 & ~n1279;
  assign w4 = n1276 | ~n1280;
  assign w5 = n3 & ~n542;
  assign n1283 = ~c & n1275;
  assign n1284 = ~n1186 & n1283;
  assign n1285 = c & ~n636;
  assign n1286 = n1186 & n1285;
  assign n1287 = e2 & n636;
  assign n1288 = c & n1277;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~n1286 & n1289;
  assign x4 = n1284 | ~n1290;
  assign n1292 = k2 & ~n1012;
  assign n1293 = k2 & ~l2;
  assign n1294 = ~n1010 & ~n1293;
  assign x5 = n1292 | ~n1294;
  assign n1296 = r & ~p3;
  assign n1297 = s2 & u0;
  assign n1298 = r & k3;
  assign n1299 = ~n1297 & ~n1298;
  assign x7 = n1296 | ~n1299;
  assign n1301 = v0 & ~x3;
  assign y4 = a | n1301;
  assign n1303 = l3 & n1008;
  assign y5 = ~n532 | n1303;
  assign y7 = j3 & p3;
  assign d6 = ~p2;
  assign l4 = ~o3;
  assign a5 = m2;
  assign a7 = y0;
  assign b7 = z0;
  assign f8 = w0;
  assign g8 = x0;
  assign k4 = s3;
  assign k5 = l2;
  assign m4 = t3;
  assign s7 = w;
  assign t7 = z;
  assign u7 = a0;
  assign v6 = z6;
  assign v7 = b0;
  assign w6 = y0;
  assign w7 = c0;
  assign x6 = e8;
  assign y6 = w0;
endmodule


