// Benchmark "term1" written by ABC on Tue May 16 16:07:53 2017

module term1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, c0, d0, e0, f0, g0, h0, i0,
    j0, k0, l0, m0, n0, o0, p0, q0, r0, s0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, c0, d0, e0, f0, g0, h0, i0;
  output j0, k0, l0, m0, n0, o0, p0, q0, r0, s0;
  wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754;
  assign n45 = c & ~i0;
  assign n46 = ~d & ~i0;
  assign n47 = c & ~d;
  assign n48 = ~n46 & ~n47;
  assign n49 = ~n45 & n48;
  assign n50 = c & n49;
  assign n51 = ~d & n49;
  assign n52 = h0 & n49;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~n50 & n53;
  assign n55 = ~c & n54;
  assign n56 = d & n54;
  assign n57 = ~h0 & n54;
  assign n58 = ~n56 & ~n57;
  assign k0 = n55 | ~n58;
  assign n60 = e & h;
  assign n61 = d & h;
  assign n62 = d & e;
  assign n63 = ~n61 & ~n62;
  assign n64 = ~n60 & n63;
  assign n65 = d & n64;
  assign n66 = e & n64;
  assign n67 = h & n64;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~n65 & n68;
  assign n70 = ~d & n69;
  assign n71 = ~h & n69;
  assign n72 = ~e & n69;
  assign n73 = ~n71 & ~n72;
  assign n74 = ~n70 & n73;
  assign n75 = ~d & h;
  assign n76 = ~d & e;
  assign n77 = ~n75 & ~n76;
  assign n78 = ~n60 & n77;
  assign n79 = ~d & n78;
  assign n80 = e & n78;
  assign n81 = h & n78;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~n79 & n82;
  assign n84 = ~h & n83;
  assign n85 = ~e & n83;
  assign n86 = ~n84 & ~n85;
  assign n87 = d & n83;
  assign n88 = n86 & ~n87;
  assign n89 = n74 & n88;
  assign n90 = c & n74;
  assign n91 = ~c & n88;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~n89 & n92;
  assign n94 = i & ~j;
  assign n95 = ~c & g;
  assign n96 = ~e & ~h;
  assign n97 = ~d & f;
  assign n98 = ~n96 & ~n97;
  assign n99 = ~n95 & n98;
  assign n100 = ~e & n99;
  assign n101 = ~h & n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = ~e & ~g;
  assign n104 = ~h & n103;
  assign n105 = c & ~e;
  assign n106 = ~h & n105;
  assign n107 = e & ~g;
  assign n108 = h & n107;
  assign n109 = c & e;
  assign n110 = h & n109;
  assign n111 = ~n108 & ~n110;
  assign n112 = ~n106 & n111;
  assign n113 = ~n104 & n112;
  assign n114 = ~f & ~h;
  assign n115 = e & n114;
  assign n116 = d & ~h;
  assign n117 = e & n116;
  assign n118 = ~n115 & ~n117;
  assign n119 = ~n60 & ~n96;
  assign n120 = n97 & n119;
  assign n121 = n118 & n120;
  assign n122 = d & n97;
  assign n123 = n118 & n122;
  assign n124 = ~f & n97;
  assign n125 = n118 & n124;
  assign n126 = e & n119;
  assign n127 = n118 & n126;
  assign n128 = n62 & n118;
  assign n129 = e & ~f;
  assign n130 = n118 & n129;
  assign n131 = ~h & n119;
  assign n132 = n118 & n131;
  assign n133 = n114 & n118;
  assign n134 = n116 & n118;
  assign n135 = ~n133 & ~n134;
  assign n136 = ~n132 & n135;
  assign n137 = ~n130 & n136;
  assign n138 = ~n128 & n137;
  assign n139 = ~n127 & n138;
  assign n140 = ~n125 & n139;
  assign n141 = ~n123 & n140;
  assign n142 = ~n121 & n141;
  assign n143 = n113 & n142;
  assign n144 = n102 & n143;
  assign n145 = c & n113;
  assign n146 = n102 & n145;
  assign n147 = ~g & n113;
  assign n148 = n102 & n147;
  assign n149 = d & n142;
  assign n150 = n102 & n149;
  assign n151 = c & d;
  assign n152 = n102 & n151;
  assign n153 = d & ~g;
  assign n154 = n102 & n153;
  assign n155 = ~f & n142;
  assign n156 = n102 & n155;
  assign n157 = ~f & ~g;
  assign n158 = n102 & n157;
  assign n159 = c & ~f;
  assign n160 = n102 & n159;
  assign n161 = ~n158 & ~n160;
  assign n162 = ~n156 & n161;
  assign n163 = ~n154 & n162;
  assign n164 = ~n152 & n163;
  assign n165 = ~n150 & n164;
  assign n166 = ~n148 & n165;
  assign n167 = ~n146 & n166;
  assign n168 = ~n144 & n167;
  assign n169 = b & n94;
  assign n170 = ~n93 & n169;
  assign n171 = ~b & n94;
  assign n172 = n168 & n171;
  assign l0 = n170 | n172;
  assign n174 = u & v;
  assign n175 = w & n174;
  assign n176 = p & v;
  assign n177 = w & n176;
  assign n178 = q & u;
  assign n179 = w & n178;
  assign n180 = p & q;
  assign n181 = w & n180;
  assign n182 = r & n174;
  assign n183 = r & n176;
  assign n184 = r & n178;
  assign n185 = r & n180;
  assign n186 = ~n184 & ~n185;
  assign n187 = ~n183 & n186;
  assign n188 = ~n182 & n187;
  assign n189 = ~n181 & n188;
  assign n190 = ~n179 & n189;
  assign n191 = ~n177 & n190;
  assign n192 = ~n175 & n191;
  assign n193 = ~t & ~y;
  assign n194 = ~s & ~x;
  assign n195 = ~n192 & ~n194;
  assign n196 = ~n193 & n195;
  assign n197 = ~n151 & ~n196;
  assign n198 = ~a0 & ~c0;
  assign n199 = z & n198;
  assign n200 = b & n199;
  assign m0 = n197 & n200;
  assign n202 = ~p & ~u;
  assign n203 = ~n193 & ~n202;
  assign n204 = ~n194 & n203;
  assign n205 = q & r;
  assign n206 = n204 & n205;
  assign n207 = q & w;
  assign n208 = n204 & n207;
  assign n209 = r & v;
  assign n210 = n204 & n209;
  assign n211 = v & w;
  assign n212 = n204 & n211;
  assign n213 = ~n210 & ~n212;
  assign n214 = ~n208 & n213;
  assign n215 = ~n206 & n214;
  assign n216 = ~d & n215;
  assign n217 = ~c & n215;
  assign n218 = ~n216 & ~n217;
  assign n219 = ~r & ~w;
  assign n220 = ~q & ~v;
  assign n221 = ~n194 & ~n220;
  assign n222 = ~n219 & n221;
  assign n223 = p & t;
  assign n224 = n222 & n223;
  assign n225 = p & y;
  assign n226 = n222 & n225;
  assign n227 = t & u;
  assign n228 = n222 & n227;
  assign n229 = u & y;
  assign n230 = n222 & n229;
  assign n231 = ~n228 & ~n230;
  assign n232 = ~n226 & n231;
  assign n233 = ~n224 & n232;
  assign n234 = ~n194 & ~n202;
  assign n235 = ~n219 & n234;
  assign n236 = q & t;
  assign n237 = n235 & n236;
  assign n238 = q & y;
  assign n239 = n235 & n238;
  assign n240 = t & v;
  assign n241 = n235 & n240;
  assign n242 = v & y;
  assign n243 = n235 & n242;
  assign n244 = ~n241 & ~n243;
  assign n245 = ~n239 & n244;
  assign n246 = ~n237 & n245;
  assign n247 = ~d & n233;
  assign n248 = ~c & n246;
  assign n249 = ~n247 & ~n248;
  assign n250 = n218 & n249;
  assign n251 = ~d0 & n218;
  assign n252 = c0 & n218;
  assign n253 = d0 & n249;
  assign n254 = ~c0 & n249;
  assign n255 = ~c0 & ~d0;
  assign n256 = c0 & d0;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~n254 & n257;
  assign n259 = ~n253 & n258;
  assign n260 = ~n252 & n259;
  assign n261 = ~n251 & n260;
  assign n262 = ~n250 & n261;
  assign n263 = z & ~a0;
  assign n264 = b & n263;
  assign n0 = n262 & n264;
  assign n266 = w & x;
  assign n267 = v & n266;
  assign n268 = s & w;
  assign n269 = v & n268;
  assign n270 = r & x;
  assign n271 = v & n270;
  assign n272 = r & s;
  assign n273 = v & n272;
  assign n274 = q & n266;
  assign n275 = q & n268;
  assign n276 = q & n270;
  assign n277 = q & n272;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~n275 & n278;
  assign n280 = ~n274 & n279;
  assign n281 = ~n273 & n280;
  assign n282 = ~n271 & n281;
  assign n283 = ~n269 & n282;
  assign n284 = ~n267 & n283;
  assign n285 = ~n193 & ~n284;
  assign n286 = ~n202 & n285;
  assign n287 = x & n174;
  assign n288 = x & n176;
  assign n289 = x & n178;
  assign n290 = x & n180;
  assign n291 = s & n174;
  assign n292 = s & n176;
  assign n293 = s & n178;
  assign n294 = s & n180;
  assign n295 = ~n293 & ~n294;
  assign n296 = ~n292 & n295;
  assign n297 = ~n291 & n296;
  assign n298 = ~n290 & n297;
  assign n299 = ~n289 & n298;
  assign n300 = ~n288 & n299;
  assign n301 = ~n287 & n300;
  assign n302 = ~n219 & ~n301;
  assign n303 = ~n193 & n302;
  assign n304 = n286 & n303;
  assign n305 = c0 & n286;
  assign n306 = d0 & n303;
  assign n307 = ~n256 & ~n306;
  assign n308 = ~n305 & n307;
  assign n309 = ~n304 & n308;
  assign n310 = ~d & e0;
  assign n311 = n309 & n310;
  assign n312 = ~n202 & ~n220;
  assign n313 = ~n194 & n312;
  assign n314 = r & t;
  assign n315 = n313 & n314;
  assign n316 = t & w;
  assign n317 = n313 & n316;
  assign n318 = r & y;
  assign n319 = n313 & n318;
  assign n320 = w & y;
  assign n321 = n313 & n320;
  assign n322 = ~n319 & ~n321;
  assign n323 = ~n317 & n322;
  assign n324 = ~n315 & n323;
  assign n325 = ~d0 & n246;
  assign n326 = ~c0 & n324;
  assign n327 = ~n325 & ~n326;
  assign n328 = d0 & ~e0;
  assign n329 = n218 & n327;
  assign n330 = ~n311 & n329;
  assign n331 = n327 & ~n328;
  assign n332 = ~n311 & n331;
  assign n333 = ~c0 & n327;
  assign n334 = ~n311 & n333;
  assign n335 = c & n218;
  assign n336 = ~n311 & n335;
  assign n337 = c & ~n328;
  assign n338 = ~n311 & n337;
  assign n339 = c & ~c0;
  assign n340 = ~n311 & n339;
  assign n341 = ~e0 & n218;
  assign n342 = ~n311 & n341;
  assign n343 = ~e0 & ~n328;
  assign n344 = ~n311 & n343;
  assign n345 = ~c0 & ~e0;
  assign n346 = ~n311 & n345;
  assign n347 = ~n344 & ~n346;
  assign n348 = ~n342 & n347;
  assign n349 = ~n340 & n348;
  assign n350 = ~n338 & n349;
  assign n351 = ~n336 & n350;
  assign n352 = ~n334 & n351;
  assign n353 = ~n332 & n352;
  assign n354 = ~n330 & n353;
  assign o0 = n264 & n354;
  assign n356 = x & n316;
  assign n357 = x & n320;
  assign n358 = e0 & n256;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n356 & n359;
  assign n361 = x & y;
  assign n362 = t & x;
  assign n363 = s & y;
  assign n364 = s & t;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n362 & n365;
  assign n367 = ~n361 & n366;
  assign n368 = n193 & n367;
  assign n369 = n360 & n368;
  assign n370 = ~s & n367;
  assign n371 = n360 & n370;
  assign n372 = ~w & n367;
  assign n373 = n360 & n372;
  assign n374 = ~r & n193;
  assign n375 = n360 & n374;
  assign n376 = ~r & ~s;
  assign n377 = n360 & n376;
  assign n378 = n219 & n360;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n375 & n379;
  assign n381 = ~n373 & n380;
  assign n382 = ~n371 & n381;
  assign n383 = ~n369 & n382;
  assign n384 = d0 & e0;
  assign n385 = c0 & n384;
  assign n386 = n174 & n383;
  assign n387 = n176 & n383;
  assign n388 = n178 & n383;
  assign n389 = n180 & n383;
  assign n390 = n383 & n385;
  assign n391 = ~n389 & ~n390;
  assign n392 = ~n388 & n391;
  assign n393 = ~n387 & n392;
  assign n394 = ~n386 & n393;
  assign n395 = ~d & f0;
  assign n396 = n394 & n395;
  assign n397 = ~n193 & ~n194;
  assign n398 = ~e0 & n193;
  assign n399 = ~d0 & n193;
  assign n400 = ~c0 & n193;
  assign n401 = ~x & ~e0;
  assign n402 = ~w & ~e0;
  assign n403 = ~x & ~d0;
  assign n404 = ~w & ~d0;
  assign n405 = ~x & ~c0;
  assign n406 = ~w & ~c0;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n404 & n407;
  assign n409 = ~n403 & n408;
  assign n410 = ~n402 & n409;
  assign n411 = ~n401 & n410;
  assign n412 = ~n400 & n411;
  assign n413 = ~n399 & n412;
  assign n414 = ~n398 & n413;
  assign n415 = ~n193 & n268;
  assign n416 = r & n397;
  assign n417 = ~n414 & ~n416;
  assign n418 = ~n415 & n417;
  assign n419 = n220 & ~n385;
  assign n420 = n202 & ~n385;
  assign n421 = ~n418 & ~n420;
  assign n422 = ~n419 & n421;
  assign n423 = e0 & ~f0;
  assign n424 = d0 & n423;
  assign n425 = n218 & n422;
  assign n426 = ~n396 & n425;
  assign n427 = n422 & ~n424;
  assign n428 = ~n396 & n427;
  assign n429 = ~c0 & n422;
  assign n430 = ~n396 & n429;
  assign n431 = n335 & ~n396;
  assign n432 = c & ~n424;
  assign n433 = ~n396 & n432;
  assign n434 = n339 & ~n396;
  assign n435 = ~f0 & n218;
  assign n436 = ~n396 & n435;
  assign n437 = ~f0 & ~n424;
  assign n438 = ~n396 & n437;
  assign n439 = ~c0 & ~f0;
  assign n440 = ~n396 & n439;
  assign n441 = ~n438 & ~n440;
  assign n442 = ~n436 & n441;
  assign n443 = ~n434 & n442;
  assign n444 = ~n433 & n443;
  assign n445 = ~n431 & n444;
  assign n446 = ~n430 & n445;
  assign n447 = ~n428 & n446;
  assign n448 = ~n426 & n447;
  assign p0 = n264 & n448;
  assign n450 = ~n219 & n397;
  assign n451 = ~n194 & n211;
  assign n452 = y & n451;
  assign n453 = t & n451;
  assign n454 = ~n452 & ~n453;
  assign n455 = w & n361;
  assign n456 = w & n362;
  assign n457 = w & n363;
  assign n458 = w & n364;
  assign n459 = r & n361;
  assign n460 = r & n362;
  assign n461 = r & n363;
  assign n462 = r & n364;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n460 & n463;
  assign n465 = ~n459 & n464;
  assign n466 = ~n458 & n465;
  assign n467 = ~n457 & n466;
  assign n468 = ~n456 & n467;
  assign n469 = ~n455 & n468;
  assign n470 = n367 & n469;
  assign n471 = n454 & n470;
  assign n472 = ~r & n469;
  assign n473 = n454 & n472;
  assign n474 = ~v & n469;
  assign n475 = n454 & n474;
  assign n476 = ~q & n367;
  assign n477 = n454 & n476;
  assign n478 = ~q & ~r;
  assign n479 = n454 & n478;
  assign n480 = n220 & n454;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n477 & n481;
  assign n483 = ~n475 & n482;
  assign n484 = ~n473 & n483;
  assign n485 = ~n471 & n484;
  assign n486 = f0 & ~g0;
  assign n487 = n385 & n486;
  assign n488 = ~c & ~a0;
  assign n489 = ~n487 & n488;
  assign n490 = ~d & ~a0;
  assign n491 = ~n487 & n490;
  assign n492 = ~n489 & ~n491;
  assign n493 = b & z;
  assign n494 = ~n492 & n493;
  assign n495 = e0 & f0;
  assign n496 = n256 & n495;
  assign n497 = n469 & n496;
  assign n498 = n494 & n497;
  assign n499 = ~u & n496;
  assign n500 = n494 & n499;
  assign n501 = ~v & n496;
  assign n502 = n494 & n501;
  assign n503 = ~g0 & n469;
  assign n504 = n494 & n503;
  assign n505 = ~u & ~g0;
  assign n506 = n494 & n505;
  assign n507 = ~v & ~g0;
  assign n508 = n494 & n507;
  assign n509 = ~n506 & ~n508;
  assign n510 = ~n504 & n509;
  assign n511 = ~n502 & n510;
  assign n512 = ~n500 & n511;
  assign n513 = ~n498 & n512;
  assign n514 = n178 & n450;
  assign n515 = p & n485;
  assign n516 = ~n513 & ~n515;
  assign q0 = n514 | ~n516;
  assign n518 = n205 & n364;
  assign n519 = ~m & n364;
  assign n520 = ~l & r;
  assign n521 = n364 & n520;
  assign n522 = ~o & s;
  assign n523 = ~n & t;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n364 & n524;
  assign n526 = ~r & ~n519;
  assign n527 = ~q & ~n521;
  assign n528 = ~n525 & ~n527;
  assign n529 = ~n526 & n528;
  assign n530 = ~k & n205;
  assign n531 = n364 & n530;
  assign n532 = ~r & ~t;
  assign n533 = g0 & ~n531;
  assign n534 = ~n532 & n533;
  assign n535 = n314 & n534;
  assign n536 = s & n534;
  assign n537 = ~n535 & ~n536;
  assign n538 = ~f0 & n255;
  assign n539 = ~e0 & ~f0;
  assign n540 = ~n537 & ~n539;
  assign n541 = ~n538 & n540;
  assign n542 = n255 & n462;
  assign n543 = n541 & n542;
  assign n544 = ~e0 & n462;
  assign n545 = n541 & n544;
  assign n546 = ~f0 & n462;
  assign n547 = n541 & n546;
  assign n548 = q & n255;
  assign n549 = n541 & n548;
  assign n550 = q & ~e0;
  assign n551 = n541 & n550;
  assign n552 = q & ~f0;
  assign n553 = n541 & n552;
  assign n554 = ~n551 & ~n553;
  assign n555 = ~n549 & n554;
  assign n556 = ~n547 & n555;
  assign n557 = ~n545 & n556;
  assign n558 = ~n543 & n557;
  assign n559 = ~p & ~n518;
  assign n560 = p & n529;
  assign n561 = ~n558 & ~n560;
  assign n562 = ~n559 & n561;
  assign n563 = p & ~q;
  assign n564 = l & n563;
  assign n565 = c0 & e0;
  assign n566 = ~f0 & ~n565;
  assign n567 = ~n384 & n566;
  assign n568 = ~n255 & n495;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~p & q;
  assign n571 = k & n570;
  assign n572 = o & p;
  assign n573 = n277 & n572;
  assign n574 = ~d0 & ~f0;
  assign n575 = ~c0 & n574;
  assign n576 = ~t & n573;
  assign n577 = ~n575 & n576;
  assign n578 = f0 & n255;
  assign n579 = n577 & n578;
  assign n580 = e0 & n255;
  assign n581 = n577 & n580;
  assign n582 = n423 & n577;
  assign n583 = ~e0 & f0;
  assign n584 = n577 & n583;
  assign n585 = ~n582 & ~n584;
  assign n586 = ~n581 & n585;
  assign n587 = ~n579 & n586;
  assign n588 = ~s & t;
  assign n589 = r & n588;
  assign n590 = ~r & n364;
  assign n591 = m & n180;
  assign n592 = n & n180;
  assign n593 = ~n538 & ~n539;
  assign n594 = n255 & n593;
  assign n595 = ~f0 & n593;
  assign n596 = ~e0 & n593;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n594 & n597;
  assign n599 = ~n589 & ~n590;
  assign n600 = n587 & n599;
  assign n601 = ~n589 & ~n591;
  assign n602 = n587 & n601;
  assign n603 = ~n590 & ~n592;
  assign n604 = n587 & n603;
  assign n605 = n587 & n598;
  assign n606 = ~n591 & ~n592;
  assign n607 = n587 & n606;
  assign n608 = ~n605 & ~n607;
  assign n609 = ~n604 & n608;
  assign n610 = ~n602 & n609;
  assign n611 = ~n600 & n610;
  assign n612 = n462 & n569;
  assign n613 = n564 & n612;
  assign n614 = n462 & n571;
  assign n615 = n569 & n614;
  assign n616 = ~n611 & ~n615;
  assign n617 = ~n613 & n616;
  assign n618 = n562 & n617;
  assign n619 = h0 & n562;
  assign n620 = ~g0 & n562;
  assign n621 = ~h0 & n617;
  assign n622 = ~g0 & ~h0;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n620 & n623;
  assign n625 = ~n619 & n624;
  assign n626 = ~n618 & n625;
  assign n627 = a & ~a0;
  assign r0 = n626 & n627;
  assign n629 = f0 & n384;
  assign n630 = f0 & n565;
  assign n631 = ~f0 & ~g0;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n629 & n632;
  assign n634 = ~k & q;
  assign n635 = n462 & n634;
  assign n636 = ~n376 & ~n633;
  assign n637 = ~n635 & n636;
  assign n638 = n272 & n637;
  assign n639 = t & n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = e0 & ~g0;
  assign n642 = ~n255 & n641;
  assign n643 = ~q & ~n462;
  assign n644 = ~n640 & ~n643;
  assign n645 = ~n642 & n644;
  assign n646 = n & ~s;
  assign n647 = ~s & ~t;
  assign n648 = o & ~t;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n646 & n649;
  assign n651 = n519 & n521;
  assign n652 = n650 & n651;
  assign n653 = q & n519;
  assign n654 = n650 & n653;
  assign n655 = n205 & n650;
  assign n656 = r & n521;
  assign n657 = n650 & n656;
  assign n658 = ~n655 & ~n657;
  assign n659 = ~n654 & n658;
  assign n660 = ~n652 & n659;
  assign n661 = n518 & n660;
  assign n662 = n645 & n661;
  assign n663 = ~p & n518;
  assign n664 = n645 & n663;
  assign n665 = p & n660;
  assign n666 = n645 & n665;
  assign n667 = ~n664 & ~n666;
  assign n668 = ~n662 & n667;
  assign n669 = i0 & n668;
  assign n670 = ~m & s;
  assign n671 = t & n670;
  assign n672 = ~m & ~r;
  assign n673 = ~n376 & ~n672;
  assign n674 = ~n532 & n673;
  assign n675 = ~n671 & n674;
  assign n676 = s & ~c0;
  assign n677 = n675 & n676;
  assign n678 = s & ~e0;
  assign n679 = n675 & n678;
  assign n680 = t & ~c0;
  assign n681 = n675 & n680;
  assign n682 = t & ~e0;
  assign n683 = n675 & n682;
  assign n684 = ~n681 & ~n683;
  assign n685 = ~n679 & n684;
  assign n686 = ~n677 & n685;
  assign n687 = r & n650;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~n384 & n688;
  assign n690 = ~n525 & ~n526;
  assign n691 = ~l & n272;
  assign n692 = t & n691;
  assign n693 = ~n376 & ~n692;
  assign n694 = ~n532 & n693;
  assign n695 = s & c0;
  assign n696 = n694 & n695;
  assign n697 = s & d0;
  assign n698 = n694 & n697;
  assign n699 = t & c0;
  assign n700 = n694 & n699;
  assign n701 = t & d0;
  assign n702 = n694 & n701;
  assign n703 = ~n700 & ~n702;
  assign n704 = ~n698 & n703;
  assign n705 = ~n696 & n704;
  assign n706 = q & n690;
  assign n707 = ~n643 & ~n705;
  assign n708 = ~n706 & n707;
  assign n709 = f0 & g0;
  assign n710 = l & ~q;
  assign n711 = n462 & n710;
  assign n712 = ~e0 & n711;
  assign n713 = n255 & n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = n631 & ~n714;
  assign n716 = q & n631;
  assign n717 = n689 & n716;
  assign n718 = e0 & n709;
  assign n719 = n708 & n718;
  assign n720 = ~n715 & ~n719;
  assign n721 = ~n717 & n720;
  assign n722 = ~n384 & ~n565;
  assign n723 = n631 & n722;
  assign n724 = ~n255 & n718;
  assign n725 = ~n723 & ~n724;
  assign n726 = t & ~i0;
  assign n727 = k & ~p;
  assign n728 = n726 & n727;
  assign n729 = n721 & n725;
  assign n730 = ~n669 & n729;
  assign n731 = ~n277 & n721;
  assign n732 = ~n669 & n731;
  assign n733 = n721 & ~n728;
  assign n734 = ~n669 & n733;
  assign n735 = ~p & n725;
  assign n736 = ~n669 & n735;
  assign n737 = ~p & ~n277;
  assign n738 = ~n669 & n737;
  assign n739 = ~p & ~n728;
  assign n740 = ~n669 & n739;
  assign n741 = i0 & n725;
  assign n742 = ~n669 & n741;
  assign n743 = i0 & ~n277;
  assign n744 = ~n669 & n743;
  assign n745 = i0 & ~n728;
  assign n746 = ~n669 & n745;
  assign n747 = ~n744 & ~n746;
  assign n748 = ~n742 & n747;
  assign n749 = ~n740 & n748;
  assign n750 = ~n738 & n749;
  assign n751 = ~n736 & n750;
  assign n752 = ~n734 & n751;
  assign n753 = ~n732 & n752;
  assign n754 = ~n730 & n753;
  assign s0 = n627 & n754;
  assign j0 = ~h0;
endmodule


