// Benchmark "TOP" written by ABC on Sun Apr 24 20:32:30 2016

module TOP ( clock, 
    PCLK, PRESET, Preset_0_0_, Pinp_0_0_, Pinp_1_1_, Pinp_2_2_, Pinp_3_3_,
    Pinp_4_4_, Pinp_5_5_, Pinp_6_6_, Pinp_7_7_, Pinp_8_8_, Pinp_9_9_,
    Pinp_10_10_, Pinp_11_11_, Pinp_12_12_, Pinp_13_13_, Pinp_14_14_,
    Pinp_15_15_,
    PDN, Pover_0_0_  );
  input  clock;
  input  PCLK, PRESET, Preset_0_0_, Pinp_0_0_, Pinp_1_1_, Pinp_2_2_,
    Pinp_3_3_, Pinp_4_4_, Pinp_5_5_, Pinp_6_6_, Pinp_7_7_, Pinp_8_8_,
    Pinp_9_9_, Pinp_10_10_, Pinp_11_11_, Pinp_12_12_, Pinp_13_13_,
    Pinp_14_14_, Pinp_15_15_;
  output PDN, Pover_0_0_;
  reg N_N8199, N_N9280, N_N8803, N_N8240, N_N8274, N_N8198, N_N8239,
    N_N8615, N_N7703, N_N8273, N_N8366, N_N8272, N_N8238, N_N8531, N_N7983,
    N_N8575, N_N7854, N_N8237, N_N8197, N_N8271, N_N8530, N_N8650, N_N7985,
    N_N8710, N_N8574, N_N8312, N_N8270, N_N8573, N_N8935, N_N8649, N_N8196,
    N_N8236, N_N9244, N_N8348, N_N9150, N_N8648, N_N8269, N_N8235, N_N9275,
    N_N8970, N_N9554, N_N9013, N_N8508, N_N8529, N_N9242, N_N8572, N_N8571,
    N_N9436, N_N8528, N_N8796, N_N7770, N_N9357, N_N8685, N_N9296, N_N9555,
    N_N7628, N_N9510, N_N9578, N_N8447, N_N9437, N_N7771, N_N8570, N_N8647,
    N_N7704, N_N8646, N_N7629, NDN3_11, NDN3_12, N_N8037, NDN3_16, NDN3_17,
    NDN3_19, NDN3_22, NDN3_25, NDN3_26, N_N7584, NDN3_28, NDN3_29, NDN3_40,
    NDN3_39, NDN3_42, NDN3_44, NDN3_46, N_N9358, N_N9539, N_N9556, N_N7306,
    NEN3_16, N_N9160, NEN3_19, NEN3_22, N_N8930, NEN3_28, N_N9438, NEN3_34,
    NEN3_36, NEN3_39, N_N7961, NLC1_2, N_N9359, N_N7476, N_N8577, N_N9289,
    N_N9557, N_N7630, N_N9161, N_N8691, N_N9439, N_N8798, N_N8869, N_N9360,
    N_N8911, N_N9290, N_N9558, N_N8993, N_N9162, N_N9034, N_N9440, N_N9361,
    N_N9298, N_N9559, N_N9163, N_N9550, PDN, N_N8171, N_N8173, N_N9011,
    N_N9552, N_N7701, N_N8964, N_N9291, N_N9560, N_N7627, N_N8913, N_N8756,
    N_N9164, N_N8016, N_N9441, N_N8847, N_N8631, N_N9362, Pover_0_0_,
    NDN1_4, N_N8561, N_N9292, N_N9561, NGFDN_3, N_N9165, N_N9442, N_N7768,
    N_N8118, NDN2_2, N_N8875, N_N7852, N_N7582, N_N9331, N_N9363, N_N9294,
    NDN3_2, NDN3_4, NDN3_7, NDN3_9, N_N9410, N_N8613, N_N8972, N_N9247,
    N_N9166, N_N8968, NAK3_13, N_N8668, N_N8923, N_N7769, N_N8933, N_N7702,
    N_N8978, N_N8141, N_N8200, N_N8929, N_N7853, N_N9031, N_N8241, N_N7583,
    NSr3_13, N_N9248, NSr3_14, NSr3_20, N_N9198, NSr3_23, NSr3_30, NSr3_35,
    NSr3_37, NSr3_38, NSr1_2, N_N8603;
  wire n604_1, n605, n606, n607, n665, n675, n676, n678_1, n681, n683_1,
    n685, n687, n689, n691, n694, n696, n698_1, n700, n702, n704, n706,
    n711, n712, n713_1, n714, n715, n716, n717, n718_1, n719, n720, n721,
    n722, n723_1, n724, n725, n726, n727, n728_1, n729, n730, n731, n732,
    n733_1, n734, n735, n736, n737, n738_1, n739, n740, n741, n742, n744,
    n746, n748_1, n750, n752_1, n753, n754, n755, n756, n757_1, n758, n759,
    n760, n761, n762_1, n763, n764, n765, n766, n767_1, n768, n769, n770,
    n771, n772_1, n773, n774, n775, n776, n777_1, n778, n779, n780, n781,
    n782_1, n783, n784, n785, n786, n787_1, n788, n789, n790, n791, n792_1,
    n793, n794, n795, n796, n797_1, n798, n799, n800, n801, n802_1, n803,
    n804, n805, n806, n807_1, n808, n809, n810, n811, n812_1, n813, n814,
    n815, n816, n817_1, n818, n819, n820, n821, n822_1, n823, n824, n825,
    n826, n827_1, n828, n829, n830, n831, n832_1, n833, n834, n835, n836,
    n837_1, n838, n839, n840, n841, n842_1, n843, n844, n845, n846, n847_1,
    n848, n849, n850, n851, n852_1, n853, n854, n855, n856, n857_1, n858,
    n859, n860, n861, n862_1, n863, n864, n865, n866, n867_1, n868, n869,
    n870, n871, n872_1, n873, n874, n875, n876, n877_1, n878, n879, n880,
    n881, n882_1, n883, n884, n885, n886, n887_1, n888, n889, n890, n891,
    n892_1, n893, n894, n895, n896, n897_1, n898, n899, n900, n901, n902_1,
    n903, n904, n905, n906, n907_1, n908, n909, n910, n911, n912_1, n913,
    n914, n915, n916, n917_1, n918, n919, n920, n921, n922_1, n923, n924,
    n925, n926, n927_1, n928, n929, n930, n931, n932_1, n933, n934, n935,
    n936, n937_1, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947_1, n948, n949, n950, n951, n952_1, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967_1, n968,
    n969, n970, n971, n972_1, n973, n974, n975, n976, n977_1, n978, n979,
    n980, n981, n982_1, n983, n984, n985, n986, n987_1, n988, n989, n990,
    n991, n992_1, n993, n994, n995, n996, n997_1, n998, n999, n1000, n1001,
    n1002_1, n1003, n1004, n1005, n1006, n1007_1, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1032, n1035, n1037, n1039, n1042, n1043, n1046, n1047, n1053, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1103, n1105,
    n1106, n1107, n1108, n1109, n1115, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1133, n1134, n1135, n1136, n1137, n1138,
    n1143, n1144, n1145, n1146, n1147, n1150, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1165, n1166, n1167, n1168,
    n1169, n1172, n1173, n1174, n1177, n1178, n1179, n1180, n1181, n1182,
    n1187, n1199, n1200, n1201, n1202, n1203, n1205, n1207, n1209, n1214,
    n1215, n1216, n1218, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1232, n1233, n1234, n1235, n1236, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1249, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1262, n1263, n1265, n1267, n1268, n1270, n1271, n1274, n1275, n1277,
    n1278, n1280, n1281, n1283, n1284, n1286, n1287, n1289, n1290, n1292,
    n1293, n1294, n1295, n1296, n44, n49, n54, n59, n64, n69, n74, n79,
    n84, n89, n94, n99, n104, n109, n114, n119, n124, n129, n134, n139,
    n144, n149, n154, n159, n164, n169, n174, n179, n184, n189, n194, n199,
    n204, n209, n214, n219, n224, n229, n234, n239, n244, n249, n254, n259,
    n264, n269, n274, n279, n284, n289, n294, n299, n304, n309, n314, n319,
    n324, n329, n334, n339, n344, n349_1, n354, n359, n364, n369, n374,
    n379, n384, n389, n394, n399, n404_1, n409, n414, n419, n424, n429,
    n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489,
    n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549,
    n554, n559, n564, n569, n574, n579, n584_1, n589, n594, n599, n604,
    n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n663,
    n668, n673, n678, n683, n688, n693, n698, n703, n708, n713, n718, n723,
    n728, n733, n738, n743, n748, n752, n757, n762, n767, n772, n777, n782,
    n787, n792, n797, n802, n807, n812, n817, n822, n827, n832, n837, n842,
    n847, n852, n857, n862, n867, n872, n877, n882, n887, n892, n897, n902,
    n907, n912, n917, n922, n927, n932, n937, n942_1, n947, n952, n957_1,
    n962_1, n967, n972, n977, n982, n987, n992, n997, n1002, n1007;
  assign n604_1 = ~NLC1_2 & NSr1_2;
  assign n605 = Preset_0_0_ & n604_1;
  assign n606 = ~NDN2_2 & n605;
  assign n607 = ~PRESET & ~n606;
  assign n44 = N_N8199 & n607;
  assign n49 = N_N9280 & n607;
  assign n54 = N_N8803 & n607;
  assign n59 = N_N8240 & n607;
  assign n64 = N_N8274 & n607;
  assign n69 = N_N8198 & n607;
  assign n74 = N_N8239 & n607;
  assign n79 = N_N8615 & n607;
  assign n84 = N_N7703 & n607;
  assign n89 = N_N8273 & n607;
  assign n94 = N_N8366 & n607;
  assign n99 = N_N8272 & n607;
  assign n104 = N_N8238 & n607;
  assign n109 = N_N8531 & n607;
  assign n114 = N_N7983 & n607;
  assign n119 = N_N8575 & n607;
  assign n124 = N_N7854 & n607;
  assign n129 = N_N8237 & n607;
  assign n134 = N_N8197 & n607;
  assign n139 = N_N8271 & n607;
  assign n144 = N_N8530 & n607;
  assign n149 = N_N8650 & n607;
  assign n154 = N_N7985 & n607;
  assign n159 = N_N8710 & n607;
  assign n164 = N_N8574 & n607;
  assign n169 = N_N8312 & n607;
  assign n174 = N_N8270 & n607;
  assign n179 = N_N8573 & n607;
  assign n184 = N_N8935 & n607;
  assign n189 = N_N8649 & n607;
  assign n194 = N_N8196 & n607;
  assign n199 = N_N8236 & n607;
  assign n204 = N_N9244 & n607;
  assign n209 = N_N8348 & n607;
  assign n214 = N_N9150 & n607;
  assign n219 = N_N8648 & n607;
  assign n224 = N_N8269 & n607;
  assign n229 = N_N8235 & n607;
  assign n234 = N_N9275 & n607;
  assign n239 = N_N8970 & n607;
  assign n244 = N_N9554 & n607;
  assign n249 = N_N9013 & n607;
  assign n254 = N_N8508 & n607;
  assign n259 = N_N8529 & n607;
  assign n264 = N_N9242 & n607;
  assign n269 = N_N8572 & n607;
  assign n274 = N_N8571 & n607;
  assign n279 = N_N9436 & n607;
  assign n284 = N_N8528 & n607;
  assign n289 = N_N8796 & n607;
  assign n294 = N_N7770 & n607;
  assign n299 = N_N9357 & n607;
  assign n304 = N_N8685 & n607;
  assign n309 = N_N9296 & n607;
  assign n314 = N_N9555 & n607;
  assign n319 = N_N7628 & n607;
  assign n324 = N_N9510 & n607;
  assign n665 = ~N_N9578 & ~n606;
  assign n329 = ~PRESET & ~n665;
  assign n334 = N_N8447 & n607;
  assign n339 = N_N9437 & n607;
  assign n344 = N_N7771 & n607;
  assign n349_1 = N_N8570 & n607;
  assign n354 = N_N8647 & n607;
  assign n359 = N_N7704 & n607;
  assign n364 = N_N8646 & n607;
  assign n369 = N_N7629 & n607;
  assign n675 = ~PRESET & ~NGFDN_3;
  assign n676 = ~NDN3_11 & ~NDN3_9;
  assign n374 = n675 & ~n676;
  assign n678_1 = ~NDN3_11 & ~NDN3_12;
  assign n379 = n675 & ~n678_1;
  assign n384 = N_N8037 & n607;
  assign n681 = ~NDN3_16 & ~NEN3_16;
  assign n389 = n675 & ~n681;
  assign n683_1 = ~NDN3_16 & ~NDN3_17;
  assign n394 = n675 & ~n683_1;
  assign n685 = ~NDN3_19 & ~NEN3_19;
  assign n399 = n675 & ~n685;
  assign n687 = ~NDN3_22 & ~NEN3_22;
  assign n404_1 = n675 & ~n687;
  assign n689 = ~NDN3_22 & ~NDN3_25;
  assign n409 = n675 & ~n689;
  assign n691 = ~NDN3_25 & ~NDN3_26;
  assign n414 = n675 & ~n691;
  assign n419 = N_N7584 & n607;
  assign n694 = ~NDN3_28 & ~NEN3_28;
  assign n424 = n675 & ~n694;
  assign n696 = ~NDN3_28 & ~NDN3_29;
  assign n429 = n675 & ~n696;
  assign n698_1 = ~NDN3_40 & ~NDN3_39;
  assign n434 = n675 & ~n698_1;
  assign n700 = ~NDN3_39 & ~NEN3_39;
  assign n439 = n675 & ~n700;
  assign n702 = ~NDN3_40 & ~NDN3_42;
  assign n444 = n675 & ~n702;
  assign n704 = ~NDN3_42 & ~NDN3_44;
  assign n449 = n675 & ~n704;
  assign n706 = ~NDN3_44 & ~NDN3_46;
  assign n454 = n675 & ~n706;
  assign n459 = N_N9358 & n607;
  assign n464 = N_N9539 & n607;
  assign n469 = N_N9556 & n607;
  assign n711 = ~N_N8847 & ~N_N8631;
  assign n712 = ~N_N8798 & N_N8603;
  assign n713_1 = ~N_N8923 & n712;
  assign n714 = ~N_N8911 & ~N_N8933;
  assign n715 = ~N_N8869 & n714;
  assign n716 = n713_1 & n715;
  assign n717 = ~N_N8978 & n716;
  assign n718_1 = ~N_N8993 & n717;
  assign n719 = ~N_N9031 & n718_1;
  assign n720 = ~N_N9034 & n719;
  assign n721 = ~N_N8561 & n720;
  assign n722 = n711 & n721;
  assign n723_1 = ~N_N8913 & n722;
  assign n724 = N_N8913 & ~n722;
  assign n725 = ~n723_1 & ~n724;
  assign n726 = ~N_N8561 & ~N_N8978;
  assign n727 = ~N_N8798 & ~N_N8993;
  assign n728_1 = n711 & n727;
  assign n729 = ~N_N8964 & n728_1;
  assign n730 = n726 & n729;
  assign n731 = N_N9247 & N_N9248;
  assign n732 = ~N_N7306 & n731;
  assign n733_1 = ~N_N8603 & n732;
  assign n734 = ~N_N9011 & ~N_N8923;
  assign n735 = ~N_N9031 & n734;
  assign n736 = n715 & n735;
  assign n737 = n733_1 & n736;
  assign n738_1 = n730 & n737;
  assign n739 = N_N9034 & ~n719;
  assign n740 = ~n720 & ~n739;
  assign n741 = n738_1 & n740;
  assign n742 = n725 & n741;
  assign n474 = ~PRESET & n742;
  assign n744 = ~NEN3_16 & NSr3_14;
  assign n479 = n675 & ~n744;
  assign n746 = ~N_N9160 & ~n606;
  assign n484 = ~PRESET & ~n746;
  assign n748_1 = ~NEN3_19 & NSr3_20;
  assign n489 = n675 & ~n748_1;
  assign n750 = ~NEN3_22 & NSr3_23;
  assign n494 = n675 & ~n750;
  assign n752_1 = NDN3_12 & NSr3_13;
  assign n753 = NDN3_17 & NSr3_20;
  assign n754 = ~n752_1 & ~n753;
  assign n755 = ~NSr3_13 & NSr3_14;
  assign n756 = NDN3_26 & NSr3_30;
  assign n757_1 = ~n755 & ~n756;
  assign n758 = NDN3_19 & NSr3_23;
  assign n759 = NDN3_29 & NSr3_35;
  assign n760 = ~n758 & ~n759;
  assign n761 = n757_1 & n760;
  assign n762_1 = NEN3_34 & NSr3_37;
  assign n763 = NEN3_36 & NSr3_38;
  assign n764 = ~n762_1 & ~n763;
  assign n765 = n761 & n764;
  assign n766 = n754 & n765;
  assign n767_1 = N_N8930 & ~N_N8929;
  assign n768 = N_N9559 & n753;
  assign n769 = N_N9555 & n762_1;
  assign n770 = N_N9557 & n756;
  assign n771 = ~n769 & ~n770;
  assign n772_1 = N_N9560 & n755;
  assign n773 = n771 & ~n772_1;
  assign n774 = ~n768 & n773;
  assign n775 = N_N9556 & n759;
  assign n776 = N_N9554 & n763;
  assign n777_1 = ~n775 & ~n776;
  assign n778 = N_N9558 & n758;
  assign n779 = N_N9561 & n752_1;
  assign n780 = ~n778 & ~n779;
  assign n781 = n777_1 & n780;
  assign n782_1 = n774 & n781;
  assign n783 = N_N7583 & n756;
  assign n784 = N_N7584 & n755;
  assign n785 = N_N7985 & n758;
  assign n786 = ~n784 & ~n785;
  assign n787_1 = N_N8016 & n763;
  assign n788 = n786 & ~n787_1;
  assign n789 = ~n783 & n788;
  assign n790 = N_N8691 & n752_1;
  assign n791 = N_N7582 & n762_1;
  assign n792_1 = ~n790 & ~n791;
  assign n793 = N_N8447 & n753;
  assign n794 = N_N8968 & n759;
  assign n795 = ~n793 & ~n794;
  assign n796 = n792_1 & n795;
  assign n797_1 = n789 & n796;
  assign n798 = n782_1 & n797_1;
  assign n799 = N_N9552 & n753;
  assign n800 = N_N9359 & n759;
  assign n801 = N_N9361 & n758;
  assign n802_1 = ~n800 & ~n801;
  assign n803 = N_N9360 & n756;
  assign n804 = n802_1 & ~n803;
  assign n805 = ~n799 & n804;
  assign n806 = N_N9358 & n762_1;
  assign n807_1 = N_N9362 & n755;
  assign n808 = ~n806 & ~n807_1;
  assign n809 = N_N9363 & n752_1;
  assign n810 = N_N9357 & n763;
  assign n811 = ~n809 & ~n810;
  assign n812_1 = n808 & n811;
  assign n813 = n805 & n812_1;
  assign n814 = N_N7768 & n762_1;
  assign n815 = N_N7771 & n755;
  assign n816 = N_N7770 & n753;
  assign n817_1 = ~n815 & ~n816;
  assign n818 = N_N7769 & n756;
  assign n819 = n817_1 & ~n818;
  assign n820 = ~n814 & n819;
  assign n821 = N_N8803 & n758;
  assign n822_1 = N_N8173 & n763;
  assign n823 = ~n821 & ~n822_1;
  assign n824 = N_N7961 & n752_1;
  assign n825 = N_N9331 & n759;
  assign n826 = ~n824 & ~n825;
  assign n827_1 = n823 & n826;
  assign n828 = n820 & n827_1;
  assign n829 = ~N_N8930 & n828;
  assign n830 = n813 & n829;
  assign n831 = n798 & n830;
  assign n832_1 = N_N8796 & n759;
  assign n833 = N_N8648 & n753;
  assign n834 = N_N8649 & n755;
  assign n835 = ~n833 & ~n834;
  assign n836 = N_N8650 & n752_1;
  assign n837_1 = n835 & ~n836;
  assign n838 = ~n832_1 & n837_1;
  assign n839 = N_N8646 & n763;
  assign n840 = N_N9242 & n756;
  assign n841 = ~n839 & ~n840;
  assign n842_1 = N_N9013 & n758;
  assign n843 = N_N8647 & n762_1;
  assign n844 = ~n842_1 & ~n843;
  assign n845 = n841 & n844;
  assign n846 = n838 & n845;
  assign n847_1 = N_N8530 & n753;
  assign n848 = N_N8935 & n758;
  assign n849 = N_N9244 & n756;
  assign n850 = ~n848 & ~n849;
  assign n851 = N_N8531 & n755;
  assign n852_1 = n850 & ~n851;
  assign n853 = ~n847_1 & n852_1;
  assign n854 = N_N8528 & n763;
  assign n855 = N_N9275 & n759;
  assign n856 = ~n854 & ~n855;
  assign n857_1 = N_N8615 & n752_1;
  assign n858 = N_N8529 & n762_1;
  assign n859 = ~n857_1 & ~n858;
  assign n860 = n856 & n859;
  assign n861 = n853 & n860;
  assign n862_1 = n846 & n861;
  assign n863 = N_N7701 & n763;
  assign n864 = N_N7703 & n758;
  assign n865 = ~n863 & ~n864;
  assign n866 = N_N7702 & n756;
  assign n867_1 = n865 & ~n866;
  assign n868 = N_N7704 & n755;
  assign n869 = N_N8577 & n752_1;
  assign n870 = ~n868 & ~n869;
  assign n871 = N_N9294 & n759;
  assign n872_1 = n870 & ~n871;
  assign n873 = N_N8685 & n753;
  assign n874 = N_N8118 & n762_1;
  assign n875 = ~n873 & ~n874;
  assign n876 = n872_1 & n875;
  assign n877_1 = n867_1 & n876;
  assign n878 = N_N9410 & n752_1;
  assign n879 = N_N9539 & n762_1;
  assign n880 = ~n878 & ~n879;
  assign n881 = N_N9298 & n758;
  assign n882_1 = n880 & ~n881;
  assign n883 = N_N9291 & n753;
  assign n884 = N_N9289 & n759;
  assign n885 = ~n883 & ~n884;
  assign n886 = N_N9296 & n763;
  assign n887_1 = n885 & ~n886;
  assign n888 = N_N9292 & n755;
  assign n889 = N_N9290 & n756;
  assign n890 = ~n888 & ~n889;
  assign n891 = n887_1 & n890;
  assign n892_1 = n882_1 & n891;
  assign n893 = n877_1 & n892_1;
  assign n894 = n862_1 & n893;
  assign n895 = N_N8236 & n762_1;
  assign n896 = N_N8312 & n759;
  assign n897_1 = ~n895 & ~n896;
  assign n898 = N_N8237 & n756;
  assign n899 = n897_1 & ~n898;
  assign n900 = N_N8241 & n752_1;
  assign n901 = N_N8235 & n763;
  assign n902_1 = ~n900 & ~n901;
  assign n903 = N_N8240 & n755;
  assign n904 = n902_1 & ~n903;
  assign n905 = N_N8238 & n758;
  assign n906 = N_N8239 & n753;
  assign n907_1 = ~n905 & ~n906;
  assign n908 = n904 & n907_1;
  assign n909 = n899 & n908;
  assign n910 = N_N7629 & n755;
  assign n911 = N_N8875 & n762_1;
  assign n912_1 = ~n910 & ~n911;
  assign n913 = N_N7983 & n758;
  assign n914 = n912_1 & ~n913;
  assign n915 = N_N8613 & n759;
  assign n916 = N_N7628 & n753;
  assign n917_1 = ~n915 & ~n916;
  assign n918 = N_N7627 & n763;
  assign n919 = n917_1 & ~n918;
  assign n920 = N_N7630 & n752_1;
  assign n921 = N_N8141 & n756;
  assign n922_1 = ~n920 & ~n921;
  assign n923 = n919 & n922_1;
  assign n924 = n914 & n923;
  assign n925 = N_N8272 & n753;
  assign n926 = N_N8269 & n762_1;
  assign n927_1 = ~n925 & ~n926;
  assign n928 = N_N8348 & n759;
  assign n929 = n927_1 & ~n928;
  assign n930 = N_N8273 & n755;
  assign n931 = N_N8508 & n763;
  assign n932_1 = ~n930 & ~n931;
  assign n933 = N_N8270 & n756;
  assign n934 = n932_1 & ~n933;
  assign n935 = N_N8274 & n752_1;
  assign n936 = N_N8271 & n758;
  assign n937_1 = ~n935 & ~n936;
  assign n938 = n934 & n937_1;
  assign n939 = n929 & n938;
  assign n940 = n924 & n939;
  assign n941 = n909 & n940;
  assign n942 = n894 & n941;
  assign n943 = N_N9165 & n755;
  assign n944 = N_N9578 & n763;
  assign n945 = N_N9162 & n756;
  assign n946 = ~n944 & ~n945;
  assign n947_1 = N_N9166 & n752_1;
  assign n948 = n946 & ~n947_1;
  assign n949 = ~n943 & n948;
  assign n950 = N_N9161 & n759;
  assign n951 = N_N9163 & n758;
  assign n952_1 = ~n950 & ~n951;
  assign n953 = N_N9164 & n753;
  assign n954 = N_N9160 & n762_1;
  assign n955 = ~n953 & ~n954;
  assign n956 = n952_1 & n955;
  assign n957 = n949 & n956;
  assign n958 = N_N7854 & n753;
  assign n959 = N_N7853 & n758;
  assign n960 = N_N9510 & n755;
  assign n961 = ~n959 & ~n960;
  assign n962 = N_N7852 & n759;
  assign n963 = n961 & ~n962;
  assign n964 = ~n958 & n963;
  assign n965 = N_N8972 & n756;
  assign n966 = N_N8037 & n752_1;
  assign n967_1 = ~n965 & ~n966;
  assign n968 = N_N8171 & n763;
  assign n969 = N_N8756 & n762_1;
  assign n970 = ~n968 & ~n969;
  assign n971 = n967_1 & n970;
  assign n972_1 = n964 & n971;
  assign n973 = n957 & n972_1;
  assign n974 = N_N9438 & n759;
  assign n975 = N_N9440 & n758;
  assign n976 = N_N9437 & n762_1;
  assign n977_1 = ~n975 & ~n976;
  assign n978 = N_N9442 & n752_1;
  assign n979 = n977_1 & ~n978;
  assign n980 = ~n974 & n979;
  assign n981 = N_N9436 & n763;
  assign n982_1 = N_N9550 & n753;
  assign n983 = ~n981 & ~n982_1;
  assign n984 = N_N9439 & n756;
  assign n985 = N_N9441 & n755;
  assign n986 = ~n984 & ~n985;
  assign n987_1 = n983 & n986;
  assign n988 = n980 & n987_1;
  assign n989 = N_N8199 & n755;
  assign n990 = N_N8710 & n762_1;
  assign n991 = N_N8366 & n756;
  assign n992_1 = ~n990 & ~n991;
  assign n993 = N_N8200 & n752_1;
  assign n994 = n992_1 & ~n993;
  assign n995 = ~n989 & n994;
  assign n996 = N_N8197 & n759;
  assign n997_1 = N_N8196 & n763;
  assign n998 = ~n996 & ~n997_1;
  assign n999 = N_N8198 & n758;
  assign n1000 = N_N9280 & n753;
  assign n1001 = ~n999 & ~n1000;
  assign n1002_1 = n998 & n1001;
  assign n1003 = n995 & n1002_1;
  assign n1004 = N_N8573 & n753;
  assign n1005 = N_N8572 & n759;
  assign n1006 = N_N8574 & n755;
  assign n1007_1 = ~n1005 & ~n1006;
  assign n1008 = N_N8970 & n756;
  assign n1009 = n1007_1 & ~n1008;
  assign n1010 = ~n1004 & n1009;
  assign n1011 = N_N8570 & n763;
  assign n1012 = N_N8571 & n762_1;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = N_N9150 & n758;
  assign n1015 = N_N8575 & n752_1;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = n1013 & n1016;
  assign n1018 = n1010 & n1017;
  assign n1019 = n1003 & n1018;
  assign n1020 = n988 & n1019;
  assign n1021 = n973 & n1020;
  assign n1022 = n942 & n1021;
  assign n1023 = n831 & n1022;
  assign n1024 = ~n767_1 & ~n1023;
  assign n1025 = ~n766 & ~n1024;
  assign n1026 = N_N9198 & ~n1025;
  assign n1027 = ~PRESET & n1026;
  assign n1028 = N_N9198 & n1024;
  assign n1029 = ~n766 & n1028;
  assign n1030 = ~N_N8930 & ~n1029;
  assign n499 = n1027 & ~n1030;
  assign n1032 = ~NEN3_28 & NSr3_30;
  assign n504 = n675 & ~n1032;
  assign n509 = N_N9438 & n607;
  assign n1035 = ~NEN3_34 & NSr3_35;
  assign n514 = n675 & ~n1035;
  assign n1037 = ~NEN3_36 & NSr3_37;
  assign n519 = n675 & ~n1037;
  assign n1039 = ~NEN3_39 & NSr3_38;
  assign n524 = n675 & ~n1039;
  assign n529 = N_N7961 & n607;
  assign n1042 = ~PRESET & ~PDN;
  assign n1043 = ~NLC1_2 & ~NSr1_2;
  assign n534 = n1042 & ~n1043;
  assign n539 = N_N9359 & n607;
  assign n1046 = ~N_N7476 & ~n604_1;
  assign n1047 = ~PRESET & ~n605;
  assign n544 = ~n1046 & n1047;
  assign n549 = N_N8577 & n607;
  assign n554 = N_N9289 & n607;
  assign n559 = N_N9557 & n607;
  assign n564 = N_N7630 & n607;
  assign n1053 = ~N_N9161 & ~n606;
  assign n569 = ~PRESET & ~n1053;
  assign n574 = N_N8691 & n607;
  assign n579 = N_N9439 & n607;
  assign n1057 = ~N_N8668 & ~n1026;
  assign n1058 = n1024 & n1057;
  assign n1059 = ~N_N9247 & n1029;
  assign n1060 = ~n732 & ~n1057;
  assign n1061 = ~n1059 & n1060;
  assign n1062 = ~n1058 & ~n1061;
  assign n1063 = ~n733_1 & n1062;
  assign n1064 = N_N8798 & ~n1063;
  assign n1065 = N_N8603 & n732;
  assign n1066 = ~N_N8798 & n1065;
  assign n1067 = ~n1024 & n1057;
  assign n1068 = ~n1059 & ~n1067;
  assign n1069 = ~n957 & ~n1068;
  assign n1070 = ~n1066 & ~n1069;
  assign n1071 = ~n1064 & n1070;
  assign n584_1 = ~PRESET & ~n1071;
  assign n1073 = ~N_N8869 & n713_1;
  assign n1074 = n732 & n1073;
  assign n1075 = ~n713_1 & n732;
  assign n1076 = n1062 & ~n1075;
  assign n1077 = N_N8869 & ~n1076;
  assign n1078 = ~n892_1 & ~n1068;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = ~n1074 & n1079;
  assign n589 = ~PRESET & ~n1080;
  assign n594 = N_N9360 & n607;
  assign n1083 = ~n813 & ~n1068;
  assign n1084 = n714 & n1074;
  assign n1085 = n732 & ~n1073;
  assign n1086 = n1062 & ~n1085;
  assign n1087 = N_N8933 & n732;
  assign n1088 = n1086 & ~n1087;
  assign n1089 = N_N8911 & ~n1088;
  assign n1090 = ~n1084 & ~n1089;
  assign n1091 = ~n1083 & n1090;
  assign n599 = ~PRESET & ~n1091;
  assign n604 = N_N9290 & n607;
  assign n609 = N_N9558 & n607;
  assign n1095 = N_N8993 & ~n1062;
  assign n1096 = ~n988 & ~n1068;
  assign n1097 = N_N8993 & ~n717;
  assign n1098 = ~n718_1 & ~n1097;
  assign n1099 = n732 & ~n1098;
  assign n1100 = ~n1096 & ~n1099;
  assign n1101 = ~n1095 & n1100;
  assign n614 = ~PRESET & ~n1101;
  assign n1103 = ~N_N9162 & ~n606;
  assign n619 = ~PRESET & ~n1103;
  assign n1105 = n732 & ~n740;
  assign n1106 = N_N9034 & ~n1062;
  assign n1107 = ~n782_1 & ~n1068;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = ~n1105 & n1108;
  assign n624 = ~PRESET & ~n1109;
  assign n629 = N_N9440 & n607;
  assign n634 = N_N9361 & n607;
  assign n639 = N_N9298 & n607;
  assign n644 = N_N9559 & n607;
  assign n1115 = ~N_N9163 & ~n606;
  assign n649 = ~PRESET & ~n1115;
  assign n654 = N_N9550 & n607;
  assign n659 = ~NSr1_2 & n1042;
  assign n663 = N_N8171 & n607;
  assign n668 = N_N8173 & n607;
  assign n1121 = ~N_N8964 & n723_1;
  assign n1122 = n732 & ~n1121;
  assign n1123 = n1062 & ~n1122;
  assign n1124 = N_N9011 & ~n1123;
  assign n1125 = ~n846 & ~n1068;
  assign n1126 = n732 & n1121;
  assign n1127 = ~N_N9011 & n1126;
  assign n1128 = ~n1125 & ~n1127;
  assign n1129 = ~n1124 & n1128;
  assign n673 = ~PRESET & ~n1129;
  assign n678 = N_N9552 & n607;
  assign n683 = N_N7701 & n607;
  assign n1133 = ~n723_1 & n732;
  assign n1134 = n1062 & ~n1133;
  assign n1135 = N_N8964 & ~n1134;
  assign n1136 = ~n1018 & ~n1068;
  assign n1137 = ~n1126 & ~n1136;
  assign n1138 = ~n1135 & n1137;
  assign n688 = ~PRESET & ~n1138;
  assign n693 = N_N9291 & n607;
  assign n698 = N_N9560 & n607;
  assign n703 = N_N7627 & n607;
  assign n1143 = ~n725 & n732;
  assign n1144 = N_N8913 & ~n1062;
  assign n1145 = ~n861 & ~n1068;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1143 & n1146;
  assign n708 = ~PRESET & ~n1147;
  assign n713 = N_N8756 & n607;
  assign n1150 = ~N_N9164 & ~n606;
  assign n718 = ~PRESET & ~n1150;
  assign n723 = N_N8016 & n607;
  assign n728 = N_N9441 & n607;
  assign n1154 = n721 & n732;
  assign n1155 = n711 & n1154;
  assign n1156 = ~n939 & ~n1068;
  assign n1157 = ~n721 & n732;
  assign n1158 = n1062 & ~n1157;
  assign n1159 = N_N8631 & n732;
  assign n1160 = n1158 & ~n1159;
  assign n1161 = N_N8847 & ~n1160;
  assign n1162 = ~n1156 & ~n1161;
  assign n1163 = ~n1155 & n1162;
  assign n733 = ~PRESET & ~n1163;
  assign n1165 = N_N8631 & ~n1158;
  assign n1166 = ~N_N8631 & n1154;
  assign n1167 = ~n909 & ~n1068;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n1165 & n1168;
  assign n738 = ~PRESET & ~n1169;
  assign n743 = N_N9362 & n607;
  assign n1172 = PDN & ~NDN1_4;
  assign n1173 = ~PRESET & Pover_0_0_;
  assign n1174 = ~n1172 & n1173;
  assign n748 = n659 | n1174;
  assign n752 = NDN1_4 & n1042;
  assign n1177 = ~n720 & n732;
  assign n1178 = n1062 & ~n1177;
  assign n1179 = N_N8561 & ~n1178;
  assign n1180 = ~n1003 & ~n1068;
  assign n1181 = ~n1154 & ~n1180;
  assign n1182 = ~n1179 & n1181;
  assign n757 = ~PRESET & ~n1182;
  assign n762 = N_N9292 & n607;
  assign n767 = N_N9561 & n607;
  assign n772 = NDN3_46 & n675;
  assign n1187 = ~N_N9165 & ~n606;
  assign n777 = ~PRESET & ~n1187;
  assign n782 = N_N9442 & n607;
  assign n787 = N_N7768 & n607;
  assign n792 = N_N8118 & n607;
  assign n797 = NDN2_2 & n1047;
  assign n802 = N_N8875 & n607;
  assign n807 = N_N7852 & n607;
  assign n812 = N_N7582 & n607;
  assign n817 = N_N9331 & n607;
  assign n822 = N_N9363 & n607;
  assign n827 = N_N9294 & n607;
  assign n1199 = NLC1_2 & NSr1_2;
  assign n1200 = N_N7476 & n1199;
  assign n1201 = ~Preset_0_0_ & n604_1;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~NDN3_2 & n1202;
  assign n832 = n675 & ~n1203;
  assign n1205 = ~NDN3_2 & ~NDN3_4;
  assign n837 = n675 & ~n1205;
  assign n1207 = ~NDN3_4 & ~NDN3_7;
  assign n842 = n675 & ~n1207;
  assign n1209 = ~NDN3_7 & ~NDN3_9;
  assign n847 = n675 & ~n1209;
  assign n852 = N_N9410 & n607;
  assign n857 = N_N8613 & n607;
  assign n862 = N_N8972 & n607;
  assign n1214 = N_N9247 & ~n742;
  assign n1215 = ~n1059 & ~n1214;
  assign n1216 = N_N9248 & ~n1215;
  assign n867 = ~PRESET & n1216;
  assign n1218 = ~N_N9166 & ~n606;
  assign n872 = ~PRESET & ~n1218;
  assign n877 = N_N8968 & n607;
  assign n882 = ~PRESET & ~n1026;
  assign n887 = N_N8668 & n1027;
  assign n1223 = ~n712 & n732;
  assign n1224 = n1062 & ~n1223;
  assign n1225 = N_N8923 & ~n1224;
  assign n1226 = ~N_N8923 & n1066;
  assign n1227 = ~n924 & ~n1068;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1225 & n1228;
  assign n892 = ~PRESET & ~n1229;
  assign n897 = N_N7769 & n607;
  assign n1232 = N_N8933 & ~n1086;
  assign n1233 = ~N_N8933 & n1074;
  assign n1234 = ~n877_1 & ~n1068;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1232 & n1235;
  assign n902 = ~PRESET & ~n1236;
  assign n907 = N_N7702 & n607;
  assign n1239 = N_N8978 & ~n1062;
  assign n1240 = ~n828 & ~n1068;
  assign n1241 = N_N8978 & ~n716;
  assign n1242 = ~n717 & ~n1241;
  assign n1243 = n732 & ~n1242;
  assign n1244 = ~n1240 & ~n1243;
  assign n1245 = ~n1239 & n1244;
  assign n912 = ~PRESET & ~n1245;
  assign n917 = N_N8141 & n607;
  assign n922 = N_N8200 & n607;
  assign n1249 = ~N_N8929 & ~n1029;
  assign n927 = ~PRESET & ~n1249;
  assign n932 = N_N7853 & n607;
  assign n1252 = ~n972_1 & ~n1068;
  assign n1253 = n719 & n732;
  assign n1254 = ~n718_1 & n732;
  assign n1255 = n1062 & ~n1254;
  assign n1256 = N_N9031 & ~n1255;
  assign n1257 = ~n1253 & ~n1256;
  assign n1258 = ~n1252 & n1257;
  assign n937 = ~PRESET & ~n1258;
  assign n942_1 = N_N8241 & n607;
  assign n947 = N_N7583 & n607;
  assign n1262 = NDN3_12 & NAK3_13;
  assign n1263 = NSr3_13 & ~n1262;
  assign n952 = ~n1042 | n1263;
  assign n1265 = N_N9248 & ~n742;
  assign n957_1 = ~n1027 | n1265;
  assign n1267 = NAK3_13 & ~NSr3_13;
  assign n1268 = NSr3_14 & ~n1267;
  assign n962_1 = ~n1042 | n1268;
  assign n1270 = NDN3_17 & NAK3_13;
  assign n1271 = NSr3_20 & ~n1270;
  assign n967 = ~n1042 | n1271;
  assign n972 = n766 | n957_1;
  assign n1274 = NDN3_19 & NAK3_13;
  assign n1275 = NSr3_23 & ~n1274;
  assign n977 = ~n1042 | n1275;
  assign n1277 = NDN3_26 & NAK3_13;
  assign n1278 = NSr3_30 & ~n1277;
  assign n982 = ~n1042 | n1278;
  assign n1280 = NDN3_29 & NAK3_13;
  assign n1281 = NSr3_35 & ~n1280;
  assign n987 = ~n1042 | n1281;
  assign n1283 = NEN3_34 & NAK3_13;
  assign n1284 = NSr3_37 & ~n1283;
  assign n992 = ~n1042 | n1284;
  assign n1286 = NEN3_36 & NAK3_13;
  assign n1287 = NSr3_38 & ~n1286;
  assign n997 = ~n1042 | n1287;
  assign n1289 = ~NGFDN_3 & NSr1_2;
  assign n1290 = ~n605 & n1289;
  assign n1002 = ~n1042 | n1290;
  assign n1292 = ~N_N8603 & ~n1062;
  assign n1293 = ~n797_1 & ~n1068;
  assign n1294 = ~n1065 & ~n1293;
  assign n1295 = ~n1061 & ~n1294;
  assign n1296 = ~n1292 & ~n1295;
  assign n1007 = PRESET | n1296;
  always @ (posedge clock) begin
    N_N8199 <= n44;
    N_N9280 <= n49;
    N_N8803 <= n54;
    N_N8240 <= n59;
    N_N8274 <= n64;
    N_N8198 <= n69;
    N_N8239 <= n74;
    N_N8615 <= n79;
    N_N7703 <= n84;
    N_N8273 <= n89;
    N_N8366 <= n94;
    N_N8272 <= n99;
    N_N8238 <= n104;
    N_N8531 <= n109;
    N_N7983 <= n114;
    N_N8575 <= n119;
    N_N7854 <= n124;
    N_N8237 <= n129;
    N_N8197 <= n134;
    N_N8271 <= n139;
    N_N8530 <= n144;
    N_N8650 <= n149;
    N_N7985 <= n154;
    N_N8710 <= n159;
    N_N8574 <= n164;
    N_N8312 <= n169;
    N_N8270 <= n174;
    N_N8573 <= n179;
    N_N8935 <= n184;
    N_N8649 <= n189;
    N_N8196 <= n194;
    N_N8236 <= n199;
    N_N9244 <= n204;
    N_N8348 <= n209;
    N_N9150 <= n214;
    N_N8648 <= n219;
    N_N8269 <= n224;
    N_N8235 <= n229;
    N_N9275 <= n234;
    N_N8970 <= n239;
    N_N9554 <= n244;
    N_N9013 <= n249;
    N_N8508 <= n254;
    N_N8529 <= n259;
    N_N9242 <= n264;
    N_N8572 <= n269;
    N_N8571 <= n274;
    N_N9436 <= n279;
    N_N8528 <= n284;
    N_N8796 <= n289;
    N_N7770 <= n294;
    N_N9357 <= n299;
    N_N8685 <= n304;
    N_N9296 <= n309;
    N_N9555 <= n314;
    N_N7628 <= n319;
    N_N9510 <= n324;
    N_N9578 <= n329;
    N_N8447 <= n334;
    N_N9437 <= n339;
    N_N7771 <= n344;
    N_N8570 <= n349_1;
    N_N8647 <= n354;
    N_N7704 <= n359;
    N_N8646 <= n364;
    N_N7629 <= n369;
    NDN3_11 <= n374;
    NDN3_12 <= n379;
    N_N8037 <= n384;
    NDN3_16 <= n389;
    NDN3_17 <= n394;
    NDN3_19 <= n399;
    NDN3_22 <= n404_1;
    NDN3_25 <= n409;
    NDN3_26 <= n414;
    N_N7584 <= n419;
    NDN3_28 <= n424;
    NDN3_29 <= n429;
    NDN3_40 <= n434;
    NDN3_39 <= n439;
    NDN3_42 <= n444;
    NDN3_44 <= n449;
    NDN3_46 <= n454;
    N_N9358 <= n459;
    N_N9539 <= n464;
    N_N9556 <= n469;
    N_N7306 <= n474;
    NEN3_16 <= n479;
    N_N9160 <= n484;
    NEN3_19 <= n489;
    NEN3_22 <= n494;
    N_N8930 <= n499;
    NEN3_28 <= n504;
    N_N9438 <= n509;
    NEN3_34 <= n514;
    NEN3_36 <= n519;
    NEN3_39 <= n524;
    N_N7961 <= n529;
    NLC1_2 <= n534;
    N_N9359 <= n539;
    N_N7476 <= n544;
    N_N8577 <= n549;
    N_N9289 <= n554;
    N_N9557 <= n559;
    N_N7630 <= n564;
    N_N9161 <= n569;
    N_N8691 <= n574;
    N_N9439 <= n579;
    N_N8798 <= n584_1;
    N_N8869 <= n589;
    N_N9360 <= n594;
    N_N8911 <= n599;
    N_N9290 <= n604;
    N_N9558 <= n609;
    N_N8993 <= n614;
    N_N9162 <= n619;
    N_N9034 <= n624;
    N_N9440 <= n629;
    N_N9361 <= n634;
    N_N9298 <= n639;
    N_N9559 <= n644;
    N_N9163 <= n649;
    N_N9550 <= n654;
    PDN <= n659;
    N_N8171 <= n663;
    N_N8173 <= n668;
    N_N9011 <= n673;
    N_N9552 <= n678;
    N_N7701 <= n683;
    N_N8964 <= n688;
    N_N9291 <= n693;
    N_N9560 <= n698;
    N_N7627 <= n703;
    N_N8913 <= n708;
    N_N8756 <= n713;
    N_N9164 <= n718;
    N_N8016 <= n723;
    N_N9441 <= n728;
    N_N8847 <= n733;
    N_N8631 <= n738;
    N_N9362 <= n743;
    Pover_0_0_ <= n748;
    NDN1_4 <= n752;
    N_N8561 <= n757;
    N_N9292 <= n762;
    N_N9561 <= n767;
    NGFDN_3 <= n772;
    N_N9165 <= n777;
    N_N9442 <= n782;
    N_N7768 <= n787;
    N_N8118 <= n792;
    NDN2_2 <= n797;
    N_N8875 <= n802;
    N_N7852 <= n807;
    N_N7582 <= n812;
    N_N9331 <= n817;
    N_N9363 <= n822;
    N_N9294 <= n827;
    NDN3_2 <= n832;
    NDN3_4 <= n837;
    NDN3_7 <= n842;
    NDN3_9 <= n847;
    N_N9410 <= n852;
    N_N8613 <= n857;
    N_N8972 <= n862;
    N_N9247 <= n867;
    N_N9166 <= n872;
    N_N8968 <= n877;
    NAK3_13 <= n882;
    N_N8668 <= n887;
    N_N8923 <= n892;
    N_N7769 <= n897;
    N_N8933 <= n902;
    N_N7702 <= n907;
    N_N8978 <= n912;
    N_N8141 <= n917;
    N_N8200 <= n922;
    N_N8929 <= n927;
    N_N7853 <= n932;
    N_N9031 <= n937;
    N_N8241 <= n942_1;
    N_N7583 <= n947;
    NSr3_13 <= n952;
    N_N9248 <= n957_1;
    NSr3_14 <= n962_1;
    NSr3_20 <= n967;
    N_N9198 <= n972;
    NSr3_23 <= n977;
    NSr3_30 <= n982;
    NSr3_35 <= n987;
    NSr3_37 <= n992;
    NSr3_38 <= n997;
    NSr1_2 <= n1002;
    N_N8603 <= n1007;
  end
endmodule


