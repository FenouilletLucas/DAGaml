// Benchmark "b9" written by ABC on Tue May 16 16:07:44 2017

module b9 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, p0, q0, r0, s0, t0, u0, v0, w0,
    x0, y0, z0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0;
  output a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, p0, q0, r0, s0, t0, u0, v0,
    w0, x0, y0, z0;
  wire n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n111, n112, n114, n116, n117, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n130, n132, n133, n134, n135,
    n136, n137, n139, n140, n141, n142, n143, n144, n146, n147, n148, n149,
    n152, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n168, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185;
  assign n63 = i & d0;
  assign n64 = o0 & n63;
  assign n65 = i & j0;
  assign n66 = ~c0 & n65;
  assign n67 = ~b0 & n66;
  assign n68 = ~c0 & j0;
  assign n69 = b0 & n68;
  assign n70 = ~e & n69;
  assign n71 = ~j & ~e0;
  assign n72 = ~n70 & n71;
  assign n73 = ~n67 & n72;
  assign n74 = ~n64 & n73;
  assign n75 = ~n0 & n73;
  assign h1 = ~n74 & ~n75;
  assign n77 = c0 & j0;
  assign n78 = ~l0 & ~n77;
  assign n79 = b0 & ~n78;
  assign n80 = c0 & ~k0;
  assign n81 = ~j0 & ~k0;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~e & n82;
  assign n84 = ~e & k;
  assign n85 = ~n83 & ~n84;
  assign n86 = ~b0 & ~n84;
  assign n87 = ~n85 & ~n86;
  assign n88 = o0 & n87;
  assign n89 = ~n0 & ~n79;
  assign n90 = ~n79 & ~n88;
  assign b1 = n89 | n90;
  assign n92 = j0 & k0;
  assign n93 = c0 & ~n92;
  assign n94 = ~e0 & ~g0;
  assign n95 = n93 & n94;
  assign n96 = ~b0 & n94;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~e & o0;
  assign n99 = ~n & n98;
  assign n100 = n97 & n99;
  assign n101 = ~t & u;
  assign n102 = ~s & n101;
  assign n103 = ~j0 & ~l0;
  assign n104 = ~c0 & ~l0;
  assign n105 = ~n103 & ~n104;
  assign n106 = b0 & n105;
  assign n107 = n102 & n106;
  assign n108 = ~n100 & ~n107;
  assign n109 = ~n0 & ~n107;
  assign c1 = ~n108 & ~n109;
  assign n111 = a0 & i0;
  assign n112 = m & b0;
  assign e1 = n111 & n112;
  assign n114 = w & ~x;
  assign f1 = b & n114;
  assign n116 = x & ~y;
  assign n117 = w & n116;
  assign g1 = b & n117;
  assign n119 = i & o0;
  assign n120 = d0 & n119;
  assign n121 = i & ~c0;
  assign n122 = j0 & n121;
  assign n123 = b0 & j0;
  assign n124 = ~n122 & ~n123;
  assign n125 = ~e0 & n124;
  assign n126 = ~j & n125;
  assign n127 = ~n120 & n126;
  assign n128 = ~n0 & n126;
  assign j1 = n127 | n128;
  assign n130 = ~p & ~b1;
  assign p0 = ~q | n130;
  assign n132 = e & ~n94;
  assign n133 = e & n123;
  assign n134 = ~c0 & n133;
  assign n135 = e & b0;
  assign n136 = k0 & n135;
  assign n137 = ~n134 & ~n136;
  assign q0 = ~n132 & n137;
  assign n139 = i & n68;
  assign n140 = ~n69 & ~n139;
  assign n141 = ~c & ~n63;
  assign n142 = e & n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = n0 & n143;
  assign r0 = ~o0 | ~n144;
  assign n146 = b0 & ~n77;
  assign n147 = ~b0 & ~l0;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~n78 & n148;
  assign s0 = ~v | ~n149;
  assign t0 = v | ~n149;
  assign n152 = b0 & c0;
  assign v0 = ~l0 & ~n152;
  assign n154 = ~p & r;
  assign n155 = ~f0 & ~n154;
  assign n156 = ~h0 & n155;
  assign n157 = o & ~n156;
  assign n158 = d & ~n157;
  assign n159 = ~a & o;
  assign n160 = ~a & ~z;
  assign n161 = o & z;
  assign n162 = ~n160 & ~n161;
  assign n163 = ~n159 & n162;
  assign n164 = ~m0 & n158;
  assign n165 = n158 & n163;
  assign w0 = n164 | n165;
  assign x0 = n0 & o0;
  assign n168 = l & b0;
  assign y0 = n111 & n168;
  assign n170 = ~e & h;
  assign n171 = b0 & n170;
  assign n172 = n82 & n171;
  assign n173 = ~n0 & n172;
  assign n174 = ~o0 & n172;
  assign n175 = ~n173 & ~n174;
  assign n176 = o0 & ~n94;
  assign n177 = o0 & n82;
  assign n178 = b0 & n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = ~e & n0;
  assign n181 = ~n179 & n180;
  assign n182 = f & n181;
  assign n183 = g & b0;
  assign n184 = l0 & n183;
  assign n185 = ~n182 & ~n184;
  assign z0 = ~n175 | ~n185;
  assign a1 = ~h1;
  assign d1 = ~c1;
  assign u0 = ~v0;
  assign i1 = a1;
endmodule


