// Benchmark "t481" written by ABC on Tue May 16 16:07:52 2017

module t481 ( 
    v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9,
    \v16.0   );
  input  v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7,
    v8, v9;
  output \v16.0 ;
  wire n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674;
  assign n18 = v2 & ~v3;
  assign n19 = v4 & n18;
  assign n20 = v7 & n19;
  assign n21 = ~v1 & n20;
  assign n22 = ~v8 & n21;
  assign n23 = v0 & n18;
  assign n24 = ~v5 & v7;
  assign n25 = n23 & n24;
  assign n26 = ~v8 & n25;
  assign n27 = ~n22 & ~n26;
  assign n28 = v0 & n20;
  assign n29 = ~v8 & n28;
  assign n30 = v10 & ~v11;
  assign n31 = ~v12 & v13;
  assign n32 = ~v14 & n31;
  assign n33 = n30 & n32;
  assign n34 = n27 & ~n29;
  assign n35 = v9 & n33;
  assign n36 = ~n34 & n35;
  assign n37 = ~v4 & v5;
  assign n38 = v6 & n37;
  assign n39 = n23 & n38;
  assign n40 = ~v7 & n39;
  assign n41 = ~v8 & v9;
  assign n42 = n30 & n41;
  assign n43 = v15 & n31;
  assign n44 = n42 & n43;
  assign n45 = n40 & n44;
  assign n46 = ~v1 & n18;
  assign n47 = n38 & n46;
  assign n48 = ~v7 & n47;
  assign n49 = n44 & n48;
  assign n50 = ~v6 & n19;
  assign n51 = v0 & n50;
  assign n52 = n44 & n51;
  assign n53 = ~v1 & n50;
  assign n54 = n44 & n53;
  assign n55 = n33 & n41;
  assign n56 = ~v0 & v1;
  assign n57 = v3 & n56;
  assign n58 = ~v7 & n57;
  assign n59 = n38 & n58;
  assign n60 = n55 & n59;
  assign n61 = v6 & ~v7;
  assign n62 = n37 & n61;
  assign n63 = ~v2 & n56;
  assign n64 = n62 & n63;
  assign n65 = n55 & n64;
  assign n66 = ~v5 & ~v6;
  assign n67 = n63 & n66;
  assign n68 = n55 & n67;
  assign n69 = v9 & n30;
  assign n70 = v4 & v7;
  assign n71 = ~n18 & n70;
  assign n72 = n56 & n71;
  assign n73 = n22 & n43;
  assign n74 = n69 & n73;
  assign n75 = n55 & n72;
  assign n76 = n29 & n43;
  assign n77 = n69 & n76;
  assign n78 = ~n75 & ~n77;
  assign n79 = ~n74 & n78;
  assign n80 = n23 & n66;
  assign n81 = n46 & n66;
  assign n82 = ~n80 & ~n81;
  assign n83 = n24 & n57;
  assign n84 = n82 & ~n83;
  assign n85 = ~n53 & n84;
  assign n86 = n55 & ~n85;
  assign n87 = v4 & ~v6;
  assign n88 = n57 & n87;
  assign n89 = n24 & n63;
  assign n90 = ~n88 & ~n89;
  assign n91 = n63 & n87;
  assign n92 = n57 & n66;
  assign n93 = ~n91 & ~n92;
  assign n94 = n90 & n93;
  assign n95 = n55 & ~n94;
  assign n96 = n40 & n55;
  assign n97 = n48 & n55;
  assign n98 = n51 & n55;
  assign n99 = n44 & n64;
  assign n100 = n57 & n70;
  assign n101 = n44 & n100;
  assign n102 = n63 & n70;
  assign n103 = n44 & n102;
  assign n104 = ~v10 & v8;
  assign n105 = n32 & n104;
  assign n106 = n28 & n105;
  assign n107 = n21 & n105;
  assign n108 = n40 & n105;
  assign n109 = n44 & n89;
  assign n110 = n44 & n88;
  assign n111 = ~n59 & ~n67;
  assign n112 = n93 & n111;
  assign n113 = n44 & ~n112;
  assign n114 = ~n64 & ~n100;
  assign n115 = n50 & ~n56;
  assign n116 = ~n48 & ~n115;
  assign n117 = n84 & ~n89;
  assign n118 = v11 & v8;
  assign n119 = n32 & n118;
  assign n120 = ~n88 & n93;
  assign n121 = n111 & n120;
  assign n122 = n117 & n121;
  assign n123 = ~n28 & n122;
  assign n124 = n116 & n123;
  assign n125 = n114 & n124;
  assign n126 = ~n28 & ~n105;
  assign n127 = ~n105 & ~n119;
  assign n128 = ~n126 & ~n127;
  assign n129 = ~n125 & n128;
  assign n130 = v11 & ~v9;
  assign n131 = n43 & n130;
  assign n132 = n40 & n131;
  assign n133 = n48 & n131;
  assign n134 = n51 & n131;
  assign n135 = n53 & n131;
  assign n136 = n59 & n119;
  assign n137 = n64 & n119;
  assign n138 = n67 & n119;
  assign n139 = n20 & ~n56;
  assign n140 = n72 & n119;
  assign n141 = n131 & n139;
  assign n142 = ~n140 & ~n141;
  assign n143 = ~n85 & n119;
  assign n144 = ~n94 & n119;
  assign n145 = ~n21 & ~n25;
  assign n146 = n24 & n46;
  assign n147 = ~n40 & ~n146;
  assign n148 = ~n48 & n147;
  assign n149 = ~n51 & n148;
  assign n150 = n102 & n105;
  assign n151 = n119 & ~n145;
  assign n152 = n119 & ~n149;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~n150 & n153;
  assign n155 = ~v10 & ~v9;
  assign n156 = n43 & n155;
  assign n157 = n88 & n156;
  assign n158 = n91 & n156;
  assign n159 = n67 & n156;
  assign n160 = n59 & n156;
  assign n161 = n64 & n156;
  assign n162 = n100 & n156;
  assign n163 = n43 & n104;
  assign n164 = n28 & n163;
  assign n165 = n51 & n156;
  assign n166 = n53 & n156;
  assign n167 = n48 & n156;
  assign n168 = ~n117 & n156;
  assign n169 = ~n83 & n90;
  assign n170 = n131 & ~n169;
  assign n171 = ~n112 & n131;
  assign n172 = ~n64 & ~n72;
  assign n173 = n131 & ~n172;
  assign n174 = n28 & n156;
  assign n175 = ~n173 & ~n174;
  assign n176 = n145 & n147;
  assign n177 = n156 & ~n176;
  assign n178 = n55 & n146;
  assign n179 = ~n81 & ~n83;
  assign n180 = ~n80 & n179;
  assign n181 = ~n146 & n180;
  assign n182 = ~n25 & n181;
  assign n183 = ~n177 & n182;
  assign n184 = n175 & n183;
  assign n185 = ~n171 & n184;
  assign n186 = ~n170 & n185;
  assign n187 = ~n168 & n186;
  assign n188 = ~n167 & n187;
  assign n189 = ~n166 & n188;
  assign n190 = ~n165 & n189;
  assign n191 = ~n164 & n190;
  assign n192 = ~n162 & n191;
  assign n193 = ~n161 & n192;
  assign n194 = ~n160 & n193;
  assign n195 = ~n159 & n194;
  assign n196 = ~n158 & n195;
  assign n197 = ~n157 & n196;
  assign n198 = n154 & n197;
  assign n199 = ~n144 & n198;
  assign n200 = ~n143 & n199;
  assign n201 = n142 & n200;
  assign n202 = ~n138 & n201;
  assign n203 = ~n137 & n202;
  assign n204 = ~n136 & n203;
  assign n205 = ~n135 & n204;
  assign n206 = ~n134 & n205;
  assign n207 = ~n133 & n206;
  assign n208 = ~n132 & n207;
  assign n209 = ~n92 & n208;
  assign n210 = ~n129 & n209;
  assign n211 = ~n113 & n210;
  assign n212 = ~n110 & n211;
  assign n213 = ~n109 & n212;
  assign n214 = ~n108 & n213;
  assign n215 = ~n107 & n214;
  assign n216 = ~n106 & n215;
  assign n217 = ~n103 & n216;
  assign n218 = ~n101 & n217;
  assign n219 = ~n99 & n218;
  assign n220 = ~n98 & n219;
  assign n221 = ~n97 & n220;
  assign n222 = ~n96 & n221;
  assign n223 = ~n95 & n222;
  assign n224 = ~n86 & n223;
  assign n225 = n79 & n224;
  assign n226 = ~n68 & n225;
  assign n227 = ~n65 & n226;
  assign n228 = ~n60 & n227;
  assign n229 = ~n54 & n228;
  assign n230 = ~n52 & n229;
  assign n231 = ~n49 & n230;
  assign n232 = ~n45 & n231;
  assign n233 = ~n36 & n232;
  assign n234 = n154 & ~n164;
  assign n235 = ~n144 & n234;
  assign n236 = ~n143 & n235;
  assign n237 = n142 & n236;
  assign n238 = ~n138 & n237;
  assign n239 = ~n137 & n238;
  assign n240 = ~n136 & n239;
  assign n241 = ~n129 & n240;
  assign n242 = ~n98 & n241;
  assign n243 = ~n97 & n242;
  assign n244 = ~n96 & n243;
  assign n245 = ~n178 & n244;
  assign n246 = ~n95 & n245;
  assign n247 = ~n86 & n246;
  assign n248 = n79 & n247;
  assign n249 = ~n68 & n248;
  assign n250 = ~n65 & n249;
  assign n251 = ~n60 & n250;
  assign n252 = ~n36 & n251;
  assign n253 = ~n156 & n252;
  assign n254 = ~n105 & n253;
  assign n255 = ~n44 & n254;
  assign n256 = ~n131 & n255;
  assign n257 = ~n233 & ~n256;
  assign n258 = n32 & n130;
  assign n259 = ~n112 & n258;
  assign n260 = n43 & n118;
  assign n261 = n40 & n260;
  assign n262 = n48 & n260;
  assign n263 = n51 & n260;
  assign n264 = n53 & n260;
  assign n265 = n59 & n163;
  assign n266 = n64 & n163;
  assign n267 = n67 & n163;
  assign n268 = n72 & n104;
  assign n269 = n118 & n139;
  assign n270 = ~n268 & ~n269;
  assign n271 = n43 & ~n270;
  assign n272 = n104 & ~n145;
  assign n273 = n102 & n156;
  assign n274 = n43 & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = ~n149 & n163;
  assign n277 = ~n85 & n163;
  assign n278 = ~n94 & n163;
  assign n279 = v14 & ~v15;
  assign n280 = ~v13 & n279;
  assign n281 = n42 & n280;
  assign n282 = n88 & n281;
  assign n283 = n91 & n281;
  assign n284 = n67 & n281;
  assign n285 = n59 & n281;
  assign n286 = n64 & n281;
  assign n287 = n100 & n281;
  assign n288 = v12 & n279;
  assign n289 = n69 & n288;
  assign n290 = n29 & n289;
  assign n291 = n51 & n281;
  assign n292 = n53 & n281;
  assign n293 = n48 & n281;
  assign n294 = ~n117 & n281;
  assign n295 = ~n169 & n260;
  assign n296 = ~n112 & n260;
  assign n297 = n29 & n280;
  assign n298 = n69 & n297;
  assign n299 = ~n172 & n260;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n27 & n281;
  assign n302 = ~n147 & n281;
  assign n303 = ~n301 & ~n302;
  assign n304 = n42 & n288;
  assign n305 = n53 & n304;
  assign n306 = n89 & n304;
  assign n307 = n88 & n304;
  assign n308 = n91 & n304;
  assign n309 = n102 & n281;
  assign n310 = n22 & n289;
  assign n311 = ~n149 & n304;
  assign n312 = ~n172 & n304;
  assign n313 = n139 & n258;
  assign n314 = ~n111 & n304;
  assign n315 = ~n313 & ~n314;
  assign n316 = ~n312 & n315;
  assign n317 = ~n47 & n316;
  assign n318 = ~n39 & n317;
  assign n319 = ~n146 & n318;
  assign n320 = ~n25 & n319;
  assign n321 = ~n50 & n320;
  assign n322 = n82 & n321;
  assign n323 = n56 & n320;
  assign n324 = n82 & n323;
  assign n325 = v7 & n316;
  assign n326 = ~n146 & n325;
  assign n327 = ~n25 & n326;
  assign n328 = ~n50 & n327;
  assign n329 = n82 & n328;
  assign n330 = n56 & n327;
  assign n331 = n82 & n330;
  assign n332 = ~n258 & n316;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n329 & n333;
  assign n335 = ~n324 & n334;
  assign n336 = ~n322 & n335;
  assign n337 = n64 & n258;
  assign n338 = n100 & n258;
  assign n339 = n130 & n280;
  assign n340 = n28 & n339;
  assign n341 = n21 & n339;
  assign n342 = n102 & n258;
  assign n343 = n40 & n339;
  assign n344 = n89 & n258;
  assign n345 = n88 & n258;
  assign n346 = n122 & n172;
  assign n347 = n116 & n346;
  assign n348 = n339 & ~n347;
  assign n349 = n83 & n258;
  assign n350 = n180 & ~n348;
  assign n351 = ~n345 & n350;
  assign n352 = ~n344 & n351;
  assign n353 = ~n343 & n352;
  assign n354 = ~n342 & n353;
  assign n355 = ~n341 & n354;
  assign n356 = ~n340 & n355;
  assign n357 = ~n338 & n356;
  assign n358 = ~n337 & n357;
  assign n359 = ~n146 & n358;
  assign n360 = ~n25 & n359;
  assign n361 = ~n336 & n360;
  assign n362 = ~n311 & n361;
  assign n363 = ~n310 & n362;
  assign n364 = ~n309 & n363;
  assign n365 = ~n308 & n364;
  assign n366 = ~n307 & n365;
  assign n367 = ~n306 & n366;
  assign n368 = ~n305 & n367;
  assign n369 = n303 & n368;
  assign n370 = n300 & n369;
  assign n371 = ~n296 & n370;
  assign n372 = ~n295 & n371;
  assign n373 = ~n294 & n372;
  assign n374 = ~n293 & n373;
  assign n375 = ~n292 & n374;
  assign n376 = ~n291 & n375;
  assign n377 = ~n290 & n376;
  assign n378 = ~n287 & n377;
  assign n379 = ~n286 & n378;
  assign n380 = ~n285 & n379;
  assign n381 = ~n284 & n380;
  assign n382 = ~n283 & n381;
  assign n383 = ~n282 & n382;
  assign n384 = ~n278 & n383;
  assign n385 = ~n277 & n384;
  assign n386 = ~n276 & n385;
  assign n387 = n275 & n386;
  assign n388 = ~n271 & n387;
  assign n389 = ~n267 & n388;
  assign n390 = ~n266 & n389;
  assign n391 = ~n265 & n390;
  assign n392 = ~n264 & n391;
  assign n393 = ~n263 & n392;
  assign n394 = ~n262 & n393;
  assign n395 = ~n261 & n394;
  assign n396 = ~n92 & n395;
  assign n397 = ~n259 & n396;
  assign n398 = ~n345 & ~n349;
  assign n399 = ~n344 & n398;
  assign n400 = ~n342 & n399;
  assign n401 = ~n338 & n400;
  assign n402 = ~n337 & n401;
  assign n403 = ~n336 & n402;
  assign n404 = ~n278 & n403;
  assign n405 = ~n277 & n404;
  assign n406 = ~n276 & n405;
  assign n407 = n275 & n406;
  assign n408 = ~n271 & n407;
  assign n409 = ~n267 & n408;
  assign n410 = ~n266 & n409;
  assign n411 = ~n265 & n410;
  assign n412 = ~n259 & n411;
  assign n413 = ~n339 & n412;
  assign n414 = ~n281 & n413;
  assign n415 = ~n260 & n414;
  assign n416 = ~n304 & n415;
  assign n417 = ~n397 & ~n416;
  assign n418 = n155 & n288;
  assign n419 = ~n117 & n418;
  assign n420 = n118 & n280;
  assign n421 = n40 & n420;
  assign n422 = n48 & n420;
  assign n423 = n51 & n420;
  assign n424 = n53 & n420;
  assign n425 = n104 & n280;
  assign n426 = n59 & n425;
  assign n427 = n64 & n425;
  assign n428 = ~n270 & n280;
  assign n429 = ~n25 & ~n139;
  assign n430 = n85 & n94;
  assign n431 = n149 & n430;
  assign n432 = n429 & n431;
  assign n433 = n425 & ~n432;
  assign n434 = n130 & n288;
  assign n435 = n91 & n434;
  assign n436 = n59 & n434;
  assign n437 = n64 & n434;
  assign n438 = n102 & n434;
  assign n439 = n51 & n434;
  assign n440 = n53 & n434;
  assign n441 = n48 & n434;
  assign n442 = ~n117 & n434;
  assign n443 = ~n172 & n420;
  assign n444 = n28 & n434;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n176 & n434;
  assign n447 = ~n83 & n111;
  assign n448 = n94 & n447;
  assign n449 = n420 & ~n448;
  assign n450 = n155 & n280;
  assign n451 = n40 & n450;
  assign n452 = n48 & n450;
  assign n453 = n51 & n450;
  assign n454 = n53 & n450;
  assign n455 = n32 & n155;
  assign n456 = n59 & n455;
  assign n457 = n64 & n455;
  assign n458 = n72 & n455;
  assign n459 = n139 & n450;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n432 & n455;
  assign n462 = n91 & n418;
  assign n463 = n59 & n418;
  assign n464 = n64 & n418;
  assign n465 = n104 & n288;
  assign n466 = n28 & n465;
  assign n467 = n51 & n418;
  assign n468 = n53 & n418;
  assign n469 = n48 & n418;
  assign n470 = n112 & n450;
  assign n471 = ~n102 & n470;
  assign n472 = n169 & n471;
  assign n473 = n114 & n472;
  assign n474 = n147 & ~n450;
  assign n475 = n429 & n474;
  assign n476 = ~n418 & ~n450;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n473 & n477;
  assign n479 = n67 & n455;
  assign n480 = ~n81 & ~n478;
  assign n481 = ~n80 & n480;
  assign n482 = ~n469 & n481;
  assign n483 = ~n468 & n482;
  assign n484 = ~n467 & n483;
  assign n485 = ~n466 & n484;
  assign n486 = ~n464 & n485;
  assign n487 = ~n463 & n486;
  assign n488 = ~n462 & n487;
  assign n489 = ~n461 & n488;
  assign n490 = n460 & n489;
  assign n491 = ~n457 & n490;
  assign n492 = ~n456 & n491;
  assign n493 = ~n454 & n492;
  assign n494 = ~n453 & n493;
  assign n495 = ~n452 & n494;
  assign n496 = ~n451 & n495;
  assign n497 = ~n449 & n496;
  assign n498 = ~n446 & n497;
  assign n499 = n445 & n498;
  assign n500 = ~n442 & n499;
  assign n501 = ~n441 & n500;
  assign n502 = ~n440 & n501;
  assign n503 = ~n439 & n502;
  assign n504 = ~n438 & n503;
  assign n505 = ~n437 & n504;
  assign n506 = ~n436 & n505;
  assign n507 = ~n435 & n506;
  assign n508 = ~n433 & n507;
  assign n509 = ~n428 & n508;
  assign n510 = ~n427 & n509;
  assign n511 = ~n426 & n510;
  assign n512 = ~n424 & n511;
  assign n513 = ~n423 & n512;
  assign n514 = ~n422 & n513;
  assign n515 = ~n421 & n514;
  assign n516 = ~n146 & n515;
  assign n517 = ~n25 & n516;
  assign n518 = ~n67 & n517;
  assign n519 = ~n92 & n518;
  assign n520 = ~n88 & n519;
  assign n521 = ~n419 & n520;
  assign n522 = ~n100 & n521;
  assign n523 = ~n461 & ~n466;
  assign n524 = n460 & n523;
  assign n525 = ~n479 & n524;
  assign n526 = ~n457 & n525;
  assign n527 = ~n456 & n526;
  assign n528 = ~n418 & n527;
  assign n529 = ~n450 & n528;
  assign n530 = ~n434 & n529;
  assign n531 = ~n425 & n530;
  assign n532 = ~n420 & n531;
  assign n533 = ~n522 & ~n532;
  assign n534 = v4 & n61;
  assign n535 = n25 & ~n26;
  assign n536 = v11 & n535;
  assign n537 = n288 & n536;
  assign n538 = n118 & n288;
  assign n539 = n146 & n538;
  assign n540 = n40 & n538;
  assign n541 = n48 & n538;
  assign n542 = n51 & n538;
  assign n543 = n53 & n538;
  assign n544 = n80 & n538;
  assign n545 = n81 & n538;
  assign n546 = n59 & n465;
  assign n547 = n64 & n465;
  assign n548 = n67 & n465;
  assign n549 = ~n270 & n288;
  assign n550 = ~n85 & n465;
  assign n551 = ~n94 & n465;
  assign n552 = ~n149 & n465;
  assign n553 = n102 & n418;
  assign n554 = n272 & n288;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n552 & n555;
  assign n557 = n31 & n279;
  assign n558 = v11 & n41;
  assign n559 = v8 & n30;
  assign n560 = ~n558 & ~n559;
  assign n561 = v12 & v15;
  assign n562 = n560 & ~n561;
  assign n563 = ~n557 & n562;
  assign n564 = n30 & ~n41;
  assign n565 = ~n30 & n41;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n31 & ~n279;
  assign n568 = n566 & ~n567;
  assign n569 = n37 & ~n62;
  assign n570 = n557 & n569;
  assign n571 = n18 & n56;
  assign n572 = ~n563 & n571;
  assign n573 = ~n568 & n569;
  assign n574 = ~n568 & n571;
  assign n575 = ~n448 & n538;
  assign n576 = ~n172 & n538;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~n574 & n577;
  assign n579 = ~n573 & n578;
  assign n580 = ~n572 & n579;
  assign n581 = ~n570 & n580;
  assign n582 = ~v6 & n37;
  assign n583 = v15 & ~n31;
  assign n584 = n560 & ~n583;
  assign n585 = ~v13 & ~v14;
  assign n586 = v3 & ~n56;
  assign n587 = ~v5 & n61;
  assign n588 = n557 & n587;
  assign n589 = ~n568 & n587;
  assign n590 = n582 & ~n584;
  assign n591 = n582 & n585;
  assign n592 = ~n566 & n582;
  assign n593 = n557 & n586;
  assign n594 = ~n568 & n586;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n592 & n595;
  assign n597 = ~n591 & n596;
  assign n598 = ~n590 & n597;
  assign n599 = ~n589 & n598;
  assign n600 = ~n588 & n599;
  assign n601 = v12 & ~v14;
  assign n602 = v0 & ~v2;
  assign n603 = ~n557 & ~n601;
  assign n604 = n602 & ~n603;
  assign n605 = ~v10 & n41;
  assign n606 = ~v9 & n30;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~v1 & v3;
  assign n609 = n279 & n607;
  assign n610 = ~n557 & n609;
  assign n611 = v13 & ~n534;
  assign n612 = n607 & n611;
  assign n613 = n31 & ~n279;
  assign n614 = n534 & n613;
  assign n615 = ~n534 & ~n608;
  assign n616 = ~n614 & ~n615;
  assign n617 = ~n612 & n616;
  assign n618 = ~n610 & n617;
  assign n619 = ~n584 & n602;
  assign n620 = ~v1 & n601;
  assign n621 = ~v2 & n620;
  assign n622 = n585 & n602;
  assign n623 = n602 & ~n607;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~n621 & n624;
  assign n626 = ~v1 & ~v2;
  assign n627 = ~n563 & n626;
  assign n628 = ~v13 & ~n279;
  assign n629 = n607 & ~n628;
  assign n630 = n626 & ~n629;
  assign n631 = n41 & n534;
  assign n632 = ~n627 & ~n630;
  assign n633 = n625 & n632;
  assign n634 = ~n619 & n633;
  assign n635 = ~n618 & n634;
  assign n636 = ~n604 & n635;
  assign n637 = n600 & n636;
  assign n638 = n581 & n637;
  assign n639 = n556 & n638;
  assign n640 = ~n551 & n639;
  assign n641 = ~n550 & n640;
  assign n642 = ~n549 & n641;
  assign n643 = ~n548 & n642;
  assign n644 = ~n547 & n643;
  assign n645 = ~n546 & n644;
  assign n646 = ~n545 & n645;
  assign n647 = ~n544 & n646;
  assign n648 = ~n543 & n647;
  assign n649 = ~n542 & n648;
  assign n650 = ~n541 & n649;
  assign n651 = ~n540 & n650;
  assign n652 = ~n539 & n651;
  assign n653 = ~n537 & n652;
  assign n654 = ~n534 & n653;
  assign n655 = ~v15 & ~n618;
  assign n656 = ~n30 & n655;
  assign n657 = n534 & n656;
  assign n658 = ~n631 & n657;
  assign n659 = ~n585 & n658;
  assign n660 = n30 & n655;
  assign n661 = n631 & n660;
  assign n662 = ~n585 & n661;
  assign n663 = v13 & ~n618;
  assign n664 = ~n30 & n663;
  assign n665 = n534 & n664;
  assign n666 = ~n631 & n665;
  assign n667 = n30 & n663;
  assign n668 = n631 & n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = ~n662 & n669;
  assign n671 = ~n659 & n670;
  assign n672 = ~n654 & n671;
  assign n673 = ~n533 & ~n672;
  assign n674 = ~n417 & n673;
  assign \v16.0  = n257 | ~n674;
endmodule


