// Benchmark "i6" written by ABC on Tue May 16 16:07:50 2017

module i6 ( 
    \V32(30) , \V138(3) , \V138(2) , \V138(4) , \V138(0) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(4) , \V32(5) , \V131(27) , \V32(6) ,
    \V131(26) , \V32(7) , \V131(29) , \V32(8) , \V131(28) , \V32(9) ,
    \V96(0) , \V96(1) , \V131(21) , \V96(2) , \V131(20) , \V96(3) ,
    \V131(23) , \V96(4) , \V96(13) , \V131(22) , \V96(5) , \V96(12) ,
    \V131(25) , \V96(6) , \V97(0) , \V96(15) , \V131(24) , \V96(7) ,
    \V96(14) , \V131(17) , \V96(8) , \V131(16) , \V96(9) , \V131(19) ,
    \V96(11) , \V131(18) , \V96(10) , \V98(0) , \V96(17) , \V96(16) ,
    \V131(11) , \V96(19) , \V131(10) , \V99(0) , \V96(18) , \V131(13) ,
    \V96(23) , \V131(12) , \V96(22) , \V131(15) , \V64(13) , \V96(25) ,
    \V131(14) , \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V96(21) ,
    \V96(20) , \V64(11) , \V64(10) , \V96(27) , \V96(26) , \V64(17) ,
    \V96(29) , \V64(16) , \V96(28) , \V131(3) , \V64(19) , \V131(2) ,
    \V64(18) , \V131(5) , \V64(23) , \V131(4) , \V64(22) , \V32(13) ,
    \V64(25) , \V32(12) , \V64(24) , \V32(15) , \V131(1) , \V32(14) ,
    \V96(31) , \V131(0) , \V96(30) , \V64(21) , \V64(20) , \V32(11) ,
    \V32(10) , \V131(7) , \V131(6) , \V131(9) , \V131(31) , \V64(27) ,
    \V131(8) , \V131(30) , \V64(26) , \V32(17) , \V64(29) , \V32(16) ,
    \V64(28) , \V32(19) , \V32(18) , \V133(1) , \V32(23) , \V133(0) ,
    \V64(0) , \V32(22) , \V64(1) , \V32(25) , \V64(2) , \V32(24) ,
    \V64(3) , \V64(4) , \V64(31) , \V64(5) , \V64(30) , \V32(21) ,
    \V64(6) , \V134(0) , \V32(20) , \V64(7) , \V64(8) , \V64(9) ,
    \V32(27) , \V32(26) , \V32(29) , \V32(28) , \V32(31) ,
    \V198(7) , \V198(6) , \V198(9) , \V198(8) , \V166(3) , \V166(2) ,
    \V166(5) , \V166(4) , \V166(1) , \V166(0) , \V166(7) , \V166(6) ,
    \V166(9) , \V198(27) , \V166(8) , \V205(3) , \V198(26) , \V205(2) ,
    \V198(29) , \V205(5) , \V198(28) , \V205(4) , \V205(1) , \V205(0) ,
    \V198(21) , \V198(20) , \V198(23) , \V198(22) , \V205(6) , \V198(25) ,
    \V198(24) , \V198(17) , \V198(16) , \V166(27) , \V198(19) , \V166(26) ,
    \V198(18) , \V198(11) , \V198(10) , \V166(21) , \V198(13) , \V166(20) ,
    \V198(12) , \V166(23) , \V198(15) , \V166(22) , \V198(14) , \V166(25) ,
    \V166(24) , \V166(17) , \V166(16) , \V166(19) , \V166(18) , \V166(11) ,
    \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) , \V198(3) ,
    \V198(2) , \V198(5) , \V198(4) , \V198(31) , \V198(30) , \V198(1) ,
    \V198(0)   );
  input  \V32(30) , \V138(3) , \V138(2) , \V138(4) , \V138(0) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(4) , \V32(5) , \V131(27) , \V32(6) ,
    \V131(26) , \V32(7) , \V131(29) , \V32(8) , \V131(28) , \V32(9) ,
    \V96(0) , \V96(1) , \V131(21) , \V96(2) , \V131(20) , \V96(3) ,
    \V131(23) , \V96(4) , \V96(13) , \V131(22) , \V96(5) , \V96(12) ,
    \V131(25) , \V96(6) , \V97(0) , \V96(15) , \V131(24) , \V96(7) ,
    \V96(14) , \V131(17) , \V96(8) , \V131(16) , \V96(9) , \V131(19) ,
    \V96(11) , \V131(18) , \V96(10) , \V98(0) , \V96(17) , \V96(16) ,
    \V131(11) , \V96(19) , \V131(10) , \V99(0) , \V96(18) , \V131(13) ,
    \V96(23) , \V131(12) , \V96(22) , \V131(15) , \V64(13) , \V96(25) ,
    \V131(14) , \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V96(21) ,
    \V96(20) , \V64(11) , \V64(10) , \V96(27) , \V96(26) , \V64(17) ,
    \V96(29) , \V64(16) , \V96(28) , \V131(3) , \V64(19) , \V131(2) ,
    \V64(18) , \V131(5) , \V64(23) , \V131(4) , \V64(22) , \V32(13) ,
    \V64(25) , \V32(12) , \V64(24) , \V32(15) , \V131(1) , \V32(14) ,
    \V96(31) , \V131(0) , \V96(30) , \V64(21) , \V64(20) , \V32(11) ,
    \V32(10) , \V131(7) , \V131(6) , \V131(9) , \V131(31) , \V64(27) ,
    \V131(8) , \V131(30) , \V64(26) , \V32(17) , \V64(29) , \V32(16) ,
    \V64(28) , \V32(19) , \V32(18) , \V133(1) , \V32(23) , \V133(0) ,
    \V64(0) , \V32(22) , \V64(1) , \V32(25) , \V64(2) , \V32(24) ,
    \V64(3) , \V64(4) , \V64(31) , \V64(5) , \V64(30) , \V32(21) ,
    \V64(6) , \V134(0) , \V32(20) , \V64(7) , \V64(8) , \V64(9) ,
    \V32(27) , \V32(26) , \V32(29) , \V32(28) , \V32(31) ;
  output \V198(7) , \V198(6) , \V198(9) , \V198(8) , \V166(3) , \V166(2) ,
    \V166(5) , \V166(4) , \V166(1) , \V166(0) , \V166(7) , \V166(6) ,
    \V166(9) , \V198(27) , \V166(8) , \V205(3) , \V198(26) , \V205(2) ,
    \V198(29) , \V205(5) , \V198(28) , \V205(4) , \V205(1) , \V205(0) ,
    \V198(21) , \V198(20) , \V198(23) , \V198(22) , \V205(6) , \V198(25) ,
    \V198(24) , \V198(17) , \V198(16) , \V166(27) , \V198(19) , \V166(26) ,
    \V198(18) , \V198(11) , \V198(10) , \V166(21) , \V198(13) , \V166(20) ,
    \V198(12) , \V166(23) , \V198(15) , \V166(22) , \V198(14) , \V166(25) ,
    \V166(24) , \V166(17) , \V166(16) , \V166(19) , \V166(18) , \V166(11) ,
    \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) , \V198(3) ,
    \V198(2) , \V198(5) , \V198(4) , \V198(31) , \V198(30) , \V198(1) ,
    \V198(0) ;
  wire n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n219, n220, n221, n222, n223, n225, n226, n227, n228, n229, n231,
    n232, n233, n234, n235, n237, n238, n239, n240, n242, n243, n244, n245,
    n247, n248, n249, n250, n252, n253, n254, n255, n257, n258, n259, n260,
    n262, n263, n264, n265, n267, n268, n269, n270, n272, n273, n274, n275,
    n277, n278, n279, n280, n282, n283, n284, n285, n286, n288, n289, n290,
    n291, n293, n294, n295, n296, n297, n298, n299, n300, n301, n303, n304,
    n305, n306, n307, n309, n310, n311, n312, n313, n315, n316, n317, n318,
    n319, n321, n322, n323, n324, n325, n327, n328, n329, n330, n331, n333,
    n334, n335, n336, n337, n339, n340, n341, n342, n343, n345, n346, n347,
    n348, n349, n351, n352, n353, n354, n355, n357, n358, n359, n360, n361,
    n363, n364, n365, n366, n367, n369, n370, n371, n372, n373, n375, n376,
    n377, n378, n379, n380, n381, n383, n384, n385, n386, n387, n389, n390,
    n391, n392, n393, n395, n396, n397, n398, n399, n401, n402, n403, n404,
    n405, n407, n408, n409, n410, n412, n413, n414, n415, n416, n418, n419,
    n420, n421, n423, n424, n425, n426, n427, n429, n430, n431, n432, n433,
    n435, n436, n437, n438, n439, n441, n442, n443, n444, n446, n447, n448,
    n449, n450, n452, n453, n454, n455, n457, n458, n459, n460, n461, n463,
    n464, n465, n466, n468, n469, n470, n471, n472, n474, n475, n476, n477,
    n479, n480, n481, n482, n483, n485, n486, n487, n488, n490, n491, n492,
    n493, n495, n496, n497, n498, n500, n501, n502, n503, n505, n506, n507,
    n508, n510, n511, n512, n513, n515, n516, n517, n518, n520, n521, n522,
    n523, n525, n526, n527, n528, n530, n531, n532, n533, n535, n536, n537,
    n538, n540, n541, n542, n543, n545, n546, n547, n548, n549, n551, n552,
    n553, n554, n555, n557, n558, n559, n560, n561, n563, n564, n565, n566,
    n567, n569, n570, n571, n572, n573, n574, n576, n577, n578, n579, n580,
    n582, n583, n584, n585, n586, n588, n589, n590, n591, n592;
  assign n206 = \V138(2)  & ~\V138(4) ;
  assign n207 = \V138(2)  & \V138(0) ;
  assign n208 = \V138(4)  & n207;
  assign n209 = ~\V131(3)  & n208;
  assign n210 = ~\V138(2)  & \V138(0) ;
  assign n211 = \V138(4)  & n210;
  assign n212 = \V131(3)  & n211;
  assign n213 = ~\V138(2)  & ~\V138(0) ;
  assign n214 = \V138(4)  & n213;
  assign n215 = \V96(3)  & n214;
  assign n216 = ~n212 & ~n215;
  assign n217 = ~n209 & n216;
  assign \V198(7)  = n206 | ~n217;
  assign n219 = ~\V131(2)  & n208;
  assign n220 = \V131(2)  & n211;
  assign n221 = \V96(2)  & n214;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~n219 & n222;
  assign \V198(6)  = n206 | ~n223;
  assign n225 = ~\V131(5)  & n208;
  assign n226 = \V131(5)  & n211;
  assign n227 = \V96(5)  & n214;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n225 & n228;
  assign \V198(9)  = n206 | ~n229;
  assign n231 = ~\V131(4)  & n208;
  assign n232 = \V131(4)  & n211;
  assign n233 = \V96(4)  & n214;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n231 & n234;
  assign \V198(8)  = n206 | ~n235;
  assign n237 = ~\V64(3)  & n207;
  assign n238 = \V64(3)  & n210;
  assign n239 = \V32(3)  & n213;
  assign n240 = ~n238 & ~n239;
  assign \V166(3)  = n237 | ~n240;
  assign n242 = ~\V64(2)  & n207;
  assign n243 = \V64(2)  & n210;
  assign n244 = \V32(2)  & n213;
  assign n245 = ~n243 & ~n244;
  assign \V166(2)  = n242 | ~n245;
  assign n247 = ~\V64(5)  & n207;
  assign n248 = \V64(5)  & n210;
  assign n249 = \V32(5)  & n213;
  assign n250 = ~n248 & ~n249;
  assign \V166(5)  = n247 | ~n250;
  assign n252 = ~\V64(4)  & n207;
  assign n253 = \V64(4)  & n210;
  assign n254 = \V32(4)  & n213;
  assign n255 = ~n253 & ~n254;
  assign \V166(4)  = n252 | ~n255;
  assign n257 = ~\V64(1)  & n207;
  assign n258 = \V64(1)  & n210;
  assign n259 = \V32(1)  & n213;
  assign n260 = ~n258 & ~n259;
  assign \V166(1)  = n257 | ~n260;
  assign n262 = ~\V64(0)  & n207;
  assign n263 = \V64(0)  & n210;
  assign n264 = \V32(0)  & n213;
  assign n265 = ~n263 & ~n264;
  assign \V166(0)  = n262 | ~n265;
  assign n267 = ~\V64(7)  & n207;
  assign n268 = \V64(7)  & n210;
  assign n269 = \V32(7)  & n213;
  assign n270 = ~n268 & ~n269;
  assign \V166(7)  = n267 | ~n270;
  assign n272 = ~\V64(6)  & n207;
  assign n273 = \V64(6)  & n210;
  assign n274 = \V32(6)  & n213;
  assign n275 = ~n273 & ~n274;
  assign \V166(6)  = n272 | ~n275;
  assign n277 = ~\V64(9)  & n207;
  assign n278 = \V64(9)  & n210;
  assign n279 = \V32(9)  & n213;
  assign n280 = ~n278 & ~n279;
  assign \V166(9)  = n277 | ~n280;
  assign n282 = ~\V131(23)  & n208;
  assign n283 = \V131(23)  & n211;
  assign n284 = \V96(23)  & n214;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n282 & n285;
  assign \V198(27)  = n206 | ~n286;
  assign n288 = ~\V64(8)  & n207;
  assign n289 = \V64(8)  & n210;
  assign n290 = \V32(8)  & n213;
  assign n291 = ~n289 & ~n290;
  assign \V166(8)  = n288 | ~n291;
  assign n293 = ~\V138(3)  & \V138(2) ;
  assign n294 = \V138(3)  & n207;
  assign n295 = ~\V131(31)  & n294;
  assign n296 = \V138(3)  & n210;
  assign n297 = \V131(31)  & n296;
  assign n298 = \V138(3)  & n213;
  assign n299 = \V96(31)  & n298;
  assign n300 = ~n297 & ~n299;
  assign n301 = ~n295 & n300;
  assign \V205(3)  = n293 | ~n301;
  assign n303 = ~\V131(22)  & n208;
  assign n304 = \V131(22)  & n211;
  assign n305 = \V96(22)  & n214;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & n306;
  assign \V198(26)  = n206 | ~n307;
  assign n309 = ~\V131(30)  & n294;
  assign n310 = \V131(30)  & n296;
  assign n311 = \V96(30)  & n298;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~n309 & n312;
  assign \V205(2)  = n293 | ~n313;
  assign n315 = ~\V131(25)  & n208;
  assign n316 = \V131(25)  & n211;
  assign n317 = \V96(25)  & n214;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n315 & n318;
  assign \V198(29)  = n206 | ~n319;
  assign n321 = ~\V133(1)  & n294;
  assign n322 = \V133(1)  & n296;
  assign n323 = \V98(0)  & n298;
  assign n324 = ~n322 & ~n323;
  assign n325 = ~n321 & n324;
  assign \V205(5)  = n293 | ~n325;
  assign n327 = ~\V131(24)  & n208;
  assign n328 = \V131(24)  & n211;
  assign n329 = \V96(24)  & n214;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~n327 & n330;
  assign \V198(28)  = n206 | ~n331;
  assign n333 = ~\V133(0)  & n294;
  assign n334 = \V133(0)  & n296;
  assign n335 = \V97(0)  & n298;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~n333 & n336;
  assign \V205(4)  = n293 | ~n337;
  assign n339 = ~\V131(29)  & n294;
  assign n340 = \V131(29)  & n296;
  assign n341 = \V96(29)  & n298;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~n339 & n342;
  assign \V205(1)  = n293 | ~n343;
  assign n345 = ~\V131(28)  & n294;
  assign n346 = \V131(28)  & n296;
  assign n347 = \V96(28)  & n298;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n345 & n348;
  assign \V205(0)  = n293 | ~n349;
  assign n351 = ~\V131(17)  & n208;
  assign n352 = \V131(17)  & n211;
  assign n353 = \V96(17)  & n214;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n351 & n354;
  assign \V198(21)  = n206 | ~n355;
  assign n357 = ~\V131(16)  & n208;
  assign n358 = \V131(16)  & n211;
  assign n359 = \V96(16)  & n214;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign \V198(20)  = n206 | ~n361;
  assign n363 = ~\V131(19)  & n208;
  assign n364 = \V131(19)  & n211;
  assign n365 = \V96(19)  & n214;
  assign n366 = ~n364 & ~n365;
  assign n367 = ~n363 & n366;
  assign \V198(23)  = n206 | ~n367;
  assign n369 = ~\V131(18)  & n208;
  assign n370 = \V131(18)  & n211;
  assign n371 = \V96(18)  & n214;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n369 & n372;
  assign \V198(22)  = n206 | ~n373;
  assign n375 = \V138(0)  & \V134(0) ;
  assign n376 = \V138(2)  & n375;
  assign n377 = \V138(3)  & n376;
  assign n378 = \V134(0)  & n296;
  assign n379 = \V99(0)  & n213;
  assign n380 = \V138(3)  & n379;
  assign n381 = ~n378 & ~n380;
  assign \V205(6)  = n377 | ~n381;
  assign n383 = ~\V131(21)  & n208;
  assign n384 = \V131(21)  & n211;
  assign n385 = \V96(21)  & n214;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n383 & n386;
  assign \V198(25)  = n206 | ~n387;
  assign n389 = ~\V131(20)  & n208;
  assign n390 = \V131(20)  & n211;
  assign n391 = \V96(20)  & n214;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n389 & n392;
  assign \V198(24)  = n206 | ~n393;
  assign n395 = ~\V131(13)  & n208;
  assign n396 = \V131(13)  & n211;
  assign n397 = \V96(13)  & n214;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n395 & n398;
  assign \V198(17)  = n206 | ~n399;
  assign n401 = ~\V131(12)  & n208;
  assign n402 = \V131(12)  & n211;
  assign n403 = \V96(12)  & n214;
  assign n404 = ~n402 & ~n403;
  assign n405 = ~n401 & n404;
  assign \V198(16)  = n206 | ~n405;
  assign n407 = ~\V64(27)  & n207;
  assign n408 = \V64(27)  & n210;
  assign n409 = \V32(27)  & n213;
  assign n410 = ~n408 & ~n409;
  assign \V166(27)  = n407 | ~n410;
  assign n412 = ~\V131(15)  & n208;
  assign n413 = \V131(15)  & n211;
  assign n414 = \V96(15)  & n214;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~n412 & n415;
  assign \V198(19)  = n206 | ~n416;
  assign n418 = ~\V64(26)  & n207;
  assign n419 = \V64(26)  & n210;
  assign n420 = \V32(26)  & n213;
  assign n421 = ~n419 & ~n420;
  assign \V166(26)  = n418 | ~n421;
  assign n423 = ~\V131(14)  & n208;
  assign n424 = \V131(14)  & n211;
  assign n425 = \V96(14)  & n214;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n423 & n426;
  assign \V198(18)  = n206 | ~n427;
  assign n429 = ~\V131(7)  & n208;
  assign n430 = \V131(7)  & n211;
  assign n431 = \V96(7)  & n214;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~n429 & n432;
  assign \V198(11)  = n206 | ~n433;
  assign n435 = ~\V131(6)  & n208;
  assign n436 = \V131(6)  & n211;
  assign n437 = \V96(6)  & n214;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n435 & n438;
  assign \V198(10)  = n206 | ~n439;
  assign n441 = ~\V64(21)  & n207;
  assign n442 = \V64(21)  & n210;
  assign n443 = \V32(21)  & n213;
  assign n444 = ~n442 & ~n443;
  assign \V166(21)  = n441 | ~n444;
  assign n446 = ~\V131(9)  & n208;
  assign n447 = \V131(9)  & n211;
  assign n448 = \V96(9)  & n214;
  assign n449 = ~n447 & ~n448;
  assign n450 = ~n446 & n449;
  assign \V198(13)  = n206 | ~n450;
  assign n452 = ~\V64(20)  & n207;
  assign n453 = \V64(20)  & n210;
  assign n454 = \V32(20)  & n213;
  assign n455 = ~n453 & ~n454;
  assign \V166(20)  = n452 | ~n455;
  assign n457 = ~\V131(8)  & n208;
  assign n458 = \V131(8)  & n211;
  assign n459 = \V96(8)  & n214;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n457 & n460;
  assign \V198(12)  = n206 | ~n461;
  assign n463 = ~\V64(23)  & n207;
  assign n464 = \V64(23)  & n210;
  assign n465 = \V32(23)  & n213;
  assign n466 = ~n464 & ~n465;
  assign \V166(23)  = n463 | ~n466;
  assign n468 = ~\V131(11)  & n208;
  assign n469 = \V131(11)  & n211;
  assign n470 = \V96(11)  & n214;
  assign n471 = ~n469 & ~n470;
  assign n472 = ~n468 & n471;
  assign \V198(15)  = n206 | ~n472;
  assign n474 = ~\V64(22)  & n207;
  assign n475 = \V64(22)  & n210;
  assign n476 = \V32(22)  & n213;
  assign n477 = ~n475 & ~n476;
  assign \V166(22)  = n474 | ~n477;
  assign n479 = ~\V131(10)  & n208;
  assign n480 = \V131(10)  & n211;
  assign n481 = \V96(10)  & n214;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n479 & n482;
  assign \V198(14)  = n206 | ~n483;
  assign n485 = ~\V64(25)  & n207;
  assign n486 = \V64(25)  & n210;
  assign n487 = \V32(25)  & n213;
  assign n488 = ~n486 & ~n487;
  assign \V166(25)  = n485 | ~n488;
  assign n490 = ~\V64(24)  & n207;
  assign n491 = \V64(24)  & n210;
  assign n492 = \V32(24)  & n213;
  assign n493 = ~n491 & ~n492;
  assign \V166(24)  = n490 | ~n493;
  assign n495 = ~\V64(17)  & n207;
  assign n496 = \V64(17)  & n210;
  assign n497 = \V32(17)  & n213;
  assign n498 = ~n496 & ~n497;
  assign \V166(17)  = n495 | ~n498;
  assign n500 = ~\V64(16)  & n207;
  assign n501 = \V64(16)  & n210;
  assign n502 = \V32(16)  & n213;
  assign n503 = ~n501 & ~n502;
  assign \V166(16)  = n500 | ~n503;
  assign n505 = ~\V64(19)  & n207;
  assign n506 = \V64(19)  & n210;
  assign n507 = \V32(19)  & n213;
  assign n508 = ~n506 & ~n507;
  assign \V166(19)  = n505 | ~n508;
  assign n510 = ~\V64(18)  & n207;
  assign n511 = \V64(18)  & n210;
  assign n512 = \V32(18)  & n213;
  assign n513 = ~n511 & ~n512;
  assign \V166(18)  = n510 | ~n513;
  assign n515 = ~\V64(11)  & n207;
  assign n516 = \V64(11)  & n210;
  assign n517 = \V32(11)  & n213;
  assign n518 = ~n516 & ~n517;
  assign \V166(11)  = n515 | ~n518;
  assign n520 = ~\V64(10)  & n207;
  assign n521 = \V64(10)  & n210;
  assign n522 = \V32(10)  & n213;
  assign n523 = ~n521 & ~n522;
  assign \V166(10)  = n520 | ~n523;
  assign n525 = ~\V64(13)  & n207;
  assign n526 = \V64(13)  & n210;
  assign n527 = \V32(13)  & n213;
  assign n528 = ~n526 & ~n527;
  assign \V166(13)  = n525 | ~n528;
  assign n530 = ~\V64(12)  & n207;
  assign n531 = \V64(12)  & n210;
  assign n532 = \V32(12)  & n213;
  assign n533 = ~n531 & ~n532;
  assign \V166(12)  = n530 | ~n533;
  assign n535 = ~\V64(15)  & n207;
  assign n536 = \V64(15)  & n210;
  assign n537 = \V32(15)  & n213;
  assign n538 = ~n536 & ~n537;
  assign \V166(15)  = n535 | ~n538;
  assign n540 = ~\V64(14)  & n207;
  assign n541 = \V64(14)  & n210;
  assign n542 = \V32(14)  & n213;
  assign n543 = ~n541 & ~n542;
  assign \V166(14)  = n540 | ~n543;
  assign n545 = ~\V64(31)  & n208;
  assign n546 = \V64(31)  & n211;
  assign n547 = \V32(31)  & n214;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n545 & n548;
  assign \V198(3)  = n206 | ~n549;
  assign n551 = ~\V64(30)  & n208;
  assign n552 = \V64(30)  & n211;
  assign n553 = \V32(30)  & n214;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~n551 & n554;
  assign \V198(2)  = n206 | ~n555;
  assign n557 = ~\V131(1)  & n208;
  assign n558 = \V131(1)  & n211;
  assign n559 = \V96(1)  & n214;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n557 & n560;
  assign \V198(5)  = n206 | ~n561;
  assign n563 = ~\V131(0)  & n208;
  assign n564 = \V131(0)  & n211;
  assign n565 = \V96(0)  & n214;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n563 & n566;
  assign \V198(4)  = n206 | ~n567;
  assign n569 = ~\V131(27)  & n208;
  assign n570 = \V131(27)  & n211;
  assign n571 = \V96(27)  & n213;
  assign n572 = \V138(4)  & n571;
  assign n573 = ~n570 & ~n572;
  assign n574 = ~n569 & n573;
  assign \V198(31)  = n206 | ~n574;
  assign n576 = ~\V131(26)  & n208;
  assign n577 = \V131(26)  & n211;
  assign n578 = \V96(26)  & n214;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n576 & n579;
  assign \V198(30)  = n206 | ~n580;
  assign n582 = ~\V64(29)  & n208;
  assign n583 = \V64(29)  & n211;
  assign n584 = \V32(29)  & n214;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n582 & n585;
  assign \V198(1)  = n206 | ~n586;
  assign n588 = ~\V64(28)  & n208;
  assign n589 = \V64(28)  & n211;
  assign n590 = \V32(28)  & n214;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n588 & n591;
  assign \V198(0)  = n206 | ~n592;
endmodule


