// Benchmark "i4" written by ABC on Tue May 16 16:07:50 2017

module i4 ( 
    \V186(2) , \V88(11) , \V88(10) , \V186(1) , \V144(10) , \V186(0) ,
    \V144(13) , \V88(17) , \V144(12) , \V88(16) , \V88(19) , \V144(14) ,
    \V180(10) , \V88(18) , \V180(13) , \V88(23) , \V126(3) , \V180(12) ,
    \V56(0) , \V88(22) , \V126(2) , \V56(13) , \V56(1) , \V88(25) ,
    \V126(5) , \V56(12) , \V180(14) , \V56(2) , \V88(24) , \V126(4) ,
    \V56(15) , \V56(3) , \V56(14) , \V56(4) , \V56(5) , \V88(21) ,
    \V126(1) , \V56(6) , \V88(20) , \V126(0) , \V56(11) , \V56(7) ,
    \V189(2) , \V56(10) , \V56(8) , \V56(9) , \V88(27) , \V88(26) ,
    \V189(1) , \V56(17) , \V88(29) , \V189(0) , \V56(16) , \V88(28) ,
    \V56(19) , \V56(18) , \V56(23) , \V56(22) , \V56(25) , \V56(24) ,
    \V88(31) , \V88(30) , \V56(21) , \V56(20) , \V56(27) , \V56(26) ,
    \V120(27) , \V120(26) , \V120(29) , \V120(28) , \V168(10) , \V168(2) ,
    \V168(13) , \V168(5) , \V168(12) , \V168(4) , \V120(21) , \V120(20) ,
    \V168(14) , \V120(23) , \V28(13) , \V168(1) , \V120(22) , \V28(12) ,
    \V168(0) , \V120(25) , \V28(15) , \V120(24) , \V28(14) , \V120(17) ,
    \V120(16) , \V156(2) , \V120(19) , \V28(11) , \V156(5) , \V120(18) ,
    \V28(10) , \V168(6) , \V156(4) , \V168(9) , \V168(8) , \V156(1) ,
    \V156(0) , \V28(17) , \V28(16) , \V192(2) , \V120(11) , \V28(19) ,
    \V120(10) , \V28(18) , \V144(2) , \V120(13) , \V28(23) , \V144(5) ,
    \V120(12) , \V28(22) , \V156(6) , \V144(4) , \V120(15) , \V88(0) ,
    \V28(25) , \V156(9) , \V192(1) , \V120(14) , \V88(1) , \V28(24) ,
    \V156(8) , \V192(0) , \V88(2) , \V144(1) , \V88(3) , \V144(0) ,
    \V88(4) , \V28(21) , \V88(5) , \V28(20) , \V180(2) , \V88(6) ,
    \V132(3) , \V180(5) , \V88(7) , \V132(2) , \V180(4) , \V88(8) ,
    \V132(5) , \V88(9) , \V144(6) , \V132(4) , \V28(27) , \V144(9) ,
    \V180(1) , \V28(26) , \V144(8) , \V180(0) , \V28(0) , \V132(1) ,
    \V156(10) , \V28(1) , \V132(0) , \V156(13) , \V28(2) , \V156(12) ,
    \V28(3) , \V28(4) , \V120(3) , \V156(14) , \V28(5) , \V180(6) ,
    \V120(2) , \V28(6) , \V180(9) , \V120(5) , \V28(7) , \V180(8) ,
    \V120(4) , \V28(8) , \V28(9) , \V120(1) , \V120(0) , \V183(2) ,
    \V120(31) , \V120(7) , \V120(30) , \V120(6) , \V183(1) , \V120(9) ,
    \V183(0) , \V120(8) , \V88(13) , \V88(12) , \V88(15) , \V88(14) ,
    \V194(1) , \V194(0) , \V198(3) , \V198(2) , \V198(1) , \V198(0)   );
  input  \V186(2) , \V88(11) , \V88(10) , \V186(1) , \V144(10) ,
    \V186(0) , \V144(13) , \V88(17) , \V144(12) , \V88(16) , \V88(19) ,
    \V144(14) , \V180(10) , \V88(18) , \V180(13) , \V88(23) , \V126(3) ,
    \V180(12) , \V56(0) , \V88(22) , \V126(2) , \V56(13) , \V56(1) ,
    \V88(25) , \V126(5) , \V56(12) , \V180(14) , \V56(2) , \V88(24) ,
    \V126(4) , \V56(15) , \V56(3) , \V56(14) , \V56(4) , \V56(5) ,
    \V88(21) , \V126(1) , \V56(6) , \V88(20) , \V126(0) , \V56(11) ,
    \V56(7) , \V189(2) , \V56(10) , \V56(8) , \V56(9) , \V88(27) ,
    \V88(26) , \V189(1) , \V56(17) , \V88(29) , \V189(0) , \V56(16) ,
    \V88(28) , \V56(19) , \V56(18) , \V56(23) , \V56(22) , \V56(25) ,
    \V56(24) , \V88(31) , \V88(30) , \V56(21) , \V56(20) , \V56(27) ,
    \V56(26) , \V120(27) , \V120(26) , \V120(29) , \V120(28) , \V168(10) ,
    \V168(2) , \V168(13) , \V168(5) , \V168(12) , \V168(4) , \V120(21) ,
    \V120(20) , \V168(14) , \V120(23) , \V28(13) , \V168(1) , \V120(22) ,
    \V28(12) , \V168(0) , \V120(25) , \V28(15) , \V120(24) , \V28(14) ,
    \V120(17) , \V120(16) , \V156(2) , \V120(19) , \V28(11) , \V156(5) ,
    \V120(18) , \V28(10) , \V168(6) , \V156(4) , \V168(9) , \V168(8) ,
    \V156(1) , \V156(0) , \V28(17) , \V28(16) , \V192(2) , \V120(11) ,
    \V28(19) , \V120(10) , \V28(18) , \V144(2) , \V120(13) , \V28(23) ,
    \V144(5) , \V120(12) , \V28(22) , \V156(6) , \V144(4) , \V120(15) ,
    \V88(0) , \V28(25) , \V156(9) , \V192(1) , \V120(14) , \V88(1) ,
    \V28(24) , \V156(8) , \V192(0) , \V88(2) , \V144(1) , \V88(3) ,
    \V144(0) , \V88(4) , \V28(21) , \V88(5) , \V28(20) , \V180(2) ,
    \V88(6) , \V132(3) , \V180(5) , \V88(7) , \V132(2) , \V180(4) ,
    \V88(8) , \V132(5) , \V88(9) , \V144(6) , \V132(4) , \V28(27) ,
    \V144(9) , \V180(1) , \V28(26) , \V144(8) , \V180(0) , \V28(0) ,
    \V132(1) , \V156(10) , \V28(1) , \V132(0) , \V156(13) , \V28(2) ,
    \V156(12) , \V28(3) , \V28(4) , \V120(3) , \V156(14) , \V28(5) ,
    \V180(6) , \V120(2) , \V28(6) , \V180(9) , \V120(5) , \V28(7) ,
    \V180(8) , \V120(4) , \V28(8) , \V28(9) , \V120(1) , \V120(0) ,
    \V183(2) , \V120(31) , \V120(7) , \V120(30) , \V120(6) , \V183(1) ,
    \V120(9) , \V183(0) , \V120(8) , \V88(13) , \V88(12) , \V88(15) ,
    \V88(14) ;
  output \V194(1) , \V194(0) , \V198(3) , \V198(2) , \V198(1) , \V198(0) ;
  wire n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443;
  assign \V194(1)  = \V56(1)  & \V28(1) ;
  assign \V194(0)  = \V56(0)  & \V28(0) ;
  assign n201 = \V132(0)  & \V180(9) ;
  assign n202 = \V126(0)  & n201;
  assign n203 = \V180(8)  & n202;
  assign n204 = \V88(30)  & \V120(30) ;
  assign n205 = \V88(31)  & \V180(8) ;
  assign n206 = \V120(31)  & n205;
  assign n207 = \V180(10)  & \V180(8) ;
  assign n208 = \V126(1)  & n207;
  assign n209 = \V132(1)  & n208;
  assign n210 = \V180(9)  & n209;
  assign n211 = ~n206 & ~n210;
  assign n212 = ~n204 & n211;
  assign n213 = ~n203 & n212;
  assign n214 = \V192(1)  & ~n213;
  assign n215 = \V192(0)  & n214;
  assign n216 = \V180(2)  & \V180(0) ;
  assign n217 = \V88(25)  & n216;
  assign n218 = \V120(25)  & n217;
  assign n219 = \V180(1)  & n218;
  assign n220 = \V88(23)  & \V180(0) ;
  assign n221 = \V120(23)  & n220;
  assign n222 = \V88(22)  & \V120(22) ;
  assign n223 = \V120(24)  & \V180(1) ;
  assign n224 = \V88(24)  & n223;
  assign n225 = \V180(0)  & n224;
  assign n226 = \V120(28)  & \V180(5) ;
  assign n227 = \V88(28)  & n226;
  assign n228 = \V180(4)  & n227;
  assign n229 = \V88(26)  & \V120(26) ;
  assign n230 = \V88(27)  & \V180(4) ;
  assign n231 = \V120(27)  & n230;
  assign n232 = \V180(4)  & \V180(6) ;
  assign n233 = \V88(29)  & n232;
  assign n234 = \V120(29)  & n233;
  assign n235 = \V180(5)  & n234;
  assign n236 = ~n231 & ~n235;
  assign n237 = ~n229 & n236;
  assign n238 = ~n228 & n237;
  assign n239 = \V192(0)  & ~n238;
  assign n240 = \V180(13)  & \V132(4) ;
  assign n241 = \V126(4)  & n240;
  assign n242 = \V180(12)  & n241;
  assign n243 = \V126(2)  & \V132(2) ;
  assign n244 = \V126(3)  & \V180(12) ;
  assign n245 = \V132(3)  & n244;
  assign n246 = \V180(12)  & \V180(14) ;
  assign n247 = \V126(5)  & n246;
  assign n248 = \V132(5)  & n247;
  assign n249 = \V180(13)  & n248;
  assign n250 = ~n245 & ~n249;
  assign n251 = ~n243 & n250;
  assign n252 = ~n242 & n251;
  assign n253 = \V192(2)  & \V192(0) ;
  assign n254 = ~n252 & n253;
  assign n255 = \V192(1)  & n254;
  assign n256 = ~n239 & ~n255;
  assign n257 = ~n225 & n256;
  assign n258 = ~n222 & n257;
  assign n259 = ~n221 & n258;
  assign n260 = ~n219 & n259;
  assign \V198(3)  = n215 | ~n260;
  assign n262 = \V120(16)  & \V168(9) ;
  assign n263 = \V88(16)  & n262;
  assign n264 = \V168(8)  & n263;
  assign n265 = \V120(14)  & \V88(14) ;
  assign n266 = \V168(8)  & \V88(15) ;
  assign n267 = \V120(15)  & n266;
  assign n268 = \V168(10)  & \V168(8) ;
  assign n269 = \V88(17)  & n268;
  assign n270 = \V120(17)  & n269;
  assign n271 = \V168(9)  & n270;
  assign n272 = ~n267 & ~n271;
  assign n273 = ~n265 & n272;
  assign n274 = ~n264 & n273;
  assign n275 = \V189(1)  & ~n274;
  assign n276 = \V189(0)  & n275;
  assign n277 = \V168(2)  & \V168(0) ;
  assign n278 = \V88(9)  & n277;
  assign n279 = \V120(9)  & n278;
  assign n280 = \V168(1)  & n279;
  assign n281 = \V168(0)  & \V88(7) ;
  assign n282 = \V120(7)  & n281;
  assign n283 = \V88(6)  & \V120(6) ;
  assign n284 = \V168(1)  & \V120(8) ;
  assign n285 = \V88(8)  & n284;
  assign n286 = \V168(0)  & n285;
  assign n287 = \V168(5)  & \V120(12) ;
  assign n288 = \V88(12)  & n287;
  assign n289 = \V168(4)  & n288;
  assign n290 = \V88(10)  & \V120(10) ;
  assign n291 = \V88(11)  & \V168(4) ;
  assign n292 = \V120(11)  & n291;
  assign n293 = \V168(4)  & \V168(6) ;
  assign n294 = \V88(13)  & n293;
  assign n295 = \V120(13)  & n294;
  assign n296 = \V168(5)  & n295;
  assign n297 = ~n292 & ~n296;
  assign n298 = ~n290 & n297;
  assign n299 = ~n289 & n298;
  assign n300 = \V189(0)  & ~n299;
  assign n301 = \V168(13)  & \V120(20) ;
  assign n302 = \V88(20)  & n301;
  assign n303 = \V168(12)  & n302;
  assign n304 = \V88(18)  & \V120(18) ;
  assign n305 = \V88(19)  & \V168(12) ;
  assign n306 = \V120(19)  & n305;
  assign n307 = \V168(12)  & \V168(14) ;
  assign n308 = \V88(21)  & n307;
  assign n309 = \V120(21)  & n308;
  assign n310 = \V168(13)  & n309;
  assign n311 = ~n306 & ~n310;
  assign n312 = ~n304 & n311;
  assign n313 = ~n303 & n312;
  assign n314 = \V189(2)  & \V189(0) ;
  assign n315 = ~n313 & n314;
  assign n316 = \V189(1)  & n315;
  assign n317 = ~n300 & ~n316;
  assign n318 = ~n286 & n317;
  assign n319 = ~n283 & n318;
  assign n320 = ~n282 & n319;
  assign n321 = ~n280 & n320;
  assign \V198(2)  = n276 | ~n321;
  assign n323 = \V156(9)  & \V120(0) ;
  assign n324 = \V88(0)  & n323;
  assign n325 = \V156(8)  & n324;
  assign n326 = \V56(26)  & \V28(26) ;
  assign n327 = \V156(8)  & \V28(27) ;
  assign n328 = \V56(27)  & n327;
  assign n329 = \V156(8)  & \V156(10) ;
  assign n330 = \V88(1)  & n329;
  assign n331 = \V120(1)  & n330;
  assign n332 = \V156(9)  & n331;
  assign n333 = ~n328 & ~n332;
  assign n334 = ~n326 & n333;
  assign n335 = ~n325 & n334;
  assign n336 = \V186(1)  & ~n335;
  assign n337 = \V186(0)  & n336;
  assign n338 = \V156(2)  & \V156(0) ;
  assign n339 = \V28(21)  & n338;
  assign n340 = \V56(21)  & n339;
  assign n341 = \V156(1)  & n340;
  assign n342 = \V156(0)  & \V28(19) ;
  assign n343 = \V56(19)  & n342;
  assign n344 = \V56(18)  & \V28(18) ;
  assign n345 = \V56(20)  & \V156(1) ;
  assign n346 = \V28(20)  & n345;
  assign n347 = \V156(0)  & n346;
  assign n348 = \V56(24)  & \V156(5) ;
  assign n349 = \V28(24)  & n348;
  assign n350 = \V156(4)  & n349;
  assign n351 = \V56(22)  & \V28(22) ;
  assign n352 = \V156(4)  & \V28(23) ;
  assign n353 = \V56(23)  & n352;
  assign n354 = \V156(4)  & \V156(6) ;
  assign n355 = \V28(25)  & n354;
  assign n356 = \V56(25)  & n355;
  assign n357 = \V156(5)  & n356;
  assign n358 = ~n353 & ~n357;
  assign n359 = ~n351 & n358;
  assign n360 = ~n350 & n359;
  assign n361 = \V186(0)  & ~n360;
  assign n362 = \V156(13)  & \V120(4) ;
  assign n363 = \V88(4)  & n362;
  assign n364 = \V156(12)  & n363;
  assign n365 = \V88(2)  & \V120(2) ;
  assign n366 = \V88(3)  & \V156(12) ;
  assign n367 = \V120(3)  & n366;
  assign n368 = \V156(12)  & \V156(14) ;
  assign n369 = \V88(5)  & n368;
  assign n370 = \V120(5)  & n369;
  assign n371 = \V156(13)  & n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~n365 & n372;
  assign n374 = ~n364 & n373;
  assign n375 = \V186(2)  & \V186(0) ;
  assign n376 = ~n374 & n375;
  assign n377 = \V186(1)  & n376;
  assign n378 = ~n361 & ~n377;
  assign n379 = ~n347 & n378;
  assign n380 = ~n344 & n379;
  assign n381 = ~n343 & n380;
  assign n382 = ~n341 & n381;
  assign \V198(1)  = n337 | ~n382;
  assign n384 = \V56(12)  & \V144(9) ;
  assign n385 = \V28(12)  & n384;
  assign n386 = \V144(8)  & n385;
  assign n387 = \V56(10)  & \V28(10) ;
  assign n388 = \V28(11)  & \V144(8) ;
  assign n389 = \V56(11)  & n388;
  assign n390 = \V144(10)  & \V144(8) ;
  assign n391 = \V28(13)  & n390;
  assign n392 = \V56(13)  & n391;
  assign n393 = \V144(9)  & n392;
  assign n394 = ~n389 & ~n393;
  assign n395 = ~n387 & n394;
  assign n396 = ~n386 & n395;
  assign n397 = \V183(1)  & ~n396;
  assign n398 = \V183(0)  & n397;
  assign n399 = \V144(2)  & \V144(0) ;
  assign n400 = \V28(5)  & n399;
  assign n401 = \V56(5)  & n400;
  assign n402 = \V144(1)  & n401;
  assign n403 = \V144(0)  & \V28(3) ;
  assign n404 = \V56(3)  & n403;
  assign n405 = \V56(2)  & \V28(2) ;
  assign n406 = \V56(4)  & \V144(1) ;
  assign n407 = \V28(4)  & n406;
  assign n408 = \V144(0)  & n407;
  assign n409 = \V56(8)  & \V144(5) ;
  assign n410 = \V28(8)  & n409;
  assign n411 = \V144(4)  & n410;
  assign n412 = \V56(6)  & \V28(6) ;
  assign n413 = \V144(4)  & \V28(7) ;
  assign n414 = \V56(7)  & n413;
  assign n415 = \V144(4)  & \V144(6) ;
  assign n416 = \V28(9)  & n415;
  assign n417 = \V56(9)  & n416;
  assign n418 = \V144(5)  & n417;
  assign n419 = ~n414 & ~n418;
  assign n420 = ~n412 & n419;
  assign n421 = ~n411 & n420;
  assign n422 = \V183(0)  & ~n421;
  assign n423 = \V144(13)  & \V56(16) ;
  assign n424 = \V28(16)  & n423;
  assign n425 = \V144(12)  & n424;
  assign n426 = \V56(14)  & \V28(14) ;
  assign n427 = \V144(12)  & \V28(15) ;
  assign n428 = \V56(15)  & n427;
  assign n429 = \V144(12)  & \V144(14) ;
  assign n430 = \V28(17)  & n429;
  assign n431 = \V56(17)  & n430;
  assign n432 = \V144(13)  & n431;
  assign n433 = ~n428 & ~n432;
  assign n434 = ~n426 & n433;
  assign n435 = ~n425 & n434;
  assign n436 = \V183(2)  & \V183(0) ;
  assign n437 = ~n435 & n436;
  assign n438 = \V183(1)  & n437;
  assign n439 = ~n422 & ~n438;
  assign n440 = ~n408 & n439;
  assign n441 = ~n405 & n440;
  assign n442 = ~n404 & n441;
  assign n443 = ~n402 & n442;
  assign \V198(0)  = n398 | ~n443;
endmodule


