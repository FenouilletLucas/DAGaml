// Benchmark "DES" written by ABC on Tue May 16 16:07:49 2017

module DES ( 
    \data<63> , \data<61> , \data<62> , \reset<0> , \outreg<58> ,
    \inreg<0> , \outreg<57> , \inreg<1> , \outreg<56> , \inreg<2> ,
    \outreg<55> , \inreg<3> , \inreg<4> , \inreg<5> , \inreg<6> ,
    \outreg<59> , \inreg<7> , \outreg<50> , \inreg<8> , \inreg<9> ,
    \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \load_key<0> ,
    \outreg<60> , \outreg<63> , \outreg<62> , \outreg<61> , \D<0> , \D<1> ,
    \D<2> , \D<3> , \D<4> , \D<5> , \D<6> , \C<10> , \D<7> , \C<11> ,
    \D<8> , \C<12> , \D<9> , \C<13> , \C<14> , \C<15> , \C<16> , \C<17> ,
    \C<18> , \C<19> , \outreg<18> , \outreg<17> , \outreg<16> ,
    \outreg<15> , \C<20> , \outreg<19> , \C<21> , \outreg<10> , \C<22> ,
    \C<23> , \C<24> , \C<25> , \outreg<14> , \C<26> , \outreg<13> ,
    \C<27> , \outreg<12> , \outreg<11> , \outreg<28> , \outreg<27> ,
    \outreg<26> , \outreg<25> , \outreg<29> , \outreg<20> , \data<3> ,
    \data<4> , \data<1> , \outreg<24> , \data<2> , \outreg<23> ,
    \outreg<22> , \data<0> , \outreg<21> , \outreg<38> , \outreg<37> ,
    \outreg<36> , \outreg<35> , \data<9> , \data<7> , \data<8> ,
    \outreg<39> , \data<5> , \outreg<30> , \data<6> , \outreg<34> ,
    \outreg<33> , \outreg<32> , \outreg<31> , \outreg<48> , \outreg<47> ,
    \outreg<46> , \outreg<45> , \outreg<49> , \outreg<40> , \outreg<44> ,
    \outreg<43> , \outreg<42> , \outreg<41> , \D<10> , \D<11> , \D<12> ,
    \D<13> , \D<14> , \D<15> , \D<16> , \D<17> , \D<18> , \D<19> , \D<20> ,
    \D<21> , \data_in<7> , \D<22> , \D<23> , \data_in<5> , \D<24> ,
    \data_in<6> , \D<25> , \D<26> , \D<27> , \data_in<0> , \data_in<3> ,
    \data_in<4> , \data_in<1> , \data_in<2> , \data<37> , \data<38> ,
    \data<35> , \data<36> , \data<39> , \data<30> , \data<33> , \data<34> ,
    \data<31> , \data<32> , \data<47> , \data<48> , \data<45> , \data<46> ,
    \data<49> , \data<40> , \data<43> , \data<44> , \data<41> , \data<42> ,
    \data<17> , \data<18> , \data<15> , \count<0> , \data<16> , \count<3> ,
    \data<19> , \count<1> , \count<2> , \data<10> , \data<13> , \data<14> ,
    \data<11> , \data<12> , \data<27> , \data<28> , \data<25> , \data<26> ,
    \data<29> , \data<20> , \data<23> , \data<24> , \data<21> , \data<22> ,
    \C<0> , \C<1> , \C<2> , \C<3> , \C<4> , \C<5> , \C<6> , \C<7> , \C<8> ,
    \C<9> , \inreg<12> , \inreg<11> , \inreg<14> , \inreg<13> ,
    \inreg<10> , \inreg<19> , \inreg<16> , \inreg<15> , \inreg<18> ,
    \inreg<17> , \inreg<22> , \inreg<21> , \inreg<24> , \inreg<23> ,
    \inreg<20> , \inreg<29> , \inreg<26> , \inreg<25> , \outreg<9> ,
    \inreg<28> , \inreg<27> , \inreg<32> , \inreg<31> , \outreg<5> ,
    \inreg<34> , \outreg<6> , \inreg<33> , \outreg<7> , \outreg<8> ,
    \outreg<1> , \inreg<30> , \outreg<2> , \outreg<3> , \outreg<4> ,
    \inreg<39> , \inreg<36> , \outreg<0> , \inreg<35> , \inreg<38> ,
    \inreg<37> , \inreg<42> , \inreg<41> , \inreg<44> , \inreg<43> ,
    \inreg<40> , \inreg<49> , \inreg<46> , \inreg<45> , \encrypt_mode<0> ,
    \inreg<48> , \inreg<47> , \inreg<52> , \inreg<51> , \inreg<54> ,
    \inreg<53> , \inreg<50> , \inreg<55> , \data<57> , \data<58> ,
    \data<55> , \data<56> , \encrypt<0> , \data<59> , \data<50> ,
    \data<53> , \data<54> , \data<51> , \data<52> , \data<60> ,
    \data_new<25> , \inreg_new<45> , \data_new<26> , \data_new<13> ,
    \data_new<14> , \data_new<11> , \inreg_new<49> , \data_new<12> ,
    \inreg_new<30> , \outreg_new<11> , \count_new<0> , \outreg_new<12> ,
    \data_new<10> , \outreg_new<13> , \outreg_new<14> , \inreg_new<34> ,
    \count_new<3> , \inreg_new<33> , \inreg_new<32> , \count_new<1> ,
    \data_new<19> , \inreg_new<31> , \count_new<2> , \outreg_new<10> ,
    \inreg_new<38> , \outreg_new<19> , \data_new<17> , \inreg_new<37> ,
    \data_new<18> , \inreg_new<36> , \data_new<15> , \inreg_new<35> ,
    \data_new<16> , \outreg_new<15> , \outreg_new<16> , \outreg_new<17> ,
    \inreg_new<39> , \outreg_new<18> , \outreg_new<21> , \outreg_new<22> ,
    \outreg_new<23> , \outreg_new<24> , \outreg_new<20> , \outreg_new<29> ,
    \outreg_new<25> , \outreg_new<26> , \outreg_new<27> , \outreg_new<28> ,
    \outreg_new<31> , \outreg_new<32> , \outreg_new<33> , \outreg_new<34> ,
    \outreg_new<30> , \outreg_new<39> , \outreg_new<35> , \outreg_new<36> ,
    \outreg_new<37> , \outreg_new<38> , \outreg_new<41> , \outreg_new<42> ,
    \outreg_new<43> , \outreg_new<44> , \outreg_new<40> , \outreg_new<49> ,
    \outreg_new<45> , \outreg_new<46> , \outreg_new<47> , \outreg_new<48> ,
    \C_new<23> , \C_new<24> , \C_new<21> , \C_new<22> , \C_new<20> ,
    \data_new<4> , \data_new<3> , \C_new<27> , \data_new<2> ,
    \data_new<1> , \C_new<25> , \data_new<0> , \C_new<26> , \C_new<13> ,
    \C_new<14> , \C_new<11> , \C_new<12> , \C_new<10> , \data_new<9> ,
    \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> ,
    \C_new<19> , \C_new<17> , \C_new<18> , \C_new<15> , \C_new<16> ,
    \D_new<13> , \D_new<14> , \D_new<11> , \D_new<12> , \D_new<10> ,
    \data_new<63> , \data_new<61> , \data_new<62> , \D_new<19> ,
    \data_new<60> , \D_new<17> , \D_new<18> , \D_new<15> , \D_new<16> ,
    \D_new<23> , \D_new<24> , \D_new<21> , \D_new<22> , \D_new<20> ,
    \data_new<53> , \data_new<54> , \data_new<51> , \data_new<52> ,
    \data_new<50> , \D_new<27> , \D_new<25> , \D_new<26> , \data_new<59> ,
    \data_new<57> , \data_new<58> , \data_new<55> , \data_new<56> ,
    \D_new<7> , \C_new<6> , \D_new<8> , \C_new<5> , \D_new<5> , \C_new<8> ,
    \D_new<6> , \C_new<7> , \C_new<9> , \D_new<9> , \D_new<0> , \C_new<0> ,
    \D_new<3> , \C_new<2> , \D_new<4> , \C_new<1> , \D_new<1> , \C_new<4> ,
    \D_new<2> , \C_new<3> , \inreg_new<50> , \inreg_new<9> ,
    \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<6> ,
    \inreg_new<51> , \inreg_new<5> , \inreg_new<8> , \inreg_new<7> ,
    \inreg_new<2> , \inreg_new<55> , \inreg_new<1> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<0> , \encrypt_mode_new<0> , \outreg_new<9> ,
    \outreg_new<51> , \outreg_new<52> , \outreg_new<53> , \outreg_new<5> ,
    \outreg_new<54> , \outreg_new<6> , \outreg_new<7> , \outreg_new<8> ,
    \outreg_new<1> , \outreg_new<50> , \outreg_new<2> , \outreg_new<59> ,
    \outreg_new<3> , \outreg_new<4> , \outreg_new<55> , \data_new<43> ,
    \outreg_new<56> , \data_new<44> , \outreg_new<0> , \outreg_new<57> ,
    \data_new<41> , \outreg_new<58> , \data_new<42> , \inreg_new<20> ,
    \outreg_new<61> , \outreg_new<62> , \data_new<40> , \outreg_new<63> ,
    \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \data_new<49> ,
    \inreg_new<21> , \outreg_new<60> , \inreg_new<28> , \data_new<47> ,
    \inreg_new<27> , \data_new<48> , \inreg_new<26> , \data_new<45> ,
    \inreg_new<25> , \data_new<46> , \data_new<33> , \data_new<34> ,
    \data_new<31> , \inreg_new<29> , \data_new<32> , \inreg_new<10> ,
    \data_new<30> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \data_new<39> , \inreg_new<11> , \inreg_new<18> , \data_new<37> ,
    \inreg_new<17> , \data_new<38> , \inreg_new<16> , \data_new<35> ,
    \inreg_new<15> , \data_new<36> , \data_new<23> , \data_new<24> ,
    \data_new<21> , \inreg_new<19> , \data_new<22> , \inreg_new<40> ,
    \data_new<20> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> ,
    \data_new<29> , \inreg_new<41> , \inreg_new<48> , \data_new<27> ,
    \inreg_new<47> , \data_new<28> , \inreg_new<46>   );
  input  \data<63> , \data<61> , \data<62> , \reset<0> , \outreg<58> ,
    \inreg<0> , \outreg<57> , \inreg<1> , \outreg<56> , \inreg<2> ,
    \outreg<55> , \inreg<3> , \inreg<4> , \inreg<5> , \inreg<6> ,
    \outreg<59> , \inreg<7> , \outreg<50> , \inreg<8> , \inreg<9> ,
    \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \load_key<0> ,
    \outreg<60> , \outreg<63> , \outreg<62> , \outreg<61> , \D<0> , \D<1> ,
    \D<2> , \D<3> , \D<4> , \D<5> , \D<6> , \C<10> , \D<7> , \C<11> ,
    \D<8> , \C<12> , \D<9> , \C<13> , \C<14> , \C<15> , \C<16> , \C<17> ,
    \C<18> , \C<19> , \outreg<18> , \outreg<17> , \outreg<16> ,
    \outreg<15> , \C<20> , \outreg<19> , \C<21> , \outreg<10> , \C<22> ,
    \C<23> , \C<24> , \C<25> , \outreg<14> , \C<26> , \outreg<13> ,
    \C<27> , \outreg<12> , \outreg<11> , \outreg<28> , \outreg<27> ,
    \outreg<26> , \outreg<25> , \outreg<29> , \outreg<20> , \data<3> ,
    \data<4> , \data<1> , \outreg<24> , \data<2> , \outreg<23> ,
    \outreg<22> , \data<0> , \outreg<21> , \outreg<38> , \outreg<37> ,
    \outreg<36> , \outreg<35> , \data<9> , \data<7> , \data<8> ,
    \outreg<39> , \data<5> , \outreg<30> , \data<6> , \outreg<34> ,
    \outreg<33> , \outreg<32> , \outreg<31> , \outreg<48> , \outreg<47> ,
    \outreg<46> , \outreg<45> , \outreg<49> , \outreg<40> , \outreg<44> ,
    \outreg<43> , \outreg<42> , \outreg<41> , \D<10> , \D<11> , \D<12> ,
    \D<13> , \D<14> , \D<15> , \D<16> , \D<17> , \D<18> , \D<19> , \D<20> ,
    \D<21> , \data_in<7> , \D<22> , \D<23> , \data_in<5> , \D<24> ,
    \data_in<6> , \D<25> , \D<26> , \D<27> , \data_in<0> , \data_in<3> ,
    \data_in<4> , \data_in<1> , \data_in<2> , \data<37> , \data<38> ,
    \data<35> , \data<36> , \data<39> , \data<30> , \data<33> , \data<34> ,
    \data<31> , \data<32> , \data<47> , \data<48> , \data<45> , \data<46> ,
    \data<49> , \data<40> , \data<43> , \data<44> , \data<41> , \data<42> ,
    \data<17> , \data<18> , \data<15> , \count<0> , \data<16> , \count<3> ,
    \data<19> , \count<1> , \count<2> , \data<10> , \data<13> , \data<14> ,
    \data<11> , \data<12> , \data<27> , \data<28> , \data<25> , \data<26> ,
    \data<29> , \data<20> , \data<23> , \data<24> , \data<21> , \data<22> ,
    \C<0> , \C<1> , \C<2> , \C<3> , \C<4> , \C<5> , \C<6> , \C<7> , \C<8> ,
    \C<9> , \inreg<12> , \inreg<11> , \inreg<14> , \inreg<13> ,
    \inreg<10> , \inreg<19> , \inreg<16> , \inreg<15> , \inreg<18> ,
    \inreg<17> , \inreg<22> , \inreg<21> , \inreg<24> , \inreg<23> ,
    \inreg<20> , \inreg<29> , \inreg<26> , \inreg<25> , \outreg<9> ,
    \inreg<28> , \inreg<27> , \inreg<32> , \inreg<31> , \outreg<5> ,
    \inreg<34> , \outreg<6> , \inreg<33> , \outreg<7> , \outreg<8> ,
    \outreg<1> , \inreg<30> , \outreg<2> , \outreg<3> , \outreg<4> ,
    \inreg<39> , \inreg<36> , \outreg<0> , \inreg<35> , \inreg<38> ,
    \inreg<37> , \inreg<42> , \inreg<41> , \inreg<44> , \inreg<43> ,
    \inreg<40> , \inreg<49> , \inreg<46> , \inreg<45> , \encrypt_mode<0> ,
    \inreg<48> , \inreg<47> , \inreg<52> , \inreg<51> , \inreg<54> ,
    \inreg<53> , \inreg<50> , \inreg<55> , \data<57> , \data<58> ,
    \data<55> , \data<56> , \encrypt<0> , \data<59> , \data<50> ,
    \data<53> , \data<54> , \data<51> , \data<52> , \data<60> ;
  output \data_new<25> , \inreg_new<45> , \data_new<26> , \data_new<13> ,
    \data_new<14> , \data_new<11> , \inreg_new<49> , \data_new<12> ,
    \inreg_new<30> , \outreg_new<11> , \count_new<0> , \outreg_new<12> ,
    \data_new<10> , \outreg_new<13> , \outreg_new<14> , \inreg_new<34> ,
    \count_new<3> , \inreg_new<33> , \inreg_new<32> , \count_new<1> ,
    \data_new<19> , \inreg_new<31> , \count_new<2> , \outreg_new<10> ,
    \inreg_new<38> , \outreg_new<19> , \data_new<17> , \inreg_new<37> ,
    \data_new<18> , \inreg_new<36> , \data_new<15> , \inreg_new<35> ,
    \data_new<16> , \outreg_new<15> , \outreg_new<16> , \outreg_new<17> ,
    \inreg_new<39> , \outreg_new<18> , \outreg_new<21> , \outreg_new<22> ,
    \outreg_new<23> , \outreg_new<24> , \outreg_new<20> , \outreg_new<29> ,
    \outreg_new<25> , \outreg_new<26> , \outreg_new<27> , \outreg_new<28> ,
    \outreg_new<31> , \outreg_new<32> , \outreg_new<33> , \outreg_new<34> ,
    \outreg_new<30> , \outreg_new<39> , \outreg_new<35> , \outreg_new<36> ,
    \outreg_new<37> , \outreg_new<38> , \outreg_new<41> , \outreg_new<42> ,
    \outreg_new<43> , \outreg_new<44> , \outreg_new<40> , \outreg_new<49> ,
    \outreg_new<45> , \outreg_new<46> , \outreg_new<47> , \outreg_new<48> ,
    \C_new<23> , \C_new<24> , \C_new<21> , \C_new<22> , \C_new<20> ,
    \data_new<4> , \data_new<3> , \C_new<27> , \data_new<2> ,
    \data_new<1> , \C_new<25> , \data_new<0> , \C_new<26> , \C_new<13> ,
    \C_new<14> , \C_new<11> , \C_new<12> , \C_new<10> , \data_new<9> ,
    \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> ,
    \C_new<19> , \C_new<17> , \C_new<18> , \C_new<15> , \C_new<16> ,
    \D_new<13> , \D_new<14> , \D_new<11> , \D_new<12> , \D_new<10> ,
    \data_new<63> , \data_new<61> , \data_new<62> , \D_new<19> ,
    \data_new<60> , \D_new<17> , \D_new<18> , \D_new<15> , \D_new<16> ,
    \D_new<23> , \D_new<24> , \D_new<21> , \D_new<22> , \D_new<20> ,
    \data_new<53> , \data_new<54> , \data_new<51> , \data_new<52> ,
    \data_new<50> , \D_new<27> , \D_new<25> , \D_new<26> , \data_new<59> ,
    \data_new<57> , \data_new<58> , \data_new<55> , \data_new<56> ,
    \D_new<7> , \C_new<6> , \D_new<8> , \C_new<5> , \D_new<5> , \C_new<8> ,
    \D_new<6> , \C_new<7> , \C_new<9> , \D_new<9> , \D_new<0> , \C_new<0> ,
    \D_new<3> , \C_new<2> , \D_new<4> , \C_new<1> , \D_new<1> , \C_new<4> ,
    \D_new<2> , \C_new<3> , \inreg_new<50> , \inreg_new<9> ,
    \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<6> ,
    \inreg_new<51> , \inreg_new<5> , \inreg_new<8> , \inreg_new<7> ,
    \inreg_new<2> , \inreg_new<55> , \inreg_new<1> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<0> , \encrypt_mode_new<0> , \outreg_new<9> ,
    \outreg_new<51> , \outreg_new<52> , \outreg_new<53> , \outreg_new<5> ,
    \outreg_new<54> , \outreg_new<6> , \outreg_new<7> , \outreg_new<8> ,
    \outreg_new<1> , \outreg_new<50> , \outreg_new<2> , \outreg_new<59> ,
    \outreg_new<3> , \outreg_new<4> , \outreg_new<55> , \data_new<43> ,
    \outreg_new<56> , \data_new<44> , \outreg_new<0> , \outreg_new<57> ,
    \data_new<41> , \outreg_new<58> , \data_new<42> , \inreg_new<20> ,
    \outreg_new<61> , \outreg_new<62> , \data_new<40> , \outreg_new<63> ,
    \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \data_new<49> ,
    \inreg_new<21> , \outreg_new<60> , \inreg_new<28> , \data_new<47> ,
    \inreg_new<27> , \data_new<48> , \inreg_new<26> , \data_new<45> ,
    \inreg_new<25> , \data_new<46> , \data_new<33> , \data_new<34> ,
    \data_new<31> , \inreg_new<29> , \data_new<32> , \inreg_new<10> ,
    \data_new<30> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \data_new<39> , \inreg_new<11> , \inreg_new<18> , \data_new<37> ,
    \inreg_new<17> , \data_new<38> , \inreg_new<16> , \data_new<35> ,
    \inreg_new<15> , \data_new<36> , \data_new<23> , \data_new<24> ,
    \data_new<21> , \inreg_new<19> , \data_new<22> , \inreg_new<40> ,
    \data_new<20> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> ,
    \data_new<29> , \inreg_new<41> , \inreg_new<48> , \data_new<27> ,
    \inreg_new<47> , \data_new<28> , \inreg_new<46> ;
  wire n502, n503, n504, n505, n506, n508, n509, n510, n511, n513, n514,
    n516, n517, n519, n520, n522, n523, n525, n526, n528, n529, n531, n532,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n674, n675, n677, n678, n679,
    n680, n682, n683, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n827, n828, n829, n830, n832, n833, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n846, n847, n849, n850, n852, n853, n854, n856,
    n857, n859, n860, n862, n863, n864, n865, n866, n867, n868, n870, n871,
    n872, n873, n875, n876, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1025,
    n1026, n1028, n1029, n1031, n1032, n1034, n1035, n1037, n1038, n1040,
    n1041, n1043, n1044, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1110, n1111, n1112, n1113,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1261, n1262, n1264, n1265, n1266,
    n1267, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1413, n1414, n1415, n1416, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1478, n1479, n1480,
    n1481, n1483, n1484, n1485, n1486, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1600, n1601, n1602, n1603, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1750, n1751, n1752, n1753, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1901, n1902, n1903, n1904, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1966, n1967, n1968, n1969, n1971,
    n1972, n1973, n1974, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2097, n2098, n2099, n2100, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2243, n2244, n2245, n2246,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2306, n2307, n2308,
    n2309, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2359, n2360,
    n2361, n2362, n2364, n2365, n2366, n2367, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2460, n2461, n2462, n2463, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2509, n2510, n2511, n2512, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2665, n2666, n2668, n2669, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2702, n2703, n2705, n2706,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2732, n2733, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2889, n2890, n2892, n2893, n2895, n2896, n2898,
    n2899, n2901, n2902, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3201,
    n3202, n3203, n3204, n3205, n3206, n3208, n3209, n3210, n3211, n3212,
    n3213, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3248, n3249, n3250, n3251, n3252, n3253, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
    n3401, n3402, n3403, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
    n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3473, n3474,
    n3475, n3476, n3477, n3478, n3480, n3481, n3482, n3483, n3484, n3485,
    n3487, n3488, n3489, n3490, n3491, n3492, n3494, n3495, n3496, n3497,
    n3498, n3499, n3501, n3502, n3503, n3504, n3505, n3506, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
    n3582, n3584, n3585, n3586, n3587, n3588, n3589, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3654,
    n3655, n3656, n3657, n3658, n3659, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
    n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4006, n4007,
    n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
    n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
    n4195, n4196, n4197, n4198, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4240, n4241, n4243, n4244, n4246, n4247, n4249, n4250,
    n4252, n4253, n4255, n4256, n4258, n4259, n4261, n4262, n4264, n4265,
    n4267, n4268, n4270, n4271, n4273, n4274, n4276, n4277, n4279, n4280,
    n4282, n4283, n4285, n4286, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4392, n4393, n4394, n4395, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4450, n4451, n4452, n4453, n4455, n4456, n4457, n4458, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467, n4469, n4470, n4471, n4472,
    n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4518, n4519, n4520, n4521, n4523, n4524, n4525,
    n4526, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
    n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
    n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4618,
    n4619, n4620, n4621, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4632, n4633, n4634, n4635, n4636, n4637, n4639, n4640, n4642,
    n4643, n4644, n4645, n4646, n4647, n4649, n4650, n4651, n4652, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
    n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4695,
    n4696, n4697, n4698, n4699, n4700, n4702, n4703, n4705, n4706, n4707,
    n4708, n4709, n4710, n4712, n4713, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4756, n4757, n4759, n4760, n4761,
    n4762, n4763, n4764, n4766, n4767, n4768, n4769, n4770, n4771, n4773,
    n4774, n4776, n4777, n4779, n4780, n4782, n4783, n4784, n4785, n4786,
    n4787, n4789, n4790, n4792, n4793, n4795, n4796, n4798, n4799, n4800,
    n4801, n4802, n4803, n4805, n4806, n4808, n4809, n4810, n4811, n4812,
    n4813, n4815, n4816, n4818, n4819, n4820, n4821, n4822, n4823, n4825,
    n4826, n4828, n4829, n4830, n4831, n4832, n4833, n4835, n4836, n4837,
    n4838, n4839, n4840, n4842, n4843, n4844, n4845, n4846, n4847, n4849,
    n4850, n4852, n4853, n4855, n4856, n4857, n4858, n4859, n4860, n4862,
    n4863, n4865, n4866, n4868, n4869, n4871, n4872, n4874, n4875, n4877,
    n4878, n4879, n4880, n4881, n4882, n4884, n4885, n4887, n4888, n4890,
    n4891, n4892, n4893, n4894, n4895, n4897, n4898, n4900, n4901, n4902,
    n4903, n4904, n4905, n4907, n4908, n4910, n4911, n4912, n4913, n4914,
    n4915, n4917, n4918, n4920, n4921, n4922, n4923, n4924, n4925, n4927,
    n4928, n4930, n4931, n4933, n4934, n4936, n4937, n4939, n4940, n4942,
    n4943, n4945, n4946, n4948, n4949, n4951, n4952, n4954, n4955, n4957,
    n4958, n4960, n4961, n4963, n4964, n4966, n4967, n4969, n4970, n4972,
    n4973, n4975, n4976;
  assign n502 = \count<0>  & \count<1> ;
  assign n503 = \count<2>  & n502;
  assign n504 = \count<3>  & n503;
  assign n505 = \data<57>  & ~n504;
  assign n506 = \inreg<47>  & n504;
  assign \data_new<25>  = n505 | n506;
  assign n508 = ~\count<0>  & ~n504;
  assign n509 = \inreg<45>  & n508;
  assign n510 = \count<0>  & ~n504;
  assign n511 = \inreg<37>  & n510;
  assign \inreg_new<45>  = n509 | n511;
  assign n513 = \data<58>  & ~n504;
  assign n514 = \inreg<39>  & n504;
  assign \data_new<26>  = n513 | n514;
  assign n516 = \data<45>  & ~n504;
  assign n517 = \inreg<11>  & n504;
  assign \data_new<13>  = n516 | n517;
  assign n519 = \data<46>  & ~n504;
  assign n520 = \inreg<3>  & n504;
  assign \data_new<14>  = n519 | n520;
  assign n522 = \data<43>  & ~n504;
  assign n523 = \inreg<27>  & n504;
  assign \data_new<11>  = n522 | n523;
  assign n525 = \inreg<49>  & n508;
  assign n526 = \inreg<41>  & n510;
  assign \inreg_new<49>  = n525 | n526;
  assign n528 = \data<44>  & ~n504;
  assign n529 = \inreg<19>  & n504;
  assign \data_new<12>  = n528 | n529;
  assign n531 = \inreg<30>  & n508;
  assign n532 = \inreg<22>  & n510;
  assign \inreg_new<30>  = n531 | n532;
  assign n534 = \D<3>  & ~\data<32> ;
  assign n535 = ~\D<3>  & \data<32> ;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~\data<63>  & \D<0> ;
  assign n538 = \data<63>  & ~\D<0> ;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~\data<62>  & \D<7> ;
  assign n541 = \data<62>  & ~\D<7> ;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~\data<61>  & \D<21> ;
  assign n544 = \data<61>  & ~\D<21> ;
  assign n545 = ~n543 & ~n544;
  assign n546 = \D<13>  & ~\data<60> ;
  assign n547 = ~\D<13>  & \data<60> ;
  assign n548 = ~n546 & ~n547;
  assign n549 = \D<17>  & ~\data<59> ;
  assign n550 = ~\D<17>  & \data<59> ;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n548 & ~n551;
  assign n553 = ~n545 & n552;
  assign n554 = ~n542 & n553;
  assign n555 = ~n539 & n554;
  assign n556 = ~n536 & n555;
  assign n557 = n539 & n554;
  assign n558 = ~n536 & n557;
  assign n559 = n542 & n553;
  assign n560 = n539 & n559;
  assign n561 = ~n536 & n560;
  assign n562 = n545 & n552;
  assign n563 = n542 & n562;
  assign n564 = n539 & n563;
  assign n565 = ~n536 & n564;
  assign n566 = n548 & ~n551;
  assign n567 = ~n545 & n566;
  assign n568 = n542 & n567;
  assign n569 = ~n539 & n568;
  assign n570 = ~n536 & n569;
  assign n571 = n545 & n566;
  assign n572 = ~n542 & n571;
  assign n573 = ~n539 & n572;
  assign n574 = ~n536 & n573;
  assign n575 = n539 & n572;
  assign n576 = ~n536 & n575;
  assign n577 = ~n539 & n559;
  assign n578 = n536 & n577;
  assign n579 = n536 & n560;
  assign n580 = ~n542 & n562;
  assign n581 = n539 & n580;
  assign n582 = n536 & n581;
  assign n583 = ~n539 & n563;
  assign n584 = n536 & n583;
  assign n585 = ~n542 & n567;
  assign n586 = n539 & n585;
  assign n587 = n536 & n586;
  assign n588 = n542 & n571;
  assign n589 = ~n539 & n588;
  assign n590 = n536 & n589;
  assign n591 = n539 & n588;
  assign n592 = n536 & n591;
  assign n593 = ~n548 & n551;
  assign n594 = ~n545 & n593;
  assign n595 = n542 & n594;
  assign n596 = ~n539 & n595;
  assign n597 = ~n536 & n596;
  assign n598 = n545 & n593;
  assign n599 = ~n542 & n598;
  assign n600 = ~n539 & n599;
  assign n601 = ~n536 & n600;
  assign n602 = n539 & n599;
  assign n603 = ~n536 & n602;
  assign n604 = n548 & n551;
  assign n605 = ~n545 & n604;
  assign n606 = ~n542 & n605;
  assign n607 = n539 & n606;
  assign n608 = ~n536 & n607;
  assign n609 = n542 & n605;
  assign n610 = ~n539 & n609;
  assign n611 = ~n536 & n610;
  assign n612 = n539 & n609;
  assign n613 = ~n536 & n612;
  assign n614 = n545 & n604;
  assign n615 = n542 & n614;
  assign n616 = ~n539 & n615;
  assign n617 = ~n536 & n616;
  assign n618 = ~n542 & n594;
  assign n619 = ~n539 & n618;
  assign n620 = n536 & n619;
  assign n621 = n536 & n600;
  assign n622 = n536 & n602;
  assign n623 = n542 & n598;
  assign n624 = n539 & n623;
  assign n625 = n536 & n624;
  assign n626 = n536 & n607;
  assign n627 = n536 & n610;
  assign n628 = n536 & n612;
  assign n629 = n536 & n616;
  assign n630 = ~n539 & n585;
  assign n631 = n536 & n630;
  assign n632 = ~n536 & n591;
  assign n633 = ~n627 & ~n628;
  assign n634 = ~n626 & n633;
  assign n635 = ~n625 & n634;
  assign n636 = ~n622 & n635;
  assign n637 = ~n621 & n636;
  assign n638 = ~n620 & n637;
  assign n639 = ~n617 & n638;
  assign n640 = ~n613 & n639;
  assign n641 = ~n611 & n640;
  assign n642 = ~n608 & n641;
  assign n643 = ~n603 & n642;
  assign n644 = ~n601 & n643;
  assign n645 = ~n597 & n644;
  assign n646 = ~n592 & n645;
  assign n647 = ~n590 & n646;
  assign n648 = ~n587 & n647;
  assign n649 = ~n584 & n648;
  assign n650 = ~n582 & n649;
  assign n651 = ~n579 & n650;
  assign n652 = ~n578 & n651;
  assign n653 = ~n576 & n652;
  assign n654 = ~n574 & n653;
  assign n655 = ~n570 & n654;
  assign n656 = ~n565 & n655;
  assign n657 = ~n561 & n656;
  assign n658 = ~n558 & n657;
  assign n659 = ~n556 & n658;
  assign n660 = ~n536 & n619;
  assign n661 = n659 & ~n660;
  assign n662 = ~n632 & n661;
  assign n663 = ~n631 & n662;
  assign n664 = ~n629 & n663;
  assign n665 = \data<14>  & n504;
  assign n666 = n664 & n665;
  assign n667 = ~\data<14>  & n504;
  assign n668 = ~n664 & n667;
  assign n669 = \outreg<19>  & n510;
  assign n670 = \outreg<11>  & n508;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n668 & n671;
  assign \outreg_new<11>  = n666 | ~n672;
  assign n674 = \load_key<0>  & n504;
  assign n675 = ~\reset<0>  & ~n674;
  assign \count_new<0>  = ~\count<0>  & n675;
  assign n677 = \outreg<20>  & n510;
  assign n678 = \outreg<12>  & n508;
  assign n679 = \data<54>  & n504;
  assign n680 = ~n678 & ~n679;
  assign \outreg_new<12>  = n677 | ~n680;
  assign n682 = \data<42>  & ~n504;
  assign n683 = \inreg<35>  & n504;
  assign \data_new<10>  = n682 | n683;
  assign n685 = ~\data<36>  & \C<4> ;
  assign n686 = \data<36>  & ~\C<4> ;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~\data<35>  & \C<0> ;
  assign n689 = \data<35>  & ~\C<0> ;
  assign n690 = ~n688 & ~n689;
  assign n691 = \C<23>  & ~\data<34> ;
  assign n692 = ~\C<23>  & \data<34> ;
  assign n693 = ~n691 & ~n692;
  assign n694 = \C<10>  & ~\data<33> ;
  assign n695 = ~\C<10>  & \data<33> ;
  assign n696 = ~n694 & ~n695;
  assign n697 = \C<16>  & ~\data<32> ;
  assign n698 = ~\C<16>  & \data<32> ;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~\data<63>  & \C<13> ;
  assign n701 = \data<63>  & ~\C<13> ;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~n699 & n702;
  assign n704 = n696 & n703;
  assign n705 = n693 & n704;
  assign n706 = ~n690 & n705;
  assign n707 = n687 & n706;
  assign n708 = n690 & n705;
  assign n709 = n687 & n708;
  assign n710 = n699 & n702;
  assign n711 = ~n696 & n710;
  assign n712 = ~n693 & n711;
  assign n713 = n690 & n712;
  assign n714 = n687 & n713;
  assign n715 = ~n699 & ~n702;
  assign n716 = ~n696 & n715;
  assign n717 = ~n693 & n716;
  assign n718 = n690 & n717;
  assign n719 = ~n687 & n718;
  assign n720 = n693 & n716;
  assign n721 = n690 & n720;
  assign n722 = ~n687 & n721;
  assign n723 = n693 & n711;
  assign n724 = ~n690 & n723;
  assign n725 = n687 & n724;
  assign n726 = n696 & n715;
  assign n727 = ~n693 & n726;
  assign n728 = ~n690 & n727;
  assign n729 = ~n687 & n728;
  assign n730 = n690 & n727;
  assign n731 = ~n687 & n730;
  assign n732 = n693 & n726;
  assign n733 = ~n690 & n732;
  assign n734 = ~n687 & n733;
  assign n735 = n699 & ~n702;
  assign n736 = ~n696 & n735;
  assign n737 = ~n693 & n736;
  assign n738 = ~n690 & n737;
  assign n739 = ~n687 & n738;
  assign n740 = n696 & n735;
  assign n741 = n693 & n740;
  assign n742 = n690 & n741;
  assign n743 = ~n687 & n742;
  assign n744 = ~n690 & n720;
  assign n745 = n687 & n744;
  assign n746 = n687 & n721;
  assign n747 = n687 & n728;
  assign n748 = n690 & n732;
  assign n749 = n687 & n748;
  assign n750 = n687 & n738;
  assign n751 = n693 & n736;
  assign n752 = ~n690 & n751;
  assign n753 = n687 & n752;
  assign n754 = ~n693 & n740;
  assign n755 = n690 & n754;
  assign n756 = n687 & n755;
  assign n757 = ~n696 & n703;
  assign n758 = ~n693 & n757;
  assign n759 = n690 & n758;
  assign n760 = ~n687 & n759;
  assign n761 = ~n693 & n704;
  assign n762 = ~n690 & n761;
  assign n763 = ~n687 & n762;
  assign n764 = ~n687 & n706;
  assign n765 = ~n687 & n708;
  assign n766 = n690 & n723;
  assign n767 = ~n687 & n766;
  assign n768 = n696 & n710;
  assign n769 = ~n693 & n768;
  assign n770 = n690 & n769;
  assign n771 = ~n687 & n770;
  assign n772 = n693 & n768;
  assign n773 = ~n690 & n772;
  assign n774 = ~n687 & n773;
  assign n775 = ~n690 & n758;
  assign n776 = n687 & n775;
  assign n777 = n690 & n761;
  assign n778 = n687 & n777;
  assign n779 = n690 & n772;
  assign n780 = n687 & n779;
  assign n781 = n687 & n766;
  assign n782 = n690 & n737;
  assign n783 = n687 & n782;
  assign n784 = ~n687 & n724;
  assign n785 = ~n778 & ~n780;
  assign n786 = ~n776 & n785;
  assign n787 = ~n774 & n786;
  assign n788 = ~n771 & n787;
  assign n789 = ~n767 & n788;
  assign n790 = ~n765 & n789;
  assign n791 = ~n764 & n790;
  assign n792 = ~n763 & n791;
  assign n793 = ~n760 & n792;
  assign n794 = ~n756 & n793;
  assign n795 = ~n753 & n794;
  assign n796 = ~n750 & n795;
  assign n797 = ~n749 & n796;
  assign n798 = ~n747 & n797;
  assign n799 = ~n746 & n798;
  assign n800 = ~n745 & n799;
  assign n801 = ~n743 & n800;
  assign n802 = ~n739 & n801;
  assign n803 = ~n734 & n802;
  assign n804 = ~n731 & n803;
  assign n805 = ~n729 & n804;
  assign n806 = ~n725 & n805;
  assign n807 = ~n722 & n806;
  assign n808 = ~n719 & n807;
  assign n809 = ~n714 & n808;
  assign n810 = ~n709 & n809;
  assign n811 = ~n707 & n810;
  assign n812 = ~n690 & n754;
  assign n813 = ~n687 & n812;
  assign n814 = n811 & ~n813;
  assign n815 = ~n784 & n814;
  assign n816 = ~n783 & n815;
  assign n817 = ~n781 & n816;
  assign n818 = \data<22>  & n504;
  assign n819 = n817 & n818;
  assign n820 = ~\data<22>  & n504;
  assign n821 = ~n817 & n820;
  assign n822 = \outreg<21>  & n510;
  assign n823 = \outreg<13>  & n508;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n821 & n824;
  assign \outreg_new<13>  = n819 | ~n825;
  assign n827 = \outreg<22>  & n510;
  assign n828 = \outreg<14>  & n508;
  assign n829 = \data<62>  & n504;
  assign n830 = ~n828 & ~n829;
  assign \outreg_new<14>  = n827 | ~n830;
  assign n832 = \inreg<34>  & n508;
  assign n833 = \inreg<26>  & n510;
  assign \inreg_new<34>  = n832 | n833;
  assign n835 = ~\count<3>  & n675;
  assign n836 = \count<2>  & n835;
  assign n837 = \count<0>  & n836;
  assign n838 = \count<1>  & n837;
  assign n839 = \count<3>  & n675;
  assign n840 = ~\count<1>  & n839;
  assign n841 = ~\count<2>  & n839;
  assign n842 = ~\count<0>  & n839;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n840 & n843;
  assign \count_new<3>  = n838 | ~n844;
  assign n846 = \inreg<33>  & n508;
  assign n847 = \inreg<25>  & n510;
  assign \inreg_new<33>  = n846 | n847;
  assign n849 = \inreg<32>  & n508;
  assign n850 = \inreg<24>  & n510;
  assign \inreg_new<32>  = n849 | n850;
  assign n852 = \count<0>  & n675;
  assign n853 = ~\count<1>  & n852;
  assign n854 = \count<1>  & \count_new<0> ;
  assign \count_new<1>  = n853 | n854;
  assign n856 = \data<51>  & ~n504;
  assign n857 = \inreg<29>  & n504;
  assign \data_new<19>  = n856 | n857;
  assign n859 = \inreg<31>  & n508;
  assign n860 = \inreg<23>  & n510;
  assign \inreg_new<31>  = n859 | n860;
  assign n862 = ~\count<2>  & n675;
  assign n863 = \count<0>  & n862;
  assign n864 = \count<1>  & n863;
  assign n865 = \count<2>  & n675;
  assign n866 = ~\count<1>  & n865;
  assign n867 = ~\count<0>  & n865;
  assign n868 = ~n866 & ~n867;
  assign \count_new<2>  = n864 | ~n868;
  assign n870 = \outreg<18>  & n510;
  assign n871 = \outreg<10>  & n508;
  assign n872 = \data<46>  & n504;
  assign n873 = ~n871 & ~n872;
  assign \outreg_new<10>  = n870 | ~n873;
  assign n875 = \inreg<38>  & n508;
  assign n876 = \inreg<30>  & n510;
  assign \inreg_new<38>  = n875 | n876;
  assign n878 = \D<26>  & ~\data<52> ;
  assign n879 = ~\D<26>  & \data<52> ;
  assign n880 = ~n878 & ~n879;
  assign n881 = \D<18>  & ~\data<51> ;
  assign n882 = ~\D<18>  & \data<51> ;
  assign n883 = ~n881 & ~n882;
  assign n884 = \D<8>  & ~\data<50> ;
  assign n885 = ~\D<8>  & \data<50> ;
  assign n886 = ~n884 & ~n885;
  assign n887 = \D<2>  & ~\data<49> ;
  assign n888 = ~\D<2>  & \data<49> ;
  assign n889 = ~n887 & ~n888;
  assign n890 = \D<23>  & ~\data<48> ;
  assign n891 = ~\D<23>  & \data<48> ;
  assign n892 = ~n890 & ~n891;
  assign n893 = \D<12>  & ~\data<47> ;
  assign n894 = ~\D<12>  & \data<47> ;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n892 & ~n895;
  assign n897 = ~n889 & n896;
  assign n898 = ~n886 & n897;
  assign n899 = n883 & n898;
  assign n900 = ~n880 & n899;
  assign n901 = n889 & n896;
  assign n902 = n886 & n901;
  assign n903 = ~n883 & n902;
  assign n904 = ~n880 & n903;
  assign n905 = n883 & n902;
  assign n906 = ~n880 & n905;
  assign n907 = n892 & ~n895;
  assign n908 = ~n889 & n907;
  assign n909 = ~n886 & n908;
  assign n910 = ~n883 & n909;
  assign n911 = ~n880 & n910;
  assign n912 = n886 & n908;
  assign n913 = ~n883 & n912;
  assign n914 = ~n880 & n913;
  assign n915 = n889 & n907;
  assign n916 = ~n886 & n915;
  assign n917 = ~n883 & n916;
  assign n918 = ~n880 & n917;
  assign n919 = n883 & n916;
  assign n920 = ~n880 & n919;
  assign n921 = ~n883 & n898;
  assign n922 = n880 & n921;
  assign n923 = n886 & n897;
  assign n924 = n883 & n923;
  assign n925 = n880 & n924;
  assign n926 = ~n886 & n901;
  assign n927 = ~n883 & n926;
  assign n928 = n880 & n927;
  assign n929 = n883 & n926;
  assign n930 = n880 & n929;
  assign n931 = n880 & n905;
  assign n932 = n883 & n909;
  assign n933 = n880 & n932;
  assign n934 = n880 & n913;
  assign n935 = ~n892 & n895;
  assign n936 = ~n889 & n935;
  assign n937 = ~n886 & n936;
  assign n938 = ~n883 & n937;
  assign n939 = ~n880 & n938;
  assign n940 = n889 & n935;
  assign n941 = ~n886 & n940;
  assign n942 = n883 & n941;
  assign n943 = ~n880 & n942;
  assign n944 = n886 & n940;
  assign n945 = n883 & n944;
  assign n946 = ~n880 & n945;
  assign n947 = n892 & n895;
  assign n948 = ~n889 & n947;
  assign n949 = ~n886 & n948;
  assign n950 = n883 & n949;
  assign n951 = ~n880 & n950;
  assign n952 = n886 & n948;
  assign n953 = ~n883 & n952;
  assign n954 = ~n880 & n953;
  assign n955 = n889 & n947;
  assign n956 = ~n886 & n955;
  assign n957 = ~n883 & n956;
  assign n958 = ~n880 & n957;
  assign n959 = n886 & n955;
  assign n960 = n883 & n959;
  assign n961 = ~n880 & n960;
  assign n962 = n883 & n937;
  assign n963 = n880 & n962;
  assign n964 = n886 & n936;
  assign n965 = n883 & n964;
  assign n966 = n880 & n965;
  assign n967 = ~n883 & n941;
  assign n968 = n880 & n967;
  assign n969 = ~n883 & n944;
  assign n970 = n880 & n969;
  assign n971 = ~n883 & n949;
  assign n972 = n880 & n971;
  assign n973 = n883 & n952;
  assign n974 = n880 & n973;
  assign n975 = ~n883 & n959;
  assign n976 = n880 & n975;
  assign n977 = n886 & n915;
  assign n978 = n883 & n977;
  assign n979 = n880 & n978;
  assign n980 = n883 & n956;
  assign n981 = n880 & n980;
  assign n982 = ~n880 & n973;
  assign n983 = ~n883 & n923;
  assign n984 = ~n880 & n983;
  assign n985 = ~n974 & ~n976;
  assign n986 = ~n972 & n985;
  assign n987 = ~n970 & n986;
  assign n988 = ~n968 & n987;
  assign n989 = ~n966 & n988;
  assign n990 = ~n963 & n989;
  assign n991 = ~n961 & n990;
  assign n992 = ~n958 & n991;
  assign n993 = ~n954 & n992;
  assign n994 = ~n951 & n993;
  assign n995 = ~n946 & n994;
  assign n996 = ~n943 & n995;
  assign n997 = ~n939 & n996;
  assign n998 = ~n934 & n997;
  assign n999 = ~n933 & n998;
  assign n1000 = ~n931 & n999;
  assign n1001 = ~n930 & n1000;
  assign n1002 = ~n928 & n1001;
  assign n1003 = ~n925 & n1002;
  assign n1004 = ~n922 & n1003;
  assign n1005 = ~n920 & n1004;
  assign n1006 = ~n918 & n1005;
  assign n1007 = ~n914 & n1006;
  assign n1008 = ~n911 & n1007;
  assign n1009 = ~n906 & n1008;
  assign n1010 = ~n904 & n1009;
  assign n1011 = ~n900 & n1010;
  assign n1012 = ~n984 & n1011;
  assign n1013 = ~n982 & n1012;
  assign n1014 = ~n981 & n1013;
  assign n1015 = ~n979 & n1014;
  assign n1016 = \data<13>  & n504;
  assign n1017 = n1015 & n1016;
  assign n1018 = ~\data<13>  & n504;
  assign n1019 = ~n1015 & n1018;
  assign n1020 = \outreg<27>  & n510;
  assign n1021 = \outreg<19>  & n508;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1019 & n1022;
  assign \outreg_new<19>  = n1017 | ~n1023;
  assign n1025 = \data<49>  & ~n504;
  assign n1026 = \inreg<45>  & n504;
  assign \data_new<17>  = n1025 | n1026;
  assign n1028 = \inreg<37>  & n508;
  assign n1029 = \inreg<29>  & n510;
  assign \inreg_new<37>  = n1028 | n1029;
  assign n1031 = \data<50>  & ~n504;
  assign n1032 = \inreg<37>  & n504;
  assign \data_new<18>  = n1031 | n1032;
  assign n1034 = \inreg<36>  & n508;
  assign n1035 = \inreg<28>  & n510;
  assign \inreg_new<36>  = n1034 | n1035;
  assign n1037 = \data<47>  & ~n504;
  assign n1038 = \data_in<3>  & n504;
  assign \data_new<15>  = n1037 | n1038;
  assign n1040 = \inreg<35>  & n508;
  assign n1041 = \inreg<27>  & n510;
  assign \inreg_new<35>  = n1040 | n1041;
  assign n1043 = \data<48>  & ~n504;
  assign n1044 = \inreg<53>  & n504;
  assign \data_new<16>  = n1043 | n1044;
  assign n1046 = ~n690 & n717;
  assign n1047 = ~n687 & n1046;
  assign n1048 = ~n687 & n748;
  assign n1049 = ~n687 & n752;
  assign n1050 = n687 & n718;
  assign n1051 = n687 & n730;
  assign n1052 = n690 & n751;
  assign n1053 = n687 & n1052;
  assign n1054 = n687 & n770;
  assign n1055 = n693 & n757;
  assign n1056 = ~n690 & n1055;
  assign n1057 = ~n687 & n1056;
  assign n1058 = n690 & n1055;
  assign n1059 = ~n687 & n1058;
  assign n1060 = ~n687 & n713;
  assign n1061 = n687 & n1056;
  assign n1062 = n687 & n1058;
  assign n1063 = ~n690 & n741;
  assign n1064 = n687 & n1063;
  assign n1065 = ~n690 & n769;
  assign n1066 = n687 & n1065;
  assign n1067 = ~n687 & n782;
  assign n1068 = ~n690 & n712;
  assign n1069 = ~n687 & n1068;
  assign n1070 = ~n1061 & ~n1062;
  assign n1071 = ~n776 & n1070;
  assign n1072 = ~n774 & n1071;
  assign n1073 = ~n771 & n1072;
  assign n1074 = ~n1060 & n1073;
  assign n1075 = ~n763 & n1074;
  assign n1076 = ~n1059 & n1075;
  assign n1077 = ~n1057 & n1076;
  assign n1078 = ~n1054 & n1077;
  assign n1079 = ~n760 & n1078;
  assign n1080 = ~n1053 & n1079;
  assign n1081 = ~n750 & n1080;
  assign n1082 = ~n749 & n1081;
  assign n1083 = ~n1051 & n1082;
  assign n1084 = ~n747 & n1083;
  assign n1085 = ~n746 & n1084;
  assign n1086 = ~n1050 & n1085;
  assign n1087 = ~n743 & n1086;
  assign n1088 = ~n1049 & n1087;
  assign n1089 = ~n739 & n1088;
  assign n1090 = ~n1048 & n1089;
  assign n1091 = ~n734 & n1090;
  assign n1092 = ~n731 & n1091;
  assign n1093 = ~n725 & n1092;
  assign n1094 = ~n1047 & n1093;
  assign n1095 = ~n714 & n1094;
  assign n1096 = ~n709 & n1095;
  assign n1097 = ~n1069 & n1096;
  assign n1098 = ~n1067 & n1097;
  assign n1099 = ~n1066 & n1098;
  assign n1100 = ~n1064 & n1099;
  assign n1101 = \data<30>  & n504;
  assign n1102 = n1100 & n1101;
  assign n1103 = ~\data<30>  & n504;
  assign n1104 = ~n1100 & n1103;
  assign n1105 = \outreg<23>  & n510;
  assign n1106 = \outreg<15>  & n508;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = ~n1104 & n1107;
  assign \outreg_new<15>  = n1102 | ~n1108;
  assign n1110 = \outreg<24>  & n510;
  assign n1111 = \outreg<16>  & n508;
  assign n1112 = \data<37>  & n504;
  assign n1113 = ~n1111 & ~n1112;
  assign \outreg_new<16>  = n1110 | ~n1113;
  assign n1115 = ~\data<44>  & \C<7> ;
  assign n1116 = \data<44>  & ~\C<7> ;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = \C<25>  & ~\data<43> ;
  assign n1119 = ~\C<25>  & \data<43> ;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~\data<42>  & \C<3> ;
  assign n1122 = \data<42>  & ~\C<3> ;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = \C<11>  & ~\data<41> ;
  assign n1125 = ~\C<11>  & \data<41> ;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = \C<18>  & ~\data<40> ;
  assign n1128 = ~\C<18>  & \data<40> ;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = \C<22>  & ~\data<39> ;
  assign n1131 = ~\C<22>  & \data<39> ;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1129 & ~n1132;
  assign n1134 = ~n1126 & n1133;
  assign n1135 = n1123 & n1134;
  assign n1136 = ~n1120 & n1135;
  assign n1137 = ~n1117 & n1136;
  assign n1138 = n1120 & n1135;
  assign n1139 = ~n1117 & n1138;
  assign n1140 = n1126 & n1133;
  assign n1141 = ~n1123 & n1140;
  assign n1142 = ~n1120 & n1141;
  assign n1143 = ~n1117 & n1142;
  assign n1144 = n1123 & n1140;
  assign n1145 = ~n1120 & n1144;
  assign n1146 = ~n1117 & n1145;
  assign n1147 = n1129 & ~n1132;
  assign n1148 = ~n1126 & n1147;
  assign n1149 = ~n1123 & n1148;
  assign n1150 = ~n1120 & n1149;
  assign n1151 = ~n1117 & n1150;
  assign n1152 = n1123 & n1148;
  assign n1153 = ~n1120 & n1152;
  assign n1154 = ~n1117 & n1153;
  assign n1155 = n1126 & n1147;
  assign n1156 = ~n1123 & n1155;
  assign n1157 = n1120 & n1156;
  assign n1158 = ~n1117 & n1157;
  assign n1159 = ~n1123 & n1134;
  assign n1160 = ~n1120 & n1159;
  assign n1161 = n1117 & n1160;
  assign n1162 = n1117 & n1138;
  assign n1163 = n1120 & n1144;
  assign n1164 = n1117 & n1163;
  assign n1165 = n1120 & n1149;
  assign n1166 = n1117 & n1165;
  assign n1167 = n1117 & n1153;
  assign n1168 = ~n1120 & n1156;
  assign n1169 = n1117 & n1168;
  assign n1170 = n1123 & n1155;
  assign n1171 = n1120 & n1170;
  assign n1172 = n1117 & n1171;
  assign n1173 = ~n1129 & n1132;
  assign n1174 = ~n1126 & n1173;
  assign n1175 = ~n1123 & n1174;
  assign n1176 = n1120 & n1175;
  assign n1177 = ~n1117 & n1176;
  assign n1178 = n1123 & n1174;
  assign n1179 = ~n1120 & n1178;
  assign n1180 = ~n1117 & n1179;
  assign n1181 = n1126 & n1173;
  assign n1182 = ~n1123 & n1181;
  assign n1183 = n1120 & n1182;
  assign n1184 = ~n1117 & n1183;
  assign n1185 = n1129 & n1132;
  assign n1186 = ~n1126 & n1185;
  assign n1187 = n1123 & n1186;
  assign n1188 = n1120 & n1187;
  assign n1189 = ~n1117 & n1188;
  assign n1190 = n1126 & n1185;
  assign n1191 = ~n1123 & n1190;
  assign n1192 = ~n1120 & n1191;
  assign n1193 = ~n1117 & n1192;
  assign n1194 = n1123 & n1190;
  assign n1195 = ~n1120 & n1194;
  assign n1196 = ~n1117 & n1195;
  assign n1197 = n1120 & n1194;
  assign n1198 = ~n1117 & n1197;
  assign n1199 = n1120 & n1178;
  assign n1200 = n1117 & n1199;
  assign n1201 = ~n1120 & n1182;
  assign n1202 = n1117 & n1201;
  assign n1203 = n1123 & n1181;
  assign n1204 = ~n1120 & n1203;
  assign n1205 = n1117 & n1204;
  assign n1206 = ~n1123 & n1186;
  assign n1207 = ~n1120 & n1206;
  assign n1208 = n1117 & n1207;
  assign n1209 = n1120 & n1206;
  assign n1210 = n1117 & n1209;
  assign n1211 = ~n1120 & n1187;
  assign n1212 = n1117 & n1211;
  assign n1213 = n1120 & n1191;
  assign n1214 = n1117 & n1213;
  assign n1215 = n1120 & n1203;
  assign n1216 = n1117 & n1215;
  assign n1217 = n1117 & n1145;
  assign n1218 = ~n1117 & n1171;
  assign n1219 = ~n1212 & ~n1214;
  assign n1220 = ~n1210 & n1219;
  assign n1221 = ~n1208 & n1220;
  assign n1222 = ~n1205 & n1221;
  assign n1223 = ~n1202 & n1222;
  assign n1224 = ~n1200 & n1223;
  assign n1225 = ~n1198 & n1224;
  assign n1226 = ~n1196 & n1225;
  assign n1227 = ~n1193 & n1226;
  assign n1228 = ~n1189 & n1227;
  assign n1229 = ~n1184 & n1228;
  assign n1230 = ~n1180 & n1229;
  assign n1231 = ~n1177 & n1230;
  assign n1232 = ~n1172 & n1231;
  assign n1233 = ~n1169 & n1232;
  assign n1234 = ~n1167 & n1233;
  assign n1235 = ~n1166 & n1234;
  assign n1236 = ~n1164 & n1235;
  assign n1237 = ~n1162 & n1236;
  assign n1238 = ~n1161 & n1237;
  assign n1239 = ~n1158 & n1238;
  assign n1240 = ~n1154 & n1239;
  assign n1241 = ~n1151 & n1240;
  assign n1242 = ~n1146 & n1241;
  assign n1243 = ~n1143 & n1242;
  assign n1244 = ~n1139 & n1243;
  assign n1245 = ~n1137 & n1244;
  assign n1246 = ~n1120 & n1175;
  assign n1247 = ~n1117 & n1246;
  assign n1248 = n1245 & ~n1247;
  assign n1249 = ~n1218 & n1248;
  assign n1250 = ~n1217 & n1249;
  assign n1251 = ~n1216 & n1250;
  assign n1252 = \data<5>  & n504;
  assign n1253 = n1251 & n1252;
  assign n1254 = ~\data<5>  & n504;
  assign n1255 = ~n1251 & n1254;
  assign n1256 = \outreg<25>  & n510;
  assign n1257 = \outreg<17>  & n508;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n1255 & n1258;
  assign \outreg_new<17>  = n1253 | ~n1259;
  assign n1261 = \inreg<39>  & n508;
  assign n1262 = \inreg<31>  & n510;
  assign \inreg_new<39>  = n1261 | n1262;
  assign n1264 = \outreg<26>  & n510;
  assign n1265 = \outreg<18>  & n508;
  assign n1266 = \data<45>  & n504;
  assign n1267 = ~n1265 & ~n1266;
  assign \outreg_new<18>  = n1264 | ~n1267;
  assign n1269 = \D<24>  & ~\data<60> ;
  assign n1270 = ~\D<24>  & \data<60> ;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = \D<5>  & ~\data<59> ;
  assign n1273 = ~\D<5>  & \data<59> ;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = \D<27>  & ~\data<58> ;
  assign n1276 = ~\D<27>  & \data<58> ;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = \D<10>  & ~\data<57> ;
  assign n1279 = ~\D<10>  & \data<57> ;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = \D<20>  & ~\data<56> ;
  assign n1282 = ~\D<20>  & \data<56> ;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = \D<15>  & ~\data<55> ;
  assign n1285 = ~\D<15>  & \data<55> ;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1283 & ~n1286;
  assign n1288 = ~n1280 & n1287;
  assign n1289 = ~n1277 & n1288;
  assign n1290 = n1274 & n1289;
  assign n1291 = ~n1271 & n1290;
  assign n1292 = n1277 & n1288;
  assign n1293 = n1274 & n1292;
  assign n1294 = ~n1271 & n1293;
  assign n1295 = n1280 & n1287;
  assign n1296 = ~n1277 & n1295;
  assign n1297 = ~n1274 & n1296;
  assign n1298 = ~n1271 & n1297;
  assign n1299 = n1283 & ~n1286;
  assign n1300 = ~n1280 & n1299;
  assign n1301 = ~n1277 & n1300;
  assign n1302 = ~n1274 & n1301;
  assign n1303 = ~n1271 & n1302;
  assign n1304 = n1274 & n1301;
  assign n1305 = ~n1271 & n1304;
  assign n1306 = n1280 & n1299;
  assign n1307 = n1277 & n1306;
  assign n1308 = ~n1274 & n1307;
  assign n1309 = ~n1271 & n1308;
  assign n1310 = n1274 & n1307;
  assign n1311 = ~n1271 & n1310;
  assign n1312 = n1274 & n1296;
  assign n1313 = n1271 & n1312;
  assign n1314 = n1277 & n1295;
  assign n1315 = ~n1274 & n1314;
  assign n1316 = n1271 & n1315;
  assign n1317 = n1274 & n1314;
  assign n1318 = n1271 & n1317;
  assign n1319 = n1271 & n1302;
  assign n1320 = n1271 & n1304;
  assign n1321 = n1277 & n1300;
  assign n1322 = ~n1274 & n1321;
  assign n1323 = n1271 & n1322;
  assign n1324 = ~n1277 & n1306;
  assign n1325 = n1274 & n1324;
  assign n1326 = n1271 & n1325;
  assign n1327 = ~n1283 & n1286;
  assign n1328 = ~n1280 & n1327;
  assign n1329 = ~n1277 & n1328;
  assign n1330 = ~n1274 & n1329;
  assign n1331 = ~n1271 & n1330;
  assign n1332 = n1277 & n1328;
  assign n1333 = ~n1274 & n1332;
  assign n1334 = ~n1271 & n1333;
  assign n1335 = n1280 & n1327;
  assign n1336 = n1277 & n1335;
  assign n1337 = ~n1274 & n1336;
  assign n1338 = ~n1271 & n1337;
  assign n1339 = n1274 & n1336;
  assign n1340 = ~n1271 & n1339;
  assign n1341 = n1283 & n1286;
  assign n1342 = ~n1280 & n1341;
  assign n1343 = ~n1277 & n1342;
  assign n1344 = ~n1274 & n1343;
  assign n1345 = ~n1271 & n1344;
  assign n1346 = n1280 & n1341;
  assign n1347 = ~n1277 & n1346;
  assign n1348 = ~n1274 & n1347;
  assign n1349 = ~n1271 & n1348;
  assign n1350 = n1274 & n1347;
  assign n1351 = ~n1271 & n1350;
  assign n1352 = n1274 & n1329;
  assign n1353 = n1271 & n1352;
  assign n1354 = n1271 & n1333;
  assign n1355 = ~n1277 & n1335;
  assign n1356 = ~n1274 & n1355;
  assign n1357 = n1271 & n1356;
  assign n1358 = n1271 & n1339;
  assign n1359 = n1277 & n1342;
  assign n1360 = n1274 & n1359;
  assign n1361 = n1271 & n1360;
  assign n1362 = n1271 & n1348;
  assign n1363 = n1277 & n1346;
  assign n1364 = ~n1274 & n1363;
  assign n1365 = n1271 & n1364;
  assign n1366 = n1271 & n1350;
  assign n1367 = ~n1274 & n1289;
  assign n1368 = n1271 & n1367;
  assign n1369 = ~n1274 & n1292;
  assign n1370 = ~n1271 & n1369;
  assign n1371 = ~n1362 & ~n1365;
  assign n1372 = ~n1361 & n1371;
  assign n1373 = ~n1358 & n1372;
  assign n1374 = ~n1357 & n1373;
  assign n1375 = ~n1354 & n1374;
  assign n1376 = ~n1353 & n1375;
  assign n1377 = ~n1351 & n1376;
  assign n1378 = ~n1349 & n1377;
  assign n1379 = ~n1345 & n1378;
  assign n1380 = ~n1340 & n1379;
  assign n1381 = ~n1338 & n1380;
  assign n1382 = ~n1334 & n1381;
  assign n1383 = ~n1331 & n1382;
  assign n1384 = ~n1326 & n1383;
  assign n1385 = ~n1323 & n1384;
  assign n1386 = ~n1320 & n1385;
  assign n1387 = ~n1319 & n1386;
  assign n1388 = ~n1318 & n1387;
  assign n1389 = ~n1316 & n1388;
  assign n1390 = ~n1313 & n1389;
  assign n1391 = ~n1311 & n1390;
  assign n1392 = ~n1309 & n1391;
  assign n1393 = ~n1305 & n1392;
  assign n1394 = ~n1303 & n1393;
  assign n1395 = ~n1298 & n1394;
  assign n1396 = ~n1294 & n1395;
  assign n1397 = ~n1291 & n1396;
  assign n1398 = ~n1370 & n1397;
  assign n1399 = n1274 & n1332;
  assign n1400 = ~n1271 & n1399;
  assign n1401 = n1398 & ~n1400;
  assign n1402 = ~n1368 & n1401;
  assign n1403 = ~n1366 & n1402;
  assign n1404 = \data<21>  & n504;
  assign n1405 = n1403 & n1404;
  assign n1406 = ~\data<21>  & n504;
  assign n1407 = ~n1403 & n1406;
  assign n1408 = \outreg<29>  & n510;
  assign n1409 = \outreg<21>  & n508;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1407 & n1410;
  assign \outreg_new<21>  = n1405 | ~n1411;
  assign n1413 = \outreg<30>  & n510;
  assign n1414 = \outreg<22>  & n508;
  assign n1415 = \data<61>  & n504;
  assign n1416 = ~n1414 & ~n1415;
  assign \outreg_new<22>  = n1413 | ~n1416;
  assign n1418 = n1120 & n1141;
  assign n1419 = ~n1117 & n1418;
  assign n1420 = n1120 & n1152;
  assign n1421 = ~n1117 & n1420;
  assign n1422 = ~n1120 & n1170;
  assign n1423 = ~n1117 & n1422;
  assign n1424 = n1120 & n1159;
  assign n1425 = n1117 & n1424;
  assign n1426 = n1117 & n1136;
  assign n1427 = n1117 & n1422;
  assign n1428 = ~n1117 & n1201;
  assign n1429 = ~n1117 & n1207;
  assign n1430 = ~n1117 & n1209;
  assign n1431 = n1117 & n1188;
  assign n1432 = n1117 & n1192;
  assign n1433 = n1117 & n1197;
  assign n1434 = n1117 & n1418;
  assign n1435 = n1117 & n1176;
  assign n1436 = ~n1117 & n1215;
  assign n1437 = ~n1432 & ~n1433;
  assign n1438 = ~n1431 & n1437;
  assign n1439 = ~n1212 & n1438;
  assign n1440 = ~n1210 & n1439;
  assign n1441 = ~n1202 & n1440;
  assign n1442 = ~n1200 & n1441;
  assign n1443 = ~n1196 & n1442;
  assign n1444 = ~n1189 & n1443;
  assign n1445 = ~n1430 & n1444;
  assign n1446 = ~n1429 & n1445;
  assign n1447 = ~n1428 & n1446;
  assign n1448 = ~n1180 & n1447;
  assign n1449 = ~n1177 & n1448;
  assign n1450 = ~n1427 & n1449;
  assign n1451 = ~n1167 & n1450;
  assign n1452 = ~n1166 & n1451;
  assign n1453 = ~n1164 & n1452;
  assign n1454 = ~n1426 & n1453;
  assign n1455 = ~n1425 & n1454;
  assign n1456 = ~n1161 & n1455;
  assign n1457 = ~n1423 & n1456;
  assign n1458 = ~n1421 & n1457;
  assign n1459 = ~n1151 & n1458;
  assign n1460 = ~n1146 & n1459;
  assign n1461 = ~n1419 & n1460;
  assign n1462 = ~n1143 & n1461;
  assign n1463 = ~n1139 & n1462;
  assign n1464 = ~n1117 & n1424;
  assign n1465 = n1463 & ~n1464;
  assign n1466 = ~n1436 & n1465;
  assign n1467 = ~n1435 & n1466;
  assign n1468 = ~n1434 & n1467;
  assign n1469 = \data<29>  & n504;
  assign n1470 = n1468 & n1469;
  assign n1471 = ~\data<29>  & n504;
  assign n1472 = ~n1468 & n1471;
  assign n1473 = \outreg<31>  & n510;
  assign n1474 = \outreg<23>  & n508;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n1472 & n1475;
  assign \outreg_new<23>  = n1470 | ~n1476;
  assign n1478 = \outreg<32>  & n510;
  assign n1479 = \outreg<24>  & n508;
  assign n1480 = \data<36>  & n504;
  assign n1481 = ~n1479 & ~n1480;
  assign \outreg_new<24>  = n1478 | ~n1481;
  assign n1483 = \outreg<28>  & n510;
  assign n1484 = \outreg<20>  & n508;
  assign n1485 = \data<53>  & n504;
  assign n1486 = ~n1484 & ~n1485;
  assign \outreg_new<20>  = n1483 | ~n1486;
  assign n1488 = ~n536 & n577;
  assign n1489 = ~n536 & n581;
  assign n1490 = ~n536 & n630;
  assign n1491 = n536 & n557;
  assign n1492 = ~n539 & n580;
  assign n1493 = n536 & n1492;
  assign n1494 = n539 & n568;
  assign n1495 = n536 & n1494;
  assign n1496 = n539 & n618;
  assign n1497 = ~n536 & n1496;
  assign n1498 = ~n539 & n623;
  assign n1499 = ~n536 & n1498;
  assign n1500 = ~n542 & n614;
  assign n1501 = n539 & n1500;
  assign n1502 = ~n536 & n1501;
  assign n1503 = n539 & n595;
  assign n1504 = n536 & n1503;
  assign n1505 = n536 & n1498;
  assign n1506 = n539 & n615;
  assign n1507 = n536 & n1506;
  assign n1508 = n536 & n573;
  assign n1509 = ~n539 & n606;
  assign n1510 = n536 & n1509;
  assign n1511 = ~n536 & n1506;
  assign n1512 = ~n627 & ~n1507;
  assign n1513 = ~n626 & n1512;
  assign n1514 = ~n1505 & n1513;
  assign n1515 = ~n622 & n1514;
  assign n1516 = ~n1504 & n1515;
  assign n1517 = ~n620 & n1516;
  assign n1518 = ~n617 & n1517;
  assign n1519 = ~n1502 & n1518;
  assign n1520 = ~n611 & n1519;
  assign n1521 = ~n608 & n1520;
  assign n1522 = ~n1499 & n1521;
  assign n1523 = ~n601 & n1522;
  assign n1524 = ~n1497 & n1523;
  assign n1525 = ~n592 & n1524;
  assign n1526 = ~n590 & n1525;
  assign n1527 = ~n1495 & n1526;
  assign n1528 = ~n1493 & n1527;
  assign n1529 = ~n579 & n1528;
  assign n1530 = ~n578 & n1529;
  assign n1531 = ~n1491 & n1530;
  assign n1532 = ~n574 & n1531;
  assign n1533 = ~n1490 & n1532;
  assign n1534 = ~n565 & n1533;
  assign n1535 = ~n1489 & n1534;
  assign n1536 = ~n561 & n1535;
  assign n1537 = ~n1488 & n1536;
  assign n1538 = ~n556 & n1537;
  assign n1539 = ~n536 & n589;
  assign n1540 = n1538 & ~n1539;
  assign n1541 = ~n1511 & n1540;
  assign n1542 = ~n1510 & n1541;
  assign n1543 = ~n1508 & n1542;
  assign n1544 = \data<20>  & n504;
  assign n1545 = n1543 & n1544;
  assign n1546 = ~\data<20>  & n504;
  assign n1547 = ~n1543 & n1546;
  assign n1548 = \outreg<37>  & n510;
  assign n1549 = \outreg<29>  & n508;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~n1547 & n1550;
  assign \outreg_new<29>  = n1545 | ~n1551;
  assign n1553 = ~n536 & n583;
  assign n1554 = n536 & n569;
  assign n1555 = ~n536 & n624;
  assign n1556 = n536 & n1496;
  assign n1557 = n536 & n1501;
  assign n1558 = n536 & n555;
  assign n1559 = ~n536 & n586;
  assign n1560 = ~n539 & n1500;
  assign n1561 = ~n536 & n1560;
  assign n1562 = ~n625 & n1513;
  assign n1563 = ~n1505 & n1562;
  assign n1564 = ~n621 & n1563;
  assign n1565 = ~n1556 & n1564;
  assign n1566 = ~n617 & n1565;
  assign n1567 = ~n1502 & n1566;
  assign n1568 = ~n613 & n1567;
  assign n1569 = ~n1555 & n1568;
  assign n1570 = ~n601 & n1569;
  assign n1571 = ~n597 & n1570;
  assign n1572 = ~n1497 & n1571;
  assign n1573 = ~n590 & n1572;
  assign n1574 = ~n1495 & n1573;
  assign n1575 = ~n1554 & n1574;
  assign n1576 = ~n587 & n1575;
  assign n1577 = ~n582 & n1576;
  assign n1578 = ~n1493 & n1577;
  assign n1579 = ~n579 & n1578;
  assign n1580 = ~n576 & n1579;
  assign n1581 = ~n570 & n1580;
  assign n1582 = ~n1490 & n1581;
  assign n1583 = ~n565 & n1582;
  assign n1584 = ~n1553 & n1583;
  assign n1585 = ~n1489 & n1584;
  assign n1586 = ~n556 & n1585;
  assign n1587 = ~n1561 & n1586;
  assign n1588 = ~n1559 & n1587;
  assign n1589 = ~n1558 & n1588;
  assign n1590 = ~n1557 & n1589;
  assign n1591 = \data<4>  & n504;
  assign n1592 = n1590 & n1591;
  assign n1593 = ~\data<4>  & n504;
  assign n1594 = ~n1590 & n1593;
  assign n1595 = \outreg<33>  & n510;
  assign n1596 = \outreg<25>  & n508;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1594 & n1597;
  assign \outreg_new<25>  = n1592 | ~n1598;
  assign n1600 = \outreg<34>  & n510;
  assign n1601 = \outreg<26>  & n508;
  assign n1602 = \data<44>  & n504;
  assign n1603 = ~n1601 & ~n1602;
  assign \outreg_new<26>  = n1600 | ~n1603;
  assign n1605 = ~\data<38>  & \C<5> ;
  assign n1606 = \data<38>  & ~\C<5> ;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = \C<14>  & ~\data<37> ;
  assign n1609 = ~\C<14>  & \data<37> ;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = \C<27>  & ~\data<36> ;
  assign n1612 = ~\C<27>  & \data<36> ;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = ~\data<35>  & \C<2> ;
  assign n1615 = \data<35>  & ~\C<2> ;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~\data<40>  & \C<9> ;
  assign n1618 = \data<40>  & ~\C<9> ;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = \C<20>  & ~\data<39> ;
  assign n1621 = ~\C<20>  & \data<39> ;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = n1619 & ~n1622;
  assign n1624 = ~n1616 & n1623;
  assign n1625 = n1613 & n1624;
  assign n1626 = n1610 & n1625;
  assign n1627 = n1607 & n1626;
  assign n1628 = ~n1619 & n1622;
  assign n1629 = n1616 & n1628;
  assign n1630 = ~n1613 & n1629;
  assign n1631 = ~n1610 & n1630;
  assign n1632 = ~n1607 & n1631;
  assign n1633 = ~n1619 & ~n1622;
  assign n1634 = n1616 & n1633;
  assign n1635 = ~n1613 & n1634;
  assign n1636 = ~n1610 & n1635;
  assign n1637 = n1607 & n1636;
  assign n1638 = n1610 & n1635;
  assign n1639 = ~n1607 & n1638;
  assign n1640 = n1610 & n1630;
  assign n1641 = n1607 & n1640;
  assign n1642 = n1613 & n1634;
  assign n1643 = ~n1610 & n1642;
  assign n1644 = ~n1607 & n1643;
  assign n1645 = n1613 & n1629;
  assign n1646 = ~n1610 & n1645;
  assign n1647 = n1607 & n1646;
  assign n1648 = n1610 & n1642;
  assign n1649 = n1607 & n1648;
  assign n1650 = n1616 & n1623;
  assign n1651 = ~n1613 & n1650;
  assign n1652 = ~n1610 & n1651;
  assign n1653 = ~n1607 & n1652;
  assign n1654 = n1619 & n1622;
  assign n1655 = n1616 & n1654;
  assign n1656 = ~n1613 & n1655;
  assign n1657 = ~n1610 & n1656;
  assign n1658 = n1607 & n1657;
  assign n1659 = n1610 & n1651;
  assign n1660 = ~n1607 & n1659;
  assign n1661 = n1610 & n1656;
  assign n1662 = n1607 & n1661;
  assign n1663 = n1613 & n1650;
  assign n1664 = ~n1610 & n1663;
  assign n1665 = n1607 & n1664;
  assign n1666 = n1610 & n1663;
  assign n1667 = ~n1607 & n1666;
  assign n1668 = n1613 & n1655;
  assign n1669 = n1610 & n1668;
  assign n1670 = n1607 & n1669;
  assign n1671 = ~n1616 & n1633;
  assign n1672 = ~n1613 & n1671;
  assign n1673 = ~n1610 & n1672;
  assign n1674 = ~n1607 & n1673;
  assign n1675 = ~n1616 & n1628;
  assign n1676 = ~n1613 & n1675;
  assign n1677 = ~n1610 & n1676;
  assign n1678 = ~n1607 & n1677;
  assign n1679 = n1610 & n1672;
  assign n1680 = ~n1607 & n1679;
  assign n1681 = n1610 & n1676;
  assign n1682 = n1607 & n1681;
  assign n1683 = n1613 & n1671;
  assign n1684 = ~n1610 & n1683;
  assign n1685 = n1607 & n1684;
  assign n1686 = n1613 & n1675;
  assign n1687 = n1610 & n1686;
  assign n1688 = ~n1607 & n1687;
  assign n1689 = n1607 & n1687;
  assign n1690 = ~n1613 & n1624;
  assign n1691 = ~n1610 & n1690;
  assign n1692 = ~n1607 & n1691;
  assign n1693 = ~n1616 & n1654;
  assign n1694 = ~n1613 & n1693;
  assign n1695 = ~n1610 & n1694;
  assign n1696 = n1607 & n1695;
  assign n1697 = n1610 & n1694;
  assign n1698 = ~n1607 & n1697;
  assign n1699 = n1613 & n1693;
  assign n1700 = ~n1610 & n1699;
  assign n1701 = ~n1607 & n1700;
  assign n1702 = n1607 & n1700;
  assign n1703 = ~n1607 & n1626;
  assign n1704 = n1610 & n1683;
  assign n1705 = n1607 & n1704;
  assign n1706 = n1610 & n1690;
  assign n1707 = n1607 & n1706;
  assign n1708 = ~n1607 & n1669;
  assign n1709 = ~n1702 & ~n1703;
  assign n1710 = ~n1701 & n1709;
  assign n1711 = ~n1698 & n1710;
  assign n1712 = ~n1696 & n1711;
  assign n1713 = ~n1692 & n1712;
  assign n1714 = ~n1689 & n1713;
  assign n1715 = ~n1688 & n1714;
  assign n1716 = ~n1685 & n1715;
  assign n1717 = ~n1682 & n1716;
  assign n1718 = ~n1680 & n1717;
  assign n1719 = ~n1678 & n1718;
  assign n1720 = ~n1674 & n1719;
  assign n1721 = ~n1670 & n1720;
  assign n1722 = ~n1667 & n1721;
  assign n1723 = ~n1665 & n1722;
  assign n1724 = ~n1662 & n1723;
  assign n1725 = ~n1660 & n1724;
  assign n1726 = ~n1658 & n1725;
  assign n1727 = ~n1653 & n1726;
  assign n1728 = ~n1649 & n1727;
  assign n1729 = ~n1647 & n1728;
  assign n1730 = ~n1644 & n1729;
  assign n1731 = ~n1641 & n1730;
  assign n1732 = ~n1639 & n1731;
  assign n1733 = ~n1637 & n1732;
  assign n1734 = ~n1632 & n1733;
  assign n1735 = ~n1627 & n1734;
  assign n1736 = ~n1607 & n1646;
  assign n1737 = n1735 & ~n1736;
  assign n1738 = ~n1708 & n1737;
  assign n1739 = ~n1707 & n1738;
  assign n1740 = ~n1705 & n1739;
  assign n1741 = \data<12>  & n504;
  assign n1742 = n1740 & n1741;
  assign n1743 = ~\data<12>  & n504;
  assign n1744 = ~n1740 & n1743;
  assign n1745 = \outreg<35>  & n510;
  assign n1746 = \outreg<27>  & n508;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n1744 & n1747;
  assign \outreg_new<27>  = n1742 | ~n1748;
  assign n1750 = \outreg<36>  & n510;
  assign n1751 = \outreg<28>  & n508;
  assign n1752 = \data<52>  & n504;
  assign n1753 = ~n1751 & ~n1752;
  assign \outreg_new<28>  = n1750 | ~n1753;
  assign n1755 = \D<19>  & ~\data<56> ;
  assign n1756 = ~\D<19>  & \data<56> ;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = \D<4>  & ~\data<55> ;
  assign n1759 = ~\D<4>  & \data<55> ;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = \D<16>  & ~\data<54> ;
  assign n1762 = ~\D<16>  & \data<54> ;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = \D<22>  & ~\data<53> ;
  assign n1765 = ~\D<22>  & \data<53> ;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = \D<11>  & ~\data<52> ;
  assign n1768 = ~\D<11>  & \data<52> ;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = \D<1>  & ~\data<51> ;
  assign n1771 = ~\D<1>  & \data<51> ;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = ~n1769 & ~n1772;
  assign n1774 = ~n1766 & n1773;
  assign n1775 = ~n1763 & n1774;
  assign n1776 = ~n1760 & n1775;
  assign n1777 = ~n1757 & n1776;
  assign n1778 = n1763 & n1774;
  assign n1779 = n1760 & n1778;
  assign n1780 = ~n1757 & n1779;
  assign n1781 = n1766 & n1773;
  assign n1782 = ~n1763 & n1781;
  assign n1783 = ~n1760 & n1782;
  assign n1784 = ~n1757 & n1783;
  assign n1785 = n1763 & n1781;
  assign n1786 = ~n1760 & n1785;
  assign n1787 = ~n1757 & n1786;
  assign n1788 = n1769 & ~n1772;
  assign n1789 = ~n1766 & n1788;
  assign n1790 = ~n1763 & n1789;
  assign n1791 = n1760 & n1790;
  assign n1792 = ~n1757 & n1791;
  assign n1793 = n1763 & n1789;
  assign n1794 = ~n1760 & n1793;
  assign n1795 = ~n1757 & n1794;
  assign n1796 = n1766 & n1788;
  assign n1797 = ~n1763 & n1796;
  assign n1798 = ~n1760 & n1797;
  assign n1799 = ~n1757 & n1798;
  assign n1800 = n1757 & n1776;
  assign n1801 = ~n1760 & n1778;
  assign n1802 = n1757 & n1801;
  assign n1803 = n1760 & n1785;
  assign n1804 = n1757 & n1803;
  assign n1805 = n1757 & n1791;
  assign n1806 = n1757 & n1798;
  assign n1807 = n1760 & n1797;
  assign n1808 = n1757 & n1807;
  assign n1809 = n1763 & n1796;
  assign n1810 = ~n1760 & n1809;
  assign n1811 = n1757 & n1810;
  assign n1812 = ~n1769 & n1772;
  assign n1813 = n1766 & n1812;
  assign n1814 = ~n1763 & n1813;
  assign n1815 = ~n1760 & n1814;
  assign n1816 = ~n1757 & n1815;
  assign n1817 = n1760 & n1814;
  assign n1818 = ~n1757 & n1817;
  assign n1819 = n1763 & n1813;
  assign n1820 = n1760 & n1819;
  assign n1821 = ~n1757 & n1820;
  assign n1822 = n1769 & n1772;
  assign n1823 = ~n1766 & n1822;
  assign n1824 = ~n1763 & n1823;
  assign n1825 = ~n1760 & n1824;
  assign n1826 = ~n1757 & n1825;
  assign n1827 = n1763 & n1823;
  assign n1828 = ~n1760 & n1827;
  assign n1829 = ~n1757 & n1828;
  assign n1830 = n1760 & n1827;
  assign n1831 = ~n1757 & n1830;
  assign n1832 = n1766 & n1822;
  assign n1833 = n1763 & n1832;
  assign n1834 = ~n1760 & n1833;
  assign n1835 = ~n1757 & n1834;
  assign n1836 = ~n1766 & n1812;
  assign n1837 = ~n1763 & n1836;
  assign n1838 = n1760 & n1837;
  assign n1839 = n1757 & n1838;
  assign n1840 = n1763 & n1836;
  assign n1841 = ~n1760 & n1840;
  assign n1842 = n1757 & n1841;
  assign n1843 = n1760 & n1840;
  assign n1844 = n1757 & n1843;
  assign n1845 = ~n1760 & n1819;
  assign n1846 = n1757 & n1845;
  assign n1847 = n1760 & n1824;
  assign n1848 = n1757 & n1847;
  assign n1849 = ~n1763 & n1832;
  assign n1850 = ~n1760 & n1849;
  assign n1851 = n1757 & n1850;
  assign n1852 = n1760 & n1833;
  assign n1853 = n1757 & n1852;
  assign n1854 = n1760 & n1782;
  assign n1855 = n1757 & n1854;
  assign n1856 = n1757 & n1815;
  assign n1857 = n1760 & n1809;
  assign n1858 = ~n1757 & n1857;
  assign n1859 = ~n1851 & ~n1853;
  assign n1860 = ~n1848 & n1859;
  assign n1861 = ~n1846 & n1860;
  assign n1862 = ~n1844 & n1861;
  assign n1863 = ~n1842 & n1862;
  assign n1864 = ~n1839 & n1863;
  assign n1865 = ~n1835 & n1864;
  assign n1866 = ~n1831 & n1865;
  assign n1867 = ~n1829 & n1866;
  assign n1868 = ~n1826 & n1867;
  assign n1869 = ~n1821 & n1868;
  assign n1870 = ~n1818 & n1869;
  assign n1871 = ~n1816 & n1870;
  assign n1872 = ~n1811 & n1871;
  assign n1873 = ~n1808 & n1872;
  assign n1874 = ~n1806 & n1873;
  assign n1875 = ~n1805 & n1874;
  assign n1876 = ~n1804 & n1875;
  assign n1877 = ~n1802 & n1876;
  assign n1878 = ~n1800 & n1877;
  assign n1879 = ~n1799 & n1878;
  assign n1880 = ~n1795 & n1879;
  assign n1881 = ~n1792 & n1880;
  assign n1882 = ~n1787 & n1881;
  assign n1883 = ~n1784 & n1882;
  assign n1884 = ~n1780 & n1883;
  assign n1885 = ~n1777 & n1884;
  assign n1886 = n1760 & n1849;
  assign n1887 = ~n1757 & n1886;
  assign n1888 = n1885 & ~n1887;
  assign n1889 = ~n1858 & n1888;
  assign n1890 = ~n1856 & n1889;
  assign n1891 = ~n1855 & n1890;
  assign n1892 = \data<28>  & n504;
  assign n1893 = n1891 & n1892;
  assign n1894 = ~\data<28>  & n504;
  assign n1895 = ~n1891 & n1894;
  assign n1896 = \outreg<39>  & n510;
  assign n1897 = \outreg<31>  & n508;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1895 & n1898;
  assign \outreg_new<31>  = n1893 | ~n1899;
  assign n1901 = \outreg<40>  & n510;
  assign n1902 = \outreg<32>  & n508;
  assign n1903 = \data<35>  & n504;
  assign n1904 = ~n1902 & ~n1903;
  assign \outreg_new<32>  = n1901 | ~n1904;
  assign n1906 = ~n1757 & n1803;
  assign n1907 = ~n1760 & n1790;
  assign n1908 = ~n1757 & n1907;
  assign n1909 = n1760 & n1793;
  assign n1910 = ~n1757 & n1909;
  assign n1911 = n1760 & n1775;
  assign n1912 = n1757 & n1911;
  assign n1913 = n1757 & n1783;
  assign n1914 = n1757 & n1857;
  assign n1915 = ~n1757 & n1841;
  assign n1916 = ~n1757 & n1847;
  assign n1917 = ~n1757 & n1852;
  assign n1918 = ~n1760 & n1837;
  assign n1919 = n1757 & n1918;
  assign n1920 = n1757 & n1830;
  assign n1921 = n1757 & n1886;
  assign n1922 = n1757 & n1794;
  assign n1923 = n1757 & n1825;
  assign n1924 = ~n1757 & n1911;
  assign n1925 = ~n1853 & ~n1921;
  assign n1926 = ~n1851 & n1925;
  assign n1927 = ~n1920 & n1926;
  assign n1928 = ~n1846 & n1927;
  assign n1929 = ~n1844 & n1928;
  assign n1930 = ~n1919 & n1929;
  assign n1931 = ~n1917 & n1930;
  assign n1932 = ~n1835 & n1931;
  assign n1933 = ~n1829 & n1932;
  assign n1934 = ~n1916 & n1933;
  assign n1935 = ~n1818 & n1934;
  assign n1936 = ~n1816 & n1935;
  assign n1937 = ~n1915 & n1936;
  assign n1938 = ~n1914 & n1937;
  assign n1939 = ~n1811 & n1938;
  assign n1940 = ~n1808 & n1939;
  assign n1941 = ~n1805 & n1940;
  assign n1942 = ~n1913 & n1941;
  assign n1943 = ~n1802 & n1942;
  assign n1944 = ~n1912 & n1943;
  assign n1945 = ~n1799 & n1944;
  assign n1946 = ~n1910 & n1945;
  assign n1947 = ~n1792 & n1946;
  assign n1948 = ~n1908 & n1947;
  assign n1949 = ~n1906 & n1948;
  assign n1950 = ~n1787 & n1949;
  assign n1951 = ~n1777 & n1950;
  assign n1952 = ~n1757 & n1918;
  assign n1953 = n1951 & ~n1952;
  assign n1954 = ~n1924 & n1953;
  assign n1955 = ~n1923 & n1954;
  assign n1956 = ~n1922 & n1955;
  assign n1957 = \data<3>  & n504;
  assign n1958 = n1956 & n1957;
  assign n1959 = ~\data<3>  & n504;
  assign n1960 = ~n1956 & n1959;
  assign n1961 = \outreg<41>  & n510;
  assign n1962 = \outreg<33>  & n508;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~n1960 & n1963;
  assign \outreg_new<33>  = n1958 | ~n1964;
  assign n1966 = \outreg<42>  & n510;
  assign n1967 = \outreg<34>  & n508;
  assign n1968 = \data<43>  & n504;
  assign n1969 = ~n1967 & ~n1968;
  assign \outreg_new<34>  = n1966 | ~n1969;
  assign n1971 = \outreg<38>  & n510;
  assign n1972 = \outreg<30>  & n508;
  assign n1973 = \data<60>  & n504;
  assign n1974 = ~n1972 & ~n1973;
  assign \outreg_new<30>  = n1971 | ~n1974;
  assign n1976 = n1610 & n1699;
  assign n1977 = ~n1607 & n1976;
  assign n1978 = ~n1607 & n1636;
  assign n1979 = n1607 & n1631;
  assign n1980 = ~n1607 & n1648;
  assign n1981 = ~n1607 & n1657;
  assign n1982 = n1607 & n1659;
  assign n1983 = ~n1610 & n1668;
  assign n1984 = n1607 & n1983;
  assign n1985 = n1607 & n1673;
  assign n1986 = ~n1607 & n1681;
  assign n1987 = n1607 & n1679;
  assign n1988 = ~n1607 & n1706;
  assign n1989 = n1607 & n1697;
  assign n1990 = ~n1610 & n1625;
  assign n1991 = n1607 & n1990;
  assign n1992 = n1610 & n1645;
  assign n1993 = ~n1607 & n1992;
  assign n1994 = ~n1607 & n1664;
  assign n1995 = ~n1701 & ~n1989;
  assign n1996 = ~n1698 & n1995;
  assign n1997 = ~n1988 & n1996;
  assign n1998 = ~n1692 & n1997;
  assign n1999 = ~n1689 & n1998;
  assign n2000 = ~n1685 & n1999;
  assign n2001 = ~n1987 & n2000;
  assign n2002 = ~n1986 & n2001;
  assign n2003 = ~n1680 & n2002;
  assign n2004 = ~n1985 & n2003;
  assign n2005 = ~n1678 & n2004;
  assign n2006 = ~n1670 & n2005;
  assign n2007 = ~n1667 & n2006;
  assign n2008 = ~n1984 & n2007;
  assign n2009 = ~n1982 & n2008;
  assign n2010 = ~n1660 & n2009;
  assign n2011 = ~n1658 & n2010;
  assign n2012 = ~n1981 & n2011;
  assign n2013 = ~n1649 & n2012;
  assign n2014 = ~n1980 & n2013;
  assign n2015 = ~n1647 & n2014;
  assign n2016 = ~n1644 & n2015;
  assign n2017 = ~n1641 & n2016;
  assign n2018 = ~n1979 & n2017;
  assign n2019 = ~n1978 & n2018;
  assign n2020 = ~n1627 & n2019;
  assign n2021 = ~n1977 & n2020;
  assign n2022 = ~n1610 & n1686;
  assign n2023 = ~n1607 & n2022;
  assign n2024 = n2021 & ~n2023;
  assign n2025 = ~n1994 & n2024;
  assign n2026 = ~n1993 & n2025;
  assign n2027 = ~n1991 & n2026;
  assign n2028 = \data<27>  & n504;
  assign n2029 = n2027 & n2028;
  assign n2030 = ~\data<27>  & n504;
  assign n2031 = ~n2027 & n2030;
  assign n2032 = \outreg<47>  & n510;
  assign n2033 = \outreg<39>  & n508;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~n2031 & n2034;
  assign \outreg_new<39>  = n2029 | ~n2035;
  assign n2037 = ~n1271 & n1367;
  assign n2038 = ~n1271 & n1315;
  assign n2039 = ~n1271 & n1325;
  assign n2040 = n1271 & n1369;
  assign n2041 = n1274 & n1321;
  assign n2042 = n1271 & n2041;
  assign n2043 = ~n1274 & n1324;
  assign n2044 = n1271 & n2043;
  assign n2045 = ~n1271 & n1356;
  assign n2046 = n1274 & n1355;
  assign n2047 = ~n1271 & n2046;
  assign n2048 = n1274 & n1363;
  assign n2049 = ~n1271 & n2048;
  assign n2050 = n1271 & n1399;
  assign n2051 = n1271 & n1337;
  assign n2052 = n1271 & n1344;
  assign n2053 = n1271 & n2048;
  assign n2054 = n1271 & n1308;
  assign n2055 = ~n1271 & n1360;
  assign n2056 = ~n1361 & ~n1362;
  assign n2057 = ~n2052 & n2056;
  assign n2058 = ~n2051 & n2057;
  assign n2059 = ~n1357 & n2058;
  assign n2060 = ~n2050 & n2059;
  assign n2061 = ~n1353 & n2060;
  assign n2062 = ~n2049 & n2061;
  assign n2063 = ~n1349 & n2062;
  assign n2064 = ~n1340 & n2063;
  assign n2065 = ~n2047 & n2064;
  assign n2066 = ~n2045 & n2065;
  assign n2067 = ~n1334 & n2066;
  assign n2068 = ~n1331 & n2067;
  assign n2069 = ~n2044 & n2068;
  assign n2070 = ~n2042 & n2069;
  assign n2071 = ~n1320 & n2070;
  assign n2072 = ~n1319 & n2071;
  assign n2073 = ~n1316 & n2072;
  assign n2074 = ~n1313 & n2073;
  assign n2075 = ~n2040 & n2074;
  assign n2076 = ~n1311 & n2075;
  assign n2077 = ~n2039 & n2076;
  assign n2078 = ~n1303 & n2077;
  assign n2079 = ~n2038 & n2078;
  assign n2080 = ~n1298 & n2079;
  assign n2081 = ~n1294 & n2080;
  assign n2082 = ~n2037 & n2081;
  assign n2083 = ~n1271 & n1322;
  assign n2084 = n2082 & ~n2083;
  assign n2085 = ~n2055 & n2084;
  assign n2086 = ~n2054 & n2085;
  assign n2087 = ~n2053 & n2086;
  assign n2088 = \data<11>  & n504;
  assign n2089 = n2087 & n2088;
  assign n2090 = ~\data<11>  & n504;
  assign n2091 = ~n2087 & n2090;
  assign n2092 = \outreg<43>  & n510;
  assign n2093 = \outreg<35>  & n508;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = ~n2091 & n2094;
  assign \outreg_new<35>  = n2089 | ~n2095;
  assign n2097 = \outreg<44>  & n510;
  assign n2098 = \outreg<36>  & n508;
  assign n2099 = \data<51>  & n504;
  assign n2100 = ~n2098 & ~n2099;
  assign \outreg_new<36>  = n2097 | ~n2100;
  assign n2102 = ~\data<48>  & \C<1> ;
  assign n2103 = \data<48>  & ~\C<1> ;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = \C<12>  & ~\data<47> ;
  assign n2106 = ~\C<12>  & \data<47> ;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = \C<19>  & ~\data<46> ;
  assign n2109 = ~\C<19>  & \data<46> ;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = \C<26>  & ~\data<45> ;
  assign n2112 = ~\C<26>  & \data<45> ;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~\data<44>  & \C<6> ;
  assign n2115 = \data<44>  & ~\C<6> ;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = \C<15>  & ~\data<43> ;
  assign n2118 = ~\C<15>  & \data<43> ;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~n2116 & ~n2119;
  assign n2121 = ~n2113 & n2120;
  assign n2122 = ~n2110 & n2121;
  assign n2123 = ~n2107 & n2122;
  assign n2124 = ~n2104 & n2123;
  assign n2125 = n2110 & n2121;
  assign n2126 = ~n2107 & n2125;
  assign n2127 = ~n2104 & n2126;
  assign n2128 = n2107 & n2125;
  assign n2129 = ~n2104 & n2128;
  assign n2130 = n2113 & n2120;
  assign n2131 = ~n2110 & n2130;
  assign n2132 = n2107 & n2131;
  assign n2133 = ~n2104 & n2132;
  assign n2134 = n2116 & ~n2119;
  assign n2135 = ~n2113 & n2134;
  assign n2136 = ~n2110 & n2135;
  assign n2137 = n2107 & n2136;
  assign n2138 = ~n2104 & n2137;
  assign n2139 = n2113 & n2134;
  assign n2140 = ~n2110 & n2139;
  assign n2141 = ~n2107 & n2140;
  assign n2142 = ~n2104 & n2141;
  assign n2143 = n2110 & n2139;
  assign n2144 = ~n2107 & n2143;
  assign n2145 = ~n2104 & n2144;
  assign n2146 = n2104 & n2128;
  assign n2147 = ~n2107 & n2131;
  assign n2148 = n2104 & n2147;
  assign n2149 = n2110 & n2130;
  assign n2150 = n2107 & n2149;
  assign n2151 = n2104 & n2150;
  assign n2152 = ~n2107 & n2136;
  assign n2153 = n2104 & n2152;
  assign n2154 = n2104 & n2137;
  assign n2155 = n2110 & n2135;
  assign n2156 = n2107 & n2155;
  assign n2157 = n2104 & n2156;
  assign n2158 = n2104 & n2144;
  assign n2159 = ~n2116 & n2119;
  assign n2160 = ~n2113 & n2159;
  assign n2161 = ~n2110 & n2160;
  assign n2162 = n2107 & n2161;
  assign n2163 = ~n2104 & n2162;
  assign n2164 = n2113 & n2159;
  assign n2165 = ~n2110 & n2164;
  assign n2166 = ~n2107 & n2165;
  assign n2167 = ~n2104 & n2166;
  assign n2168 = n2110 & n2164;
  assign n2169 = ~n2107 & n2168;
  assign n2170 = ~n2104 & n2169;
  assign n2171 = n2116 & n2119;
  assign n2172 = ~n2113 & n2171;
  assign n2173 = n2110 & n2172;
  assign n2174 = ~n2107 & n2173;
  assign n2175 = ~n2104 & n2174;
  assign n2176 = n2107 & n2173;
  assign n2177 = ~n2104 & n2176;
  assign n2178 = n2113 & n2171;
  assign n2179 = ~n2110 & n2178;
  assign n2180 = ~n2107 & n2179;
  assign n2181 = ~n2104 & n2180;
  assign n2182 = n2110 & n2178;
  assign n2183 = n2107 & n2182;
  assign n2184 = ~n2104 & n2183;
  assign n2185 = ~n2107 & n2161;
  assign n2186 = n2104 & n2185;
  assign n2187 = n2110 & n2160;
  assign n2188 = ~n2107 & n2187;
  assign n2189 = n2104 & n2188;
  assign n2190 = n2104 & n2166;
  assign n2191 = n2104 & n2174;
  assign n2192 = n2107 & n2179;
  assign n2193 = n2104 & n2192;
  assign n2194 = ~n2107 & n2182;
  assign n2195 = n2104 & n2194;
  assign n2196 = n2104 & n2183;
  assign n2197 = n2104 & n2162;
  assign n2198 = n2104 & n2123;
  assign n2199 = n2107 & n2168;
  assign n2200 = ~n2104 & n2199;
  assign n2201 = ~n2195 & ~n2196;
  assign n2202 = ~n2193 & n2201;
  assign n2203 = ~n2191 & n2202;
  assign n2204 = ~n2190 & n2203;
  assign n2205 = ~n2189 & n2204;
  assign n2206 = ~n2186 & n2205;
  assign n2207 = ~n2184 & n2206;
  assign n2208 = ~n2181 & n2207;
  assign n2209 = ~n2177 & n2208;
  assign n2210 = ~n2175 & n2209;
  assign n2211 = ~n2170 & n2210;
  assign n2212 = ~n2167 & n2211;
  assign n2213 = ~n2163 & n2212;
  assign n2214 = ~n2158 & n2213;
  assign n2215 = ~n2157 & n2214;
  assign n2216 = ~n2154 & n2215;
  assign n2217 = ~n2153 & n2216;
  assign n2218 = ~n2151 & n2217;
  assign n2219 = ~n2148 & n2218;
  assign n2220 = ~n2146 & n2219;
  assign n2221 = ~n2145 & n2220;
  assign n2222 = ~n2142 & n2221;
  assign n2223 = ~n2138 & n2222;
  assign n2224 = ~n2133 & n2223;
  assign n2225 = ~n2129 & n2224;
  assign n2226 = ~n2127 & n2225;
  assign n2227 = ~n2124 & n2226;
  assign n2228 = ~n2107 & n2149;
  assign n2229 = ~n2104 & n2228;
  assign n2230 = n2227 & ~n2229;
  assign n2231 = ~n2200 & n2230;
  assign n2232 = ~n2198 & n2231;
  assign n2233 = ~n2197 & n2232;
  assign n2234 = \data<19>  & n504;
  assign n2235 = n2233 & n2234;
  assign n2236 = ~\data<19>  & n504;
  assign n2237 = ~n2233 & n2236;
  assign n2238 = \outreg<45>  & n510;
  assign n2239 = \outreg<37>  & n508;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n2237 & n2240;
  assign \outreg_new<37>  = n2235 | ~n2241;
  assign n2243 = \outreg<46>  & n510;
  assign n2244 = \outreg<38>  & n508;
  assign n2245 = \data<59>  & n504;
  assign n2246 = ~n2244 & ~n2245;
  assign \outreg_new<38>  = n2243 | ~n2246;
  assign n2248 = ~n880 & n921;
  assign n2249 = ~n880 & n927;
  assign n2250 = ~n880 & n978;
  assign n2251 = n880 & n983;
  assign n2252 = n880 & n903;
  assign n2253 = n880 & n917;
  assign n2254 = ~n883 & n964;
  assign n2255 = ~n880 & n2254;
  assign n2256 = ~n880 & n965;
  assign n2257 = ~n880 & n975;
  assign n2258 = n880 & n938;
  assign n2259 = n880 & n942;
  assign n2260 = n880 & n950;
  assign n2261 = n880 & n919;
  assign n2262 = n880 & n957;
  assign n2263 = n883 & n912;
  assign n2264 = ~n880 & n2263;
  assign n2265 = ~n880 & n971;
  assign n2266 = ~n974 & ~n2260;
  assign n2267 = ~n970 & n2266;
  assign n2268 = ~n2259 & n2267;
  assign n2269 = ~n968 & n2268;
  assign n2270 = ~n966 & n2269;
  assign n2271 = ~n2258 & n2270;
  assign n2272 = ~n2257 & n2271;
  assign n2273 = ~n954 & n2272;
  assign n2274 = ~n951 & n2273;
  assign n2275 = ~n946 & n2274;
  assign n2276 = ~n943 & n2275;
  assign n2277 = ~n2256 & n2276;
  assign n2278 = ~n2255 & n2277;
  assign n2279 = ~n2253 & n2278;
  assign n2280 = ~n934 & n2279;
  assign n2281 = ~n933 & n2280;
  assign n2282 = ~n931 & n2281;
  assign n2283 = ~n2252 & n2282;
  assign n2284 = ~n928 & n2283;
  assign n2285 = ~n2251 & n2284;
  assign n2286 = ~n2250 & n2285;
  assign n2287 = ~n918 & n2286;
  assign n2288 = ~n911 & n2287;
  assign n2289 = ~n904 & n2288;
  assign n2290 = ~n2249 & n2289;
  assign n2291 = ~n900 & n2290;
  assign n2292 = ~n2248 & n2291;
  assign n2293 = ~n2265 & n2292;
  assign n2294 = ~n2264 & n2293;
  assign n2295 = ~n2262 & n2294;
  assign n2296 = ~n2261 & n2295;
  assign n2297 = \data<2>  & n504;
  assign n2298 = n2296 & n2297;
  assign n2299 = ~\data<2>  & n504;
  assign n2300 = ~n2296 & n2299;
  assign n2301 = \outreg<49>  & n510;
  assign n2302 = \outreg<41>  & n508;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~n2300 & n2303;
  assign \outreg_new<41>  = n2298 | ~n2304;
  assign n2306 = \outreg<50>  & n510;
  assign n2307 = \outreg<42>  & n508;
  assign n2308 = \data<42>  & n504;
  assign n2309 = ~n2307 & ~n2308;
  assign \outreg_new<42>  = n2306 | ~n2309;
  assign n2311 = ~n1757 & n1810;
  assign n2312 = n1757 & n1907;
  assign n2313 = ~n1757 & n1838;
  assign n2314 = n1757 & n1817;
  assign n2315 = n1757 & n1909;
  assign n2316 = n1757 & n1828;
  assign n2317 = ~n1757 & n1807;
  assign n2318 = ~n1757 & n1850;
  assign n2319 = ~n1851 & ~n1921;
  assign n2320 = ~n1848 & n2319;
  assign n2321 = ~n2314 & n2320;
  assign n2322 = ~n1844 & n2321;
  assign n2323 = ~n1842 & n2322;
  assign n2324 = ~n1919 & n2323;
  assign n2325 = ~n1917 & n2324;
  assign n2326 = ~n1835 & n2325;
  assign n2327 = ~n1831 & n2326;
  assign n2328 = ~n1821 & n2327;
  assign n2329 = ~n1816 & n2328;
  assign n2330 = ~n1915 & n2329;
  assign n2331 = ~n2313 & n2330;
  assign n2332 = ~n1811 & n2331;
  assign n2333 = ~n1808 & n2332;
  assign n2334 = ~n2312 & n2333;
  assign n2335 = ~n1804 & n2334;
  assign n2336 = ~n1913 & n2335;
  assign n2337 = ~n1912 & n2336;
  assign n2338 = ~n1800 & n2337;
  assign n2339 = ~n2311 & n2338;
  assign n2340 = ~n1792 & n2339;
  assign n2341 = ~n1908 & n2340;
  assign n2342 = ~n1906 & n2341;
  assign n2343 = ~n1787 & n2342;
  assign n2344 = ~n1784 & n2343;
  assign n2345 = ~n1780 & n2344;
  assign n2346 = ~n2318 & n2345;
  assign n2347 = ~n2317 & n2346;
  assign n2348 = ~n2316 & n2347;
  assign n2349 = ~n2315 & n2348;
  assign n2350 = \data<10>  & n504;
  assign n2351 = n2349 & n2350;
  assign n2352 = ~\data<10>  & n504;
  assign n2353 = ~n2349 & n2352;
  assign n2354 = \outreg<51>  & n510;
  assign n2355 = \outreg<43>  & n508;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = ~n2353 & n2356;
  assign \outreg_new<43>  = n2351 | ~n2357;
  assign n2359 = \outreg<52>  & n510;
  assign n2360 = \outreg<44>  & n508;
  assign n2361 = \data<50>  & n504;
  assign n2362 = ~n2360 & ~n2361;
  assign \outreg_new<44>  = n2359 | ~n2362;
  assign n2364 = \outreg<48>  & n510;
  assign n2365 = \outreg<40>  & n508;
  assign n2366 = \data<34>  & n504;
  assign n2367 = ~n2365 & ~n2366;
  assign \outreg_new<40>  = n2364 | ~n2367;
  assign n2369 = n1607 & n1992;
  assign n2370 = ~n1607 & n1983;
  assign n2371 = n1607 & n2022;
  assign n2372 = n1607 & n1691;
  assign n2373 = n1607 & n1643;
  assign n2374 = ~n1607 & n1661;
  assign n2375 = ~n1607 & n1684;
  assign n2376 = ~n1607 & n1695;
  assign n2377 = n1709 & ~n1988;
  assign n2378 = ~n2372 & n2377;
  assign n2379 = ~n1692 & n2378;
  assign n2380 = ~n1688 & n2379;
  assign n2381 = ~n2371 & n2380;
  assign n2382 = ~n1685 & n2381;
  assign n2383 = ~n1682 & n2382;
  assign n2384 = ~n1987 & n2383;
  assign n2385 = ~n1986 & n2384;
  assign n2386 = ~n1678 & n2385;
  assign n2387 = ~n1670 & n2386;
  assign n2388 = ~n1667 & n2387;
  assign n2389 = ~n1984 & n2388;
  assign n2390 = ~n1665 & n2389;
  assign n2391 = ~n2370 & n2390;
  assign n2392 = ~n1982 & n2391;
  assign n2393 = ~n1653 & n2392;
  assign n2394 = ~n2369 & n2393;
  assign n2395 = ~n1980 & n2394;
  assign n2396 = ~n1647 & n2395;
  assign n2397 = ~n1644 & n2396;
  assign n2398 = ~n1639 & n2397;
  assign n2399 = ~n1979 & n2398;
  assign n2400 = ~n1632 & n2399;
  assign n2401 = ~n1627 & n2400;
  assign n2402 = ~n1977 & n2401;
  assign n2403 = ~n2376 & n2402;
  assign n2404 = ~n2375 & n2403;
  assign n2405 = ~n2374 & n2404;
  assign n2406 = ~n2373 & n2405;
  assign n2407 = \data<1>  & n504;
  assign n2408 = n2406 & n2407;
  assign n2409 = ~\data<1>  & n504;
  assign n2410 = ~n2406 & n2409;
  assign n2411 = \outreg<57>  & n510;
  assign n2412 = \outreg<49>  & n508;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2410 & n2413;
  assign \outreg_new<49>  = n2408 | ~n2414;
  assign n2416 = n1757 & n1779;
  assign n2417 = n1757 & n1834;
  assign n2418 = ~n1851 & ~n1920;
  assign n2419 = ~n1846 & n2418;
  assign n2420 = ~n2314 & n2419;
  assign n2421 = ~n1842 & n2420;
  assign n2422 = ~n1839 & n2421;
  assign n2423 = ~n1919 & n2422;
  assign n2424 = ~n1835 & n2423;
  assign n2425 = ~n1831 & n2424;
  assign n2426 = ~n1916 & n2425;
  assign n2427 = ~n1826 & n2426;
  assign n2428 = ~n1818 & n2427;
  assign n2429 = ~n1915 & n2428;
  assign n2430 = ~n2313 & n2429;
  assign n2431 = ~n1914 & n2430;
  assign n2432 = ~n1808 & n2431;
  assign n2433 = ~n1806 & n2432;
  assign n2434 = ~n2312 & n2433;
  assign n2435 = ~n1804 & n2434;
  assign n2436 = ~n1802 & n2435;
  assign n2437 = ~n1912 & n2436;
  assign n2438 = ~n2311 & n2437;
  assign n2439 = ~n1910 & n2438;
  assign n2440 = ~n1795 & n2439;
  assign n2441 = ~n1792 & n2440;
  assign n2442 = ~n1906 & n2441;
  assign n2443 = ~n1784 & n2442;
  assign n2444 = ~n1777 & n2443;
  assign n2445 = ~n1757 & n1845;
  assign n2446 = n2444 & ~n2445;
  assign n2447 = ~n1757 & n1854;
  assign n2448 = n2446 & ~n2447;
  assign n2449 = ~n2417 & n2448;
  assign n2450 = ~n2416 & n2449;
  assign n2451 = \data<18>  & n504;
  assign n2452 = n2450 & n2451;
  assign n2453 = ~\data<18>  & n504;
  assign n2454 = ~n2450 & n2453;
  assign n2455 = \outreg<53>  & n510;
  assign n2456 = \outreg<45>  & n508;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2454 & n2457;
  assign \outreg_new<45>  = n2452 | ~n2458;
  assign n2460 = \outreg<54>  & n510;
  assign n2461 = \outreg<46>  & n508;
  assign n2462 = \data<58>  & n504;
  assign n2463 = ~n2461 & ~n2462;
  assign \outreg_new<46>  = n2460 | ~n2463;
  assign n2465 = n536 & n575;
  assign n2466 = n536 & n1560;
  assign n2467 = ~n536 & n1494;
  assign n2468 = ~n536 & n1509;
  assign n2469 = ~n628 & ~n1507;
  assign n2470 = ~n627 & n2469;
  assign n2471 = ~n621 & n2470;
  assign n2472 = ~n1504 & n2471;
  assign n2473 = ~n1556 & n2472;
  assign n2474 = ~n620 & n2473;
  assign n2475 = ~n617 & n2474;
  assign n2476 = ~n1502 & n2475;
  assign n2477 = ~n608 & n2476;
  assign n2478 = ~n1555 & n2477;
  assign n2479 = ~n1499 & n2478;
  assign n2480 = ~n603 & n2479;
  assign n2481 = ~n597 & n2480;
  assign n2482 = ~n592 & n2481;
  assign n2483 = ~n1554 & n2482;
  assign n2484 = ~n587 & n2483;
  assign n2485 = ~n584 & n2484;
  assign n2486 = ~n1493 & n2485;
  assign n2487 = ~n579 & n2486;
  assign n2488 = ~n1491 & n2487;
  assign n2489 = ~n576 & n2488;
  assign n2490 = ~n574 & n2489;
  assign n2491 = ~n1490 & n2490;
  assign n2492 = ~n565 & n2491;
  assign n2493 = ~n1553 & n2492;
  assign n2494 = ~n1488 & n2493;
  assign n2495 = ~n558 & n2494;
  assign n2496 = ~n2468 & n2495;
  assign n2497 = ~n2467 & n2496;
  assign n2498 = ~n2466 & n2497;
  assign n2499 = ~n2465 & n2498;
  assign n2500 = \data<26>  & n504;
  assign n2501 = n2499 & n2500;
  assign n2502 = ~\data<26>  & n504;
  assign n2503 = ~n2499 & n2502;
  assign n2504 = \outreg<55>  & n510;
  assign n2505 = \outreg<47>  & n508;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = ~n2503 & n2506;
  assign \outreg_new<47>  = n2501 | ~n2507;
  assign n2509 = \outreg<56>  & n510;
  assign n2510 = \outreg<48>  & n508;
  assign n2511 = \data<33>  & n504;
  assign n2512 = ~n2510 & ~n2511;
  assign \outreg_new<48>  = n2509 | ~n2512;
  assign n2514 = ~\count<0>  & ~\count<1> ;
  assign n2515 = ~\count<2>  & n2514;
  assign n2516 = ~\count<3>  & n2515;
  assign n2517 = ~\count<3>  & n503;
  assign n2518 = ~\count<0>  & \count<1> ;
  assign n2519 = \count<2>  & n2518;
  assign n2520 = \count<3>  & n2519;
  assign n2521 = ~n504 & ~n2520;
  assign n2522 = ~n2517 & n2521;
  assign n2523 = ~n2516 & n2522;
  assign n2524 = \encrypt<0>  & n504;
  assign n2525 = ~\encrypt_mode<0>  & n2524;
  assign n2526 = ~\encrypt<0>  & n504;
  assign n2527 = \encrypt_mode<0>  & n2526;
  assign n2528 = ~n2525 & ~n2527;
  assign n2529 = \C<21>  & ~n674;
  assign n2530 = ~\encrypt_mode<0>  & n2529;
  assign n2531 = n2528 & n2530;
  assign n2532 = n2523 & n2531;
  assign n2533 = ~\reset<0>  & n2532;
  assign n2534 = \C<25>  & ~n674;
  assign n2535 = \encrypt_mode<0>  & n2534;
  assign n2536 = n2528 & n2535;
  assign n2537 = n2523 & n2536;
  assign n2538 = ~\reset<0>  & n2537;
  assign n2539 = \C<22>  & ~n674;
  assign n2540 = ~\encrypt_mode<0>  & n2539;
  assign n2541 = n2528 & n2540;
  assign n2542 = ~n2523 & n2541;
  assign n2543 = ~\reset<0>  & n2542;
  assign n2544 = \C<24>  & ~n674;
  assign n2545 = \encrypt_mode<0>  & n2544;
  assign n2546 = n2528 & n2545;
  assign n2547 = ~n2523 & n2546;
  assign n2548 = ~\reset<0>  & n2547;
  assign n2549 = \encrypt<0>  & n674;
  assign n2550 = \inreg<51>  & n2549;
  assign n2551 = ~\reset<0>  & n2550;
  assign n2552 = \C<23>  & ~n674;
  assign n2553 = ~n2528 & n2552;
  assign n2554 = ~\reset<0>  & n2553;
  assign n2555 = \data_in<2>  & n674;
  assign n2556 = ~\encrypt<0>  & n2555;
  assign n2557 = ~\reset<0>  & n2556;
  assign n2558 = ~n2554 & ~n2557;
  assign n2559 = ~n2551 & n2558;
  assign n2560 = ~n2548 & n2559;
  assign n2561 = ~n2543 & n2560;
  assign n2562 = ~n2538 & n2561;
  assign \C_new<23>  = n2533 | ~n2562;
  assign n2564 = n2523 & n2541;
  assign n2565 = ~\reset<0>  & n2564;
  assign n2566 = \C<26>  & ~n674;
  assign n2567 = \encrypt_mode<0>  & n2566;
  assign n2568 = n2528 & n2567;
  assign n2569 = n2523 & n2568;
  assign n2570 = ~\reset<0>  & n2569;
  assign n2571 = ~\encrypt_mode<0>  & n2552;
  assign n2572 = n2528 & n2571;
  assign n2573 = ~n2523 & n2572;
  assign n2574 = ~\reset<0>  & n2573;
  assign n2575 = ~n2523 & n2536;
  assign n2576 = ~\reset<0>  & n2575;
  assign n2577 = ~\encrypt<0>  & n674;
  assign n2578 = \inreg<51>  & n2577;
  assign n2579 = ~\reset<0>  & n2578;
  assign n2580 = ~n2528 & n2544;
  assign n2581 = ~\reset<0>  & n2580;
  assign n2582 = \inreg<43>  & n2549;
  assign n2583 = ~\reset<0>  & n2582;
  assign n2584 = ~n2581 & ~n2583;
  assign n2585 = ~n2579 & n2584;
  assign n2586 = ~n2576 & n2585;
  assign n2587 = ~n2574 & n2586;
  assign n2588 = ~n2570 & n2587;
  assign \C_new<24>  = n2565 | ~n2588;
  assign n2590 = \C<19>  & ~n674;
  assign n2591 = ~\encrypt_mode<0>  & n2590;
  assign n2592 = n2528 & n2591;
  assign n2593 = n2523 & n2592;
  assign n2594 = ~\reset<0>  & n2593;
  assign n2595 = \encrypt_mode<0>  & n2552;
  assign n2596 = n2528 & n2595;
  assign n2597 = n2523 & n2596;
  assign n2598 = ~\reset<0>  & n2597;
  assign n2599 = \C<20>  & ~n674;
  assign n2600 = ~\encrypt_mode<0>  & n2599;
  assign n2601 = n2528 & n2600;
  assign n2602 = ~n2523 & n2601;
  assign n2603 = ~\reset<0>  & n2602;
  assign n2604 = \encrypt_mode<0>  & n2539;
  assign n2605 = n2528 & n2604;
  assign n2606 = ~n2523 & n2605;
  assign n2607 = ~\reset<0>  & n2606;
  assign n2608 = \inreg<2>  & n2549;
  assign n2609 = ~\reset<0>  & n2608;
  assign n2610 = \inreg<10>  & n2577;
  assign n2611 = ~\reset<0>  & n2610;
  assign n2612 = ~n2528 & n2529;
  assign n2613 = ~\reset<0>  & n2612;
  assign n2614 = ~n2611 & ~n2613;
  assign n2615 = ~n2609 & n2614;
  assign n2616 = ~n2607 & n2615;
  assign n2617 = ~n2603 & n2616;
  assign n2618 = ~n2598 & n2617;
  assign \C_new<21>  = n2594 | ~n2618;
  assign n2620 = n2523 & n2601;
  assign n2621 = ~\reset<0>  & n2620;
  assign n2622 = n2523 & n2546;
  assign n2623 = ~\reset<0>  & n2622;
  assign n2624 = ~n2523 & n2531;
  assign n2625 = ~\reset<0>  & n2624;
  assign n2626 = ~n2523 & n2596;
  assign n2627 = ~\reset<0>  & n2626;
  assign n2628 = \inreg<2>  & n2577;
  assign n2629 = ~\reset<0>  & n2628;
  assign n2630 = ~n2528 & n2539;
  assign n2631 = ~\reset<0>  & n2630;
  assign n2632 = \encrypt<0>  & n2555;
  assign n2633 = ~\reset<0>  & n2632;
  assign n2634 = ~n2631 & ~n2633;
  assign n2635 = ~n2629 & n2634;
  assign n2636 = ~n2627 & n2635;
  assign n2637 = ~n2625 & n2636;
  assign n2638 = ~n2623 & n2637;
  assign \C_new<22>  = n2621 | ~n2638;
  assign n2640 = \C<18>  & ~n674;
  assign n2641 = ~\encrypt_mode<0>  & n2640;
  assign n2642 = n2528 & n2641;
  assign n2643 = n2523 & n2642;
  assign n2644 = ~\reset<0>  & n2643;
  assign n2645 = n2523 & n2605;
  assign n2646 = ~\reset<0>  & n2645;
  assign n2647 = ~n2523 & n2592;
  assign n2648 = ~\reset<0>  & n2647;
  assign n2649 = \encrypt_mode<0>  & n2529;
  assign n2650 = n2528 & n2649;
  assign n2651 = ~n2523 & n2650;
  assign n2652 = ~\reset<0>  & n2651;
  assign n2653 = \inreg<18>  & n2577;
  assign n2654 = ~\reset<0>  & n2653;
  assign n2655 = ~n2528 & n2599;
  assign n2656 = ~\reset<0>  & n2655;
  assign n2657 = \inreg<10>  & n2549;
  assign n2658 = ~\reset<0>  & n2657;
  assign n2659 = ~n2656 & ~n2658;
  assign n2660 = ~n2654 & n2659;
  assign n2661 = ~n2652 & n2660;
  assign n2662 = ~n2648 & n2661;
  assign n2663 = ~n2646 & n2662;
  assign \C_new<20>  = n2644 | ~n2663;
  assign n2665 = \data<36>  & ~n504;
  assign n2666 = \inreg<17>  & n504;
  assign \data_new<4>  = n2665 | n2666;
  assign n2668 = \data<35>  & ~n504;
  assign n2669 = \inreg<25>  & n504;
  assign \data_new<3>  = n2668 | n2669;
  assign n2671 = ~\encrypt_mode<0>  & n2534;
  assign n2672 = n2528 & n2671;
  assign n2673 = n2523 & n2672;
  assign n2674 = ~\reset<0>  & n2673;
  assign n2675 = \C<1>  & ~n674;
  assign n2676 = \encrypt_mode<0>  & n2675;
  assign n2677 = n2528 & n2676;
  assign n2678 = n2523 & n2677;
  assign n2679 = ~\reset<0>  & n2678;
  assign n2680 = ~\encrypt_mode<0>  & n2566;
  assign n2681 = n2528 & n2680;
  assign n2682 = ~n2523 & n2681;
  assign n2683 = ~\reset<0>  & n2682;
  assign n2684 = \C<0>  & ~n674;
  assign n2685 = \encrypt_mode<0>  & n2684;
  assign n2686 = n2528 & n2685;
  assign n2687 = ~n2523 & n2686;
  assign n2688 = ~\reset<0>  & n2687;
  assign n2689 = \inreg<48>  & n2549;
  assign n2690 = ~\reset<0>  & n2689;
  assign n2691 = \inreg<27>  & n2577;
  assign n2692 = ~\reset<0>  & n2691;
  assign n2693 = \C<27>  & ~n674;
  assign n2694 = ~n2528 & n2693;
  assign n2695 = ~\reset<0>  & n2694;
  assign n2696 = ~n2692 & ~n2695;
  assign n2697 = ~n2690 & n2696;
  assign n2698 = ~n2688 & n2697;
  assign n2699 = ~n2683 & n2698;
  assign n2700 = ~n2679 & n2699;
  assign \C_new<27>  = n2674 | ~n2700;
  assign n2702 = \data<34>  & ~n504;
  assign n2703 = \inreg<33>  & n504;
  assign \data_new<2>  = n2702 | n2703;
  assign n2705 = \data<33>  & ~n504;
  assign n2706 = \inreg<41>  & n504;
  assign \data_new<1>  = n2705 | n2706;
  assign n2708 = n2523 & n2572;
  assign n2709 = ~\reset<0>  & n2708;
  assign n2710 = \encrypt_mode<0>  & n2693;
  assign n2711 = n2528 & n2710;
  assign n2712 = n2523 & n2711;
  assign n2713 = ~\reset<0>  & n2712;
  assign n2714 = ~\encrypt_mode<0>  & n2544;
  assign n2715 = n2528 & n2714;
  assign n2716 = ~n2523 & n2715;
  assign n2717 = ~\reset<0>  & n2716;
  assign n2718 = ~n2523 & n2568;
  assign n2719 = ~\reset<0>  & n2718;
  assign n2720 = \inreg<43>  & n2577;
  assign n2721 = ~\reset<0>  & n2720;
  assign n2722 = ~n2528 & n2534;
  assign n2723 = ~\reset<0>  & n2722;
  assign n2724 = \inreg<35>  & n2549;
  assign n2725 = ~\reset<0>  & n2724;
  assign n2726 = ~n2723 & ~n2725;
  assign n2727 = ~n2721 & n2726;
  assign n2728 = ~n2719 & n2727;
  assign n2729 = ~n2717 & n2728;
  assign n2730 = ~n2713 & n2729;
  assign \C_new<25>  = n2709 | ~n2730;
  assign n2732 = \data<32>  & ~n504;
  assign n2733 = \inreg<49>  & n504;
  assign \data_new<0>  = n2732 | n2733;
  assign n2735 = n2523 & n2715;
  assign n2736 = ~\reset<0>  & n2735;
  assign n2737 = n2523 & n2686;
  assign n2738 = ~\reset<0>  & n2737;
  assign n2739 = ~n2523 & n2672;
  assign n2740 = ~\reset<0>  & n2739;
  assign n2741 = ~n2523 & n2711;
  assign n2742 = ~\reset<0>  & n2741;
  assign n2743 = \inreg<35>  & n2577;
  assign n2744 = ~\reset<0>  & n2743;
  assign n2745 = ~n2528 & n2566;
  assign n2746 = ~\reset<0>  & n2745;
  assign n2747 = \inreg<27>  & n2549;
  assign n2748 = ~\reset<0>  & n2747;
  assign n2749 = ~n2746 & ~n2748;
  assign n2750 = ~n2744 & n2749;
  assign n2751 = ~n2742 & n2750;
  assign n2752 = ~n2740 & n2751;
  assign n2753 = ~n2738 & n2752;
  assign \C_new<26>  = n2736 | ~n2753;
  assign n2755 = \C<11>  & ~n674;
  assign n2756 = ~\encrypt_mode<0>  & n2755;
  assign n2757 = n2528 & n2756;
  assign n2758 = n2523 & n2757;
  assign n2759 = ~\reset<0>  & n2758;
  assign n2760 = \C<15>  & ~n674;
  assign n2761 = \encrypt_mode<0>  & n2760;
  assign n2762 = n2528 & n2761;
  assign n2763 = n2523 & n2762;
  assign n2764 = ~\reset<0>  & n2763;
  assign n2765 = \C<12>  & ~n674;
  assign n2766 = ~\encrypt_mode<0>  & n2765;
  assign n2767 = n2528 & n2766;
  assign n2768 = ~n2523 & n2767;
  assign n2769 = ~\reset<0>  & n2768;
  assign n2770 = \C<14>  & ~n674;
  assign n2771 = \encrypt_mode<0>  & n2770;
  assign n2772 = n2528 & n2771;
  assign n2773 = ~n2523 & n2772;
  assign n2774 = ~\reset<0>  & n2773;
  assign n2775 = \inreg<9>  & n2577;
  assign n2776 = ~\reset<0>  & n2775;
  assign n2777 = \C<13>  & ~n674;
  assign n2778 = ~n2528 & n2777;
  assign n2779 = ~\reset<0>  & n2778;
  assign n2780 = \inreg<1>  & n2549;
  assign n2781 = ~\reset<0>  & n2780;
  assign n2782 = ~n2779 & ~n2781;
  assign n2783 = ~n2776 & n2782;
  assign n2784 = ~n2774 & n2783;
  assign n2785 = ~n2769 & n2784;
  assign n2786 = ~n2764 & n2785;
  assign \C_new<13>  = n2759 | ~n2786;
  assign n2788 = n2523 & n2767;
  assign n2789 = ~\reset<0>  & n2788;
  assign n2790 = \C<16>  & ~n674;
  assign n2791 = \encrypt_mode<0>  & n2790;
  assign n2792 = n2528 & n2791;
  assign n2793 = n2523 & n2792;
  assign n2794 = ~\reset<0>  & n2793;
  assign n2795 = ~\encrypt_mode<0>  & n2777;
  assign n2796 = n2528 & n2795;
  assign n2797 = ~n2523 & n2796;
  assign n2798 = ~\reset<0>  & n2797;
  assign n2799 = ~n2523 & n2762;
  assign n2800 = ~\reset<0>  & n2799;
  assign n2801 = \inreg<1>  & n2577;
  assign n2802 = ~\reset<0>  & n2801;
  assign n2803 = ~n2528 & n2770;
  assign n2804 = ~\reset<0>  & n2803;
  assign n2805 = \data_in<1>  & n674;
  assign n2806 = \encrypt<0>  & n2805;
  assign n2807 = ~\reset<0>  & n2806;
  assign n2808 = ~n2804 & ~n2807;
  assign n2809 = ~n2802 & n2808;
  assign n2810 = ~n2800 & n2809;
  assign n2811 = ~n2798 & n2810;
  assign n2812 = ~n2794 & n2811;
  assign \C_new<14>  = n2789 | ~n2812;
  assign n2814 = \C<9>  & ~n674;
  assign n2815 = ~\encrypt_mode<0>  & n2814;
  assign n2816 = n2528 & n2815;
  assign n2817 = n2523 & n2816;
  assign n2818 = ~\reset<0>  & n2817;
  assign n2819 = \encrypt_mode<0>  & n2777;
  assign n2820 = n2528 & n2819;
  assign n2821 = n2523 & n2820;
  assign n2822 = ~\reset<0>  & n2821;
  assign n2823 = \C<10>  & ~n674;
  assign n2824 = ~\encrypt_mode<0>  & n2823;
  assign n2825 = n2528 & n2824;
  assign n2826 = ~n2523 & n2825;
  assign n2827 = ~\reset<0>  & n2826;
  assign n2828 = \encrypt_mode<0>  & n2765;
  assign n2829 = n2528 & n2828;
  assign n2830 = ~n2523 & n2829;
  assign n2831 = ~\reset<0>  & n2830;
  assign n2832 = \inreg<25>  & n2577;
  assign n2833 = ~\reset<0>  & n2832;
  assign n2834 = ~n2528 & n2755;
  assign n2835 = ~\reset<0>  & n2834;
  assign n2836 = \inreg<17>  & n2549;
  assign n2837 = ~\reset<0>  & n2836;
  assign n2838 = ~n2835 & ~n2837;
  assign n2839 = ~n2833 & n2838;
  assign n2840 = ~n2831 & n2839;
  assign n2841 = ~n2827 & n2840;
  assign n2842 = ~n2822 & n2841;
  assign \C_new<11>  = n2818 | ~n2842;
  assign n2844 = n2523 & n2825;
  assign n2845 = ~\reset<0>  & n2844;
  assign n2846 = n2523 & n2772;
  assign n2847 = ~\reset<0>  & n2846;
  assign n2848 = ~n2523 & n2757;
  assign n2849 = ~\reset<0>  & n2848;
  assign n2850 = ~n2523 & n2820;
  assign n2851 = ~\reset<0>  & n2850;
  assign n2852 = \inreg<9>  & n2549;
  assign n2853 = ~\reset<0>  & n2852;
  assign n2854 = \inreg<17>  & n2577;
  assign n2855 = ~\reset<0>  & n2854;
  assign n2856 = ~n2528 & n2765;
  assign n2857 = ~\reset<0>  & n2856;
  assign n2858 = ~n2855 & ~n2857;
  assign n2859 = ~n2853 & n2858;
  assign n2860 = ~n2851 & n2859;
  assign n2861 = ~n2849 & n2860;
  assign n2862 = ~n2847 & n2861;
  assign \C_new<12>  = n2845 | ~n2862;
  assign n2864 = \C<8>  & ~n674;
  assign n2865 = ~\encrypt_mode<0>  & n2864;
  assign n2866 = n2528 & n2865;
  assign n2867 = n2523 & n2866;
  assign n2868 = ~\reset<0>  & n2867;
  assign n2869 = n2523 & n2829;
  assign n2870 = ~\reset<0>  & n2869;
  assign n2871 = ~n2523 & n2816;
  assign n2872 = ~\reset<0>  & n2871;
  assign n2873 = \encrypt_mode<0>  & n2755;
  assign n2874 = n2528 & n2873;
  assign n2875 = ~n2523 & n2874;
  assign n2876 = ~\reset<0>  & n2875;
  assign n2877 = \inreg<33>  & n2577;
  assign n2878 = ~\reset<0>  & n2877;
  assign n2879 = ~n2528 & n2823;
  assign n2880 = ~\reset<0>  & n2879;
  assign n2881 = \inreg<25>  & n2549;
  assign n2882 = ~\reset<0>  & n2881;
  assign n2883 = ~n2880 & ~n2882;
  assign n2884 = ~n2878 & n2883;
  assign n2885 = ~n2876 & n2884;
  assign n2886 = ~n2872 & n2885;
  assign n2887 = ~n2870 & n2886;
  assign \C_new<10>  = n2868 | ~n2887;
  assign n2889 = \data<41>  & ~n504;
  assign n2890 = \inreg<43>  & n504;
  assign \data_new<9>  = n2889 | n2890;
  assign n2892 = \data<40>  & ~n504;
  assign n2893 = \inreg<51>  & n504;
  assign \data_new<8>  = n2892 | n2893;
  assign n2895 = \data<39>  & ~n504;
  assign n2896 = \data_in<1>  & n504;
  assign \data_new<7>  = n2895 | n2896;
  assign n2898 = \data<38>  & ~n504;
  assign n2899 = \inreg<1>  & n504;
  assign \data_new<6>  = n2898 | n2899;
  assign n2901 = \data<37>  & ~n504;
  assign n2902 = \inreg<9>  & n504;
  assign \data_new<5>  = n2901 | n2902;
  assign n2904 = \C<17>  & ~n674;
  assign n2905 = ~\encrypt_mode<0>  & n2904;
  assign n2906 = n2528 & n2905;
  assign n2907 = n2523 & n2906;
  assign n2908 = ~\reset<0>  & n2907;
  assign n2909 = n2523 & n2650;
  assign n2910 = ~\reset<0>  & n2909;
  assign n2911 = ~n2523 & n2642;
  assign n2912 = ~\reset<0>  & n2911;
  assign n2913 = \encrypt_mode<0>  & n2599;
  assign n2914 = n2528 & n2913;
  assign n2915 = ~n2523 & n2914;
  assign n2916 = ~\reset<0>  & n2915;
  assign n2917 = \inreg<26>  & n2577;
  assign n2918 = ~\reset<0>  & n2917;
  assign n2919 = ~n2528 & n2590;
  assign n2920 = ~\reset<0>  & n2919;
  assign n2921 = \inreg<18>  & n2549;
  assign n2922 = ~\reset<0>  & n2921;
  assign n2923 = ~n2920 & ~n2922;
  assign n2924 = ~n2918 & n2923;
  assign n2925 = ~n2916 & n2924;
  assign n2926 = ~n2912 & n2925;
  assign n2927 = ~n2910 & n2926;
  assign \C_new<19>  = n2908 | ~n2927;
  assign n2929 = ~\encrypt_mode<0>  & n2760;
  assign n2930 = n2528 & n2929;
  assign n2931 = n2523 & n2930;
  assign n2932 = ~\reset<0>  & n2931;
  assign n2933 = \encrypt_mode<0>  & n2590;
  assign n2934 = n2528 & n2933;
  assign n2935 = n2523 & n2934;
  assign n2936 = ~\reset<0>  & n2935;
  assign n2937 = ~\encrypt_mode<0>  & n2790;
  assign n2938 = n2528 & n2937;
  assign n2939 = ~n2523 & n2938;
  assign n2940 = ~\reset<0>  & n2939;
  assign n2941 = \encrypt_mode<0>  & n2640;
  assign n2942 = n2528 & n2941;
  assign n2943 = ~n2523 & n2942;
  assign n2944 = ~\reset<0>  & n2943;
  assign n2945 = \inreg<42>  & n2577;
  assign n2946 = ~\reset<0>  & n2945;
  assign n2947 = ~n2528 & n2904;
  assign n2948 = ~\reset<0>  & n2947;
  assign n2949 = \inreg<34>  & n2549;
  assign n2950 = ~\reset<0>  & n2949;
  assign n2951 = ~n2948 & ~n2950;
  assign n2952 = ~n2946 & n2951;
  assign n2953 = ~n2944 & n2952;
  assign n2954 = ~n2940 & n2953;
  assign n2955 = ~n2936 & n2954;
  assign \C_new<17>  = n2932 | ~n2955;
  assign n2957 = n2523 & n2938;
  assign n2958 = ~\reset<0>  & n2957;
  assign n2959 = n2523 & n2914;
  assign n2960 = ~\reset<0>  & n2959;
  assign n2961 = ~n2523 & n2906;
  assign n2962 = ~\reset<0>  & n2961;
  assign n2963 = ~n2523 & n2934;
  assign n2964 = ~\reset<0>  & n2963;
  assign n2965 = \inreg<34>  & n2577;
  assign n2966 = ~\reset<0>  & n2965;
  assign n2967 = ~n2528 & n2640;
  assign n2968 = ~\reset<0>  & n2967;
  assign n2969 = \inreg<26>  & n2549;
  assign n2970 = ~\reset<0>  & n2969;
  assign n2971 = ~n2968 & ~n2970;
  assign n2972 = ~n2966 & n2971;
  assign n2973 = ~n2964 & n2972;
  assign n2974 = ~n2962 & n2973;
  assign n2975 = ~n2960 & n2974;
  assign \C_new<18>  = n2958 | ~n2975;
  assign n2977 = n2523 & n2796;
  assign n2978 = ~\reset<0>  & n2977;
  assign n2979 = \encrypt_mode<0>  & n2904;
  assign n2980 = n2528 & n2979;
  assign n2981 = n2523 & n2980;
  assign n2982 = ~\reset<0>  & n2981;
  assign n2983 = ~\encrypt_mode<0>  & n2770;
  assign n2984 = n2528 & n2983;
  assign n2985 = ~n2523 & n2984;
  assign n2986 = ~\reset<0>  & n2985;
  assign n2987 = ~n2523 & n2792;
  assign n2988 = ~\reset<0>  & n2987;
  assign n2989 = \inreg<50>  & n2549;
  assign n2990 = ~\reset<0>  & n2989;
  assign n2991 = ~n2528 & n2760;
  assign n2992 = ~\reset<0>  & n2991;
  assign n2993 = ~\encrypt<0>  & n2805;
  assign n2994 = ~\reset<0>  & n2993;
  assign n2995 = ~n2992 & ~n2994;
  assign n2996 = ~n2990 & n2995;
  assign n2997 = ~n2988 & n2996;
  assign n2998 = ~n2986 & n2997;
  assign n2999 = ~n2982 & n2998;
  assign \C_new<15>  = n2978 | ~n2999;
  assign n3001 = n2523 & n2984;
  assign n3002 = ~\reset<0>  & n3001;
  assign n3003 = n2523 & n2942;
  assign n3004 = ~\reset<0>  & n3003;
  assign n3005 = ~n2523 & n2930;
  assign n3006 = ~\reset<0>  & n3005;
  assign n3007 = ~n2523 & n2980;
  assign n3008 = ~\reset<0>  & n3007;
  assign n3009 = \inreg<50>  & n2577;
  assign n3010 = ~\reset<0>  & n3009;
  assign n3011 = ~n2528 & n2790;
  assign n3012 = ~\reset<0>  & n3011;
  assign n3013 = \inreg<42>  & n2549;
  assign n3014 = ~\reset<0>  & n3013;
  assign n3015 = ~n3012 & ~n3014;
  assign n3016 = ~n3010 & n3015;
  assign n3017 = ~n3008 & n3016;
  assign n3018 = ~n3006 & n3017;
  assign n3019 = ~n3004 & n3018;
  assign \C_new<16>  = n3002 | ~n3019;
  assign n3021 = \D<11>  & ~n674;
  assign n3022 = ~\encrypt_mode<0>  & n3021;
  assign n3023 = n2528 & n3022;
  assign n3024 = n2523 & n3023;
  assign n3025 = ~\reset<0>  & n3024;
  assign n3026 = \D<15>  & ~n674;
  assign n3027 = \encrypt_mode<0>  & n3026;
  assign n3028 = n2528 & n3027;
  assign n3029 = n2523 & n3028;
  assign n3030 = ~\reset<0>  & n3029;
  assign n3031 = \D<12>  & ~n674;
  assign n3032 = ~\encrypt_mode<0>  & n3031;
  assign n3033 = n2528 & n3032;
  assign n3034 = ~n2523 & n3033;
  assign n3035 = ~\reset<0>  & n3034;
  assign n3036 = \D<14>  & ~n674;
  assign n3037 = \encrypt_mode<0>  & n3036;
  assign n3038 = n2528 & n3037;
  assign n3039 = ~n2523 & n3038;
  assign n3040 = ~\reset<0>  & n3039;
  assign n3041 = \inreg<5>  & n2549;
  assign n3042 = ~\reset<0>  & n3041;
  assign n3043 = \inreg<13>  & n2577;
  assign n3044 = ~\reset<0>  & n3043;
  assign n3045 = \D<13>  & ~n674;
  assign n3046 = ~n2528 & n3045;
  assign n3047 = ~\reset<0>  & n3046;
  assign n3048 = ~n3044 & ~n3047;
  assign n3049 = ~n3042 & n3048;
  assign n3050 = ~n3040 & n3049;
  assign n3051 = ~n3035 & n3050;
  assign n3052 = ~n3030 & n3051;
  assign \D_new<13>  = n3025 | ~n3052;
  assign n3054 = n2523 & n3033;
  assign n3055 = ~\reset<0>  & n3054;
  assign n3056 = \D<16>  & ~n674;
  assign n3057 = \encrypt_mode<0>  & n3056;
  assign n3058 = n2528 & n3057;
  assign n3059 = n2523 & n3058;
  assign n3060 = ~\reset<0>  & n3059;
  assign n3061 = ~\encrypt_mode<0>  & n3045;
  assign n3062 = n2528 & n3061;
  assign n3063 = ~n2523 & n3062;
  assign n3064 = ~\reset<0>  & n3063;
  assign n3065 = ~n2523 & n3028;
  assign n3066 = ~\reset<0>  & n3065;
  assign n3067 = \inreg<5>  & n2577;
  assign n3068 = ~\reset<0>  & n3067;
  assign n3069 = ~n2528 & n3036;
  assign n3070 = ~\reset<0>  & n3069;
  assign n3071 = \data_in<5>  & n674;
  assign n3072 = \encrypt<0>  & n3071;
  assign n3073 = ~\reset<0>  & n3072;
  assign n3074 = ~n3070 & ~n3073;
  assign n3075 = ~n3068 & n3074;
  assign n3076 = ~n3066 & n3075;
  assign n3077 = ~n3064 & n3076;
  assign n3078 = ~n3060 & n3077;
  assign \D_new<14>  = n3055 | ~n3078;
  assign n3080 = \D<9>  & ~n674;
  assign n3081 = ~\encrypt_mode<0>  & n3080;
  assign n3082 = n2528 & n3081;
  assign n3083 = n2523 & n3082;
  assign n3084 = ~\reset<0>  & n3083;
  assign n3085 = \encrypt_mode<0>  & n3045;
  assign n3086 = n2528 & n3085;
  assign n3087 = n2523 & n3086;
  assign n3088 = ~\reset<0>  & n3087;
  assign n3089 = \D<10>  & ~n674;
  assign n3090 = ~\encrypt_mode<0>  & n3089;
  assign n3091 = n2528 & n3090;
  assign n3092 = ~n2523 & n3091;
  assign n3093 = ~\reset<0>  & n3092;
  assign n3094 = \encrypt_mode<0>  & n3031;
  assign n3095 = n2528 & n3094;
  assign n3096 = ~n2523 & n3095;
  assign n3097 = ~\reset<0>  & n3096;
  assign n3098 = \inreg<29>  & n2577;
  assign n3099 = ~\reset<0>  & n3098;
  assign n3100 = ~n2528 & n3021;
  assign n3101 = ~\reset<0>  & n3100;
  assign n3102 = \inreg<21>  & n2549;
  assign n3103 = ~\reset<0>  & n3102;
  assign n3104 = ~n3101 & ~n3103;
  assign n3105 = ~n3099 & n3104;
  assign n3106 = ~n3097 & n3105;
  assign n3107 = ~n3093 & n3106;
  assign n3108 = ~n3088 & n3107;
  assign \D_new<11>  = n3084 | ~n3108;
  assign n3110 = n2523 & n3091;
  assign n3111 = ~\reset<0>  & n3110;
  assign n3112 = n2523 & n3038;
  assign n3113 = ~\reset<0>  & n3112;
  assign n3114 = ~n2523 & n3023;
  assign n3115 = ~\reset<0>  & n3114;
  assign n3116 = ~n2523 & n3086;
  assign n3117 = ~\reset<0>  & n3116;
  assign n3118 = \inreg<21>  & n2577;
  assign n3119 = ~\reset<0>  & n3118;
  assign n3120 = ~n2528 & n3031;
  assign n3121 = ~\reset<0>  & n3120;
  assign n3122 = \inreg<13>  & n2549;
  assign n3123 = ~\reset<0>  & n3122;
  assign n3124 = ~n3121 & ~n3123;
  assign n3125 = ~n3119 & n3124;
  assign n3126 = ~n3117 & n3125;
  assign n3127 = ~n3115 & n3126;
  assign n3128 = ~n3113 & n3127;
  assign \D_new<12>  = n3111 | ~n3128;
  assign n3130 = \D<8>  & ~n674;
  assign n3131 = ~\encrypt_mode<0>  & n3130;
  assign n3132 = n2528 & n3131;
  assign n3133 = n2523 & n3132;
  assign n3134 = ~\reset<0>  & n3133;
  assign n3135 = n2523 & n3095;
  assign n3136 = ~\reset<0>  & n3135;
  assign n3137 = ~n2523 & n3082;
  assign n3138 = ~\reset<0>  & n3137;
  assign n3139 = \encrypt_mode<0>  & n3021;
  assign n3140 = n2528 & n3139;
  assign n3141 = ~n2523 & n3140;
  assign n3142 = ~\reset<0>  & n3141;
  assign n3143 = \inreg<37>  & n2577;
  assign n3144 = ~\reset<0>  & n3143;
  assign n3145 = ~n2528 & n3089;
  assign n3146 = ~\reset<0>  & n3145;
  assign n3147 = \inreg<29>  & n2549;
  assign n3148 = ~\reset<0>  & n3147;
  assign n3149 = ~n3146 & ~n3148;
  assign n3150 = ~n3144 & n3149;
  assign n3151 = ~n3142 & n3150;
  assign n3152 = ~n3138 & n3151;
  assign n3153 = ~n3136 & n3152;
  assign \D_new<10>  = n3134 | ~n3153;
  assign n3155 = ~n1271 & n1317;
  assign n3156 = n1271 & n1290;
  assign n3157 = ~n1274 & n1359;
  assign n3158 = ~n1271 & n3157;
  assign n3159 = n1271 & n2046;
  assign n3160 = n1274 & n1343;
  assign n3161 = n1271 & n3160;
  assign n3162 = n1271 & n1297;
  assign n3163 = ~n1271 & n1352;
  assign n3164 = n1372 & ~n2052;
  assign n3165 = ~n2051 & n3164;
  assign n3166 = ~n3159 & n3165;
  assign n3167 = ~n1354 & n3166;
  assign n3168 = ~n2049 & n3167;
  assign n3169 = ~n1351 & n3168;
  assign n3170 = ~n3158 & n3169;
  assign n3171 = ~n1345 & n3170;
  assign n3172 = ~n1340 & n3171;
  assign n3173 = ~n2045 & n3172;
  assign n3174 = ~n1334 & n3173;
  assign n3175 = ~n1326 & n3174;
  assign n3176 = ~n2044 & n3175;
  assign n3177 = ~n2042 & n3176;
  assign n3178 = ~n1319 & n3177;
  assign n3179 = ~n1318 & n3178;
  assign n3180 = ~n1316 & n3179;
  assign n3181 = ~n3156 & n3180;
  assign n3182 = ~n1309 & n3181;
  assign n3183 = ~n2039 & n3182;
  assign n3184 = ~n1305 & n3183;
  assign n3185 = ~n3155 & n3184;
  assign n3186 = ~n1298 & n3185;
  assign n3187 = ~n1294 & n3186;
  assign n3188 = ~n2037 & n3187;
  assign n3189 = ~n1271 & n2043;
  assign n3190 = n3188 & ~n3189;
  assign n3191 = ~n3163 & n3190;
  assign n3192 = ~n3162 & n3191;
  assign n3193 = ~n3161 & n3192;
  assign n3194 = \data<31>  & ~n504;
  assign n3195 = n3193 & n3194;
  assign n3196 = ~\data<31>  & ~n504;
  assign n3197 = ~n3193 & n3196;
  assign n3198 = \data_in<6>  & n504;
  assign n3199 = ~n3197 & ~n3198;
  assign \data_new<63>  = n3195 | ~n3199;
  assign n3201 = \data<29>  & ~n504;
  assign n3202 = n1468 & n3201;
  assign n3203 = ~\data<29>  & ~n504;
  assign n3204 = ~n1468 & n3203;
  assign n3205 = \inreg<14>  & n504;
  assign n3206 = ~n3204 & ~n3205;
  assign \data_new<61>  = n3202 | ~n3206;
  assign n3208 = \data<30>  & ~n504;
  assign n3209 = n1100 & n3208;
  assign n3210 = ~\data<30>  & ~n504;
  assign n3211 = ~n1100 & n3210;
  assign n3212 = \inreg<6>  & n504;
  assign n3213 = ~n3211 & ~n3212;
  assign \data_new<62>  = n3209 | ~n3213;
  assign n3215 = \D<17>  & ~n674;
  assign n3216 = ~\encrypt_mode<0>  & n3215;
  assign n3217 = n2528 & n3216;
  assign n3218 = n2523 & n3217;
  assign n3219 = ~\reset<0>  & n3218;
  assign n3220 = \D<21>  & ~n674;
  assign n3221 = \encrypt_mode<0>  & n3220;
  assign n3222 = n2528 & n3221;
  assign n3223 = n2523 & n3222;
  assign n3224 = ~\reset<0>  & n3223;
  assign n3225 = \D<18>  & ~n674;
  assign n3226 = ~\encrypt_mode<0>  & n3225;
  assign n3227 = n2528 & n3226;
  assign n3228 = ~n2523 & n3227;
  assign n3229 = ~\reset<0>  & n3228;
  assign n3230 = \D<20>  & ~n674;
  assign n3231 = \encrypt_mode<0>  & n3230;
  assign n3232 = n2528 & n3231;
  assign n3233 = ~n2523 & n3232;
  assign n3234 = ~\reset<0>  & n3233;
  assign n3235 = \inreg<28>  & n2577;
  assign n3236 = ~\reset<0>  & n3235;
  assign n3237 = \D<19>  & ~n674;
  assign n3238 = ~n2528 & n3237;
  assign n3239 = ~\reset<0>  & n3238;
  assign n3240 = \inreg<20>  & n2549;
  assign n3241 = ~\reset<0>  & n3240;
  assign n3242 = ~n3239 & ~n3241;
  assign n3243 = ~n3236 & n3242;
  assign n3244 = ~n3234 & n3243;
  assign n3245 = ~n3229 & n3244;
  assign n3246 = ~n3224 & n3245;
  assign \D_new<19>  = n3219 | ~n3246;
  assign n3248 = \data<28>  & ~n504;
  assign n3249 = n1891 & n3248;
  assign n3250 = ~\data<28>  & ~n504;
  assign n3251 = ~n1891 & n3250;
  assign n3252 = \inreg<22>  & n504;
  assign n3253 = ~n3251 & ~n3252;
  assign \data_new<60>  = n3249 | ~n3253;
  assign n3255 = ~\encrypt_mode<0>  & n3026;
  assign n3256 = n2528 & n3255;
  assign n3257 = n2523 & n3256;
  assign n3258 = ~\reset<0>  & n3257;
  assign n3259 = \encrypt_mode<0>  & n3237;
  assign n3260 = n2528 & n3259;
  assign n3261 = n2523 & n3260;
  assign n3262 = ~\reset<0>  & n3261;
  assign n3263 = ~\encrypt_mode<0>  & n3056;
  assign n3264 = n2528 & n3263;
  assign n3265 = ~n2523 & n3264;
  assign n3266 = ~\reset<0>  & n3265;
  assign n3267 = \encrypt_mode<0>  & n3225;
  assign n3268 = n2528 & n3267;
  assign n3269 = ~n2523 & n3268;
  assign n3270 = ~\reset<0>  & n3269;
  assign n3271 = \inreg<44>  & n2577;
  assign n3272 = ~\reset<0>  & n3271;
  assign n3273 = ~n2528 & n3215;
  assign n3274 = ~\reset<0>  & n3273;
  assign n3275 = \inreg<36>  & n2549;
  assign n3276 = ~\reset<0>  & n3275;
  assign n3277 = ~n3274 & ~n3276;
  assign n3278 = ~n3272 & n3277;
  assign n3279 = ~n3270 & n3278;
  assign n3280 = ~n3266 & n3279;
  assign n3281 = ~n3262 & n3280;
  assign \D_new<17>  = n3258 | ~n3281;
  assign n3283 = n2523 & n3264;
  assign n3284 = ~\reset<0>  & n3283;
  assign n3285 = n2523 & n3232;
  assign n3286 = ~\reset<0>  & n3285;
  assign n3287 = ~n2523 & n3217;
  assign n3288 = ~\reset<0>  & n3287;
  assign n3289 = ~n2523 & n3260;
  assign n3290 = ~\reset<0>  & n3289;
  assign n3291 = \inreg<36>  & n2577;
  assign n3292 = ~\reset<0>  & n3291;
  assign n3293 = ~n2528 & n3225;
  assign n3294 = ~\reset<0>  & n3293;
  assign n3295 = \inreg<28>  & n2549;
  assign n3296 = ~\reset<0>  & n3295;
  assign n3297 = ~n3294 & ~n3296;
  assign n3298 = ~n3292 & n3297;
  assign n3299 = ~n3290 & n3298;
  assign n3300 = ~n3288 & n3299;
  assign n3301 = ~n3286 & n3300;
  assign \D_new<18>  = n3284 | ~n3301;
  assign n3303 = n2523 & n3062;
  assign n3304 = ~\reset<0>  & n3303;
  assign n3305 = \encrypt_mode<0>  & n3215;
  assign n3306 = n2528 & n3305;
  assign n3307 = n2523 & n3306;
  assign n3308 = ~\reset<0>  & n3307;
  assign n3309 = ~\encrypt_mode<0>  & n3036;
  assign n3310 = n2528 & n3309;
  assign n3311 = ~n2523 & n3310;
  assign n3312 = ~\reset<0>  & n3311;
  assign n3313 = ~n2523 & n3058;
  assign n3314 = ~\reset<0>  & n3313;
  assign n3315 = \inreg<52>  & n2549;
  assign n3316 = ~\reset<0>  & n3315;
  assign n3317 = ~n2528 & n3026;
  assign n3318 = ~\reset<0>  & n3317;
  assign n3319 = ~\encrypt<0>  & n3071;
  assign n3320 = ~\reset<0>  & n3319;
  assign n3321 = ~n3318 & ~n3320;
  assign n3322 = ~n3316 & n3321;
  assign n3323 = ~n3314 & n3322;
  assign n3324 = ~n3312 & n3323;
  assign n3325 = ~n3308 & n3324;
  assign \D_new<15>  = n3304 | ~n3325;
  assign n3327 = n2523 & n3310;
  assign n3328 = ~\reset<0>  & n3327;
  assign n3329 = n2523 & n3268;
  assign n3330 = ~\reset<0>  & n3329;
  assign n3331 = ~n2523 & n3256;
  assign n3332 = ~\reset<0>  & n3331;
  assign n3333 = ~n2523 & n3306;
  assign n3334 = ~\reset<0>  & n3333;
  assign n3335 = \inreg<52>  & n2577;
  assign n3336 = ~\reset<0>  & n3335;
  assign n3337 = ~n2528 & n3056;
  assign n3338 = ~\reset<0>  & n3337;
  assign n3339 = \inreg<44>  & n2549;
  assign n3340 = ~\reset<0>  & n3339;
  assign n3341 = ~n3338 & ~n3340;
  assign n3342 = ~n3336 & n3341;
  assign n3343 = ~n3334 & n3342;
  assign n3344 = ~n3332 & n3343;
  assign n3345 = ~n3330 & n3344;
  assign \D_new<16>  = n3328 | ~n3345;
  assign n3347 = ~\encrypt_mode<0>  & n3220;
  assign n3348 = n2528 & n3347;
  assign n3349 = n2523 & n3348;
  assign n3350 = ~\reset<0>  & n3349;
  assign n3351 = \D<25>  & ~n674;
  assign n3352 = \encrypt_mode<0>  & n3351;
  assign n3353 = n2528 & n3352;
  assign n3354 = n2523 & n3353;
  assign n3355 = ~\reset<0>  & n3354;
  assign n3356 = \D<22>  & ~n674;
  assign n3357 = ~\encrypt_mode<0>  & n3356;
  assign n3358 = n2528 & n3357;
  assign n3359 = ~n2523 & n3358;
  assign n3360 = ~\reset<0>  & n3359;
  assign n3361 = \D<24>  & ~n674;
  assign n3362 = \encrypt_mode<0>  & n3361;
  assign n3363 = n2528 & n3362;
  assign n3364 = ~n2523 & n3363;
  assign n3365 = ~\reset<0>  & n3364;
  assign n3366 = \inreg<19>  & n2549;
  assign n3367 = ~\reset<0>  & n3366;
  assign n3368 = \D<23>  & ~n674;
  assign n3369 = ~n2528 & n3368;
  assign n3370 = ~\reset<0>  & n3369;
  assign n3371 = \data_in<4>  & n674;
  assign n3372 = ~\encrypt<0>  & n3371;
  assign n3373 = ~\reset<0>  & n3372;
  assign n3374 = ~n3370 & ~n3373;
  assign n3375 = ~n3367 & n3374;
  assign n3376 = ~n3365 & n3375;
  assign n3377 = ~n3360 & n3376;
  assign n3378 = ~n3355 & n3377;
  assign \D_new<23>  = n3350 | ~n3378;
  assign n3380 = n2523 & n3358;
  assign n3381 = ~\reset<0>  & n3380;
  assign n3382 = \D<26>  & ~n674;
  assign n3383 = \encrypt_mode<0>  & n3382;
  assign n3384 = n2528 & n3383;
  assign n3385 = n2523 & n3384;
  assign n3386 = ~\reset<0>  & n3385;
  assign n3387 = ~\encrypt_mode<0>  & n3368;
  assign n3388 = n2528 & n3387;
  assign n3389 = ~n2523 & n3388;
  assign n3390 = ~\reset<0>  & n3389;
  assign n3391 = ~n2523 & n3353;
  assign n3392 = ~\reset<0>  & n3391;
  assign n3393 = \inreg<19>  & n2577;
  assign n3394 = ~\reset<0>  & n3393;
  assign n3395 = ~n2528 & n3361;
  assign n3396 = ~\reset<0>  & n3395;
  assign n3397 = \inreg<11>  & n2549;
  assign n3398 = ~\reset<0>  & n3397;
  assign n3399 = ~n3396 & ~n3398;
  assign n3400 = ~n3394 & n3399;
  assign n3401 = ~n3392 & n3400;
  assign n3402 = ~n3390 & n3401;
  assign n3403 = ~n3386 & n3402;
  assign \D_new<24>  = n3381 | ~n3403;
  assign n3405 = ~\encrypt_mode<0>  & n3237;
  assign n3406 = n2528 & n3405;
  assign n3407 = n2523 & n3406;
  assign n3408 = ~\reset<0>  & n3407;
  assign n3409 = \encrypt_mode<0>  & n3368;
  assign n3410 = n2528 & n3409;
  assign n3411 = n2523 & n3410;
  assign n3412 = ~\reset<0>  & n3411;
  assign n3413 = ~\encrypt_mode<0>  & n3230;
  assign n3414 = n2528 & n3413;
  assign n3415 = ~n2523 & n3414;
  assign n3416 = ~\reset<0>  & n3415;
  assign n3417 = \encrypt_mode<0>  & n3356;
  assign n3418 = n2528 & n3417;
  assign n3419 = ~n2523 & n3418;
  assign n3420 = ~\reset<0>  & n3419;
  assign n3421 = \inreg<4>  & n2549;
  assign n3422 = ~\reset<0>  & n3421;
  assign n3423 = \inreg<12>  & n2577;
  assign n3424 = ~\reset<0>  & n3423;
  assign n3425 = ~n2528 & n3220;
  assign n3426 = ~\reset<0>  & n3425;
  assign n3427 = ~n3424 & ~n3426;
  assign n3428 = ~n3422 & n3427;
  assign n3429 = ~n3420 & n3428;
  assign n3430 = ~n3416 & n3429;
  assign n3431 = ~n3412 & n3430;
  assign \D_new<21>  = n3408 | ~n3431;
  assign n3433 = n2523 & n3414;
  assign n3434 = ~\reset<0>  & n3433;
  assign n3435 = n2523 & n3363;
  assign n3436 = ~\reset<0>  & n3435;
  assign n3437 = ~n2523 & n3348;
  assign n3438 = ~\reset<0>  & n3437;
  assign n3439 = ~n2523 & n3410;
  assign n3440 = ~\reset<0>  & n3439;
  assign n3441 = \inreg<4>  & n2577;
  assign n3442 = ~\reset<0>  & n3441;
  assign n3443 = ~n2528 & n3356;
  assign n3444 = ~\reset<0>  & n3443;
  assign n3445 = \encrypt<0>  & n3371;
  assign n3446 = ~\reset<0>  & n3445;
  assign n3447 = ~n3444 & ~n3446;
  assign n3448 = ~n3442 & n3447;
  assign n3449 = ~n3440 & n3448;
  assign n3450 = ~n3438 & n3449;
  assign n3451 = ~n3436 & n3450;
  assign \D_new<22>  = n3434 | ~n3451;
  assign n3453 = n2523 & n3227;
  assign n3454 = ~\reset<0>  & n3453;
  assign n3455 = n2523 & n3418;
  assign n3456 = ~\reset<0>  & n3455;
  assign n3457 = ~n2523 & n3406;
  assign n3458 = ~\reset<0>  & n3457;
  assign n3459 = ~n2523 & n3222;
  assign n3460 = ~\reset<0>  & n3459;
  assign n3461 = \inreg<20>  & n2577;
  assign n3462 = ~\reset<0>  & n3461;
  assign n3463 = ~n2528 & n3230;
  assign n3464 = ~\reset<0>  & n3463;
  assign n3465 = \inreg<12>  & n2549;
  assign n3466 = ~\reset<0>  & n3465;
  assign n3467 = ~n3464 & ~n3466;
  assign n3468 = ~n3462 & n3467;
  assign n3469 = ~n3460 & n3468;
  assign n3470 = ~n3458 & n3469;
  assign n3471 = ~n3456 & n3470;
  assign \D_new<20>  = n3454 | ~n3471;
  assign n3473 = \data<21>  & ~n504;
  assign n3474 = n1403 & n3473;
  assign n3475 = ~\data<21>  & ~n504;
  assign n3476 = ~n1403 & n3475;
  assign n3477 = \inreg<12>  & n504;
  assign n3478 = ~n3476 & ~n3477;
  assign \data_new<53>  = n3474 | ~n3478;
  assign n3480 = \data<22>  & ~n504;
  assign n3481 = n817 & n3480;
  assign n3482 = ~\data<22>  & ~n504;
  assign n3483 = ~n817 & n3482;
  assign n3484 = \inreg<4>  & n504;
  assign n3485 = ~n3483 & ~n3484;
  assign \data_new<54>  = n3481 | ~n3485;
  assign n3487 = \data<19>  & ~n504;
  assign n3488 = n2233 & n3487;
  assign n3489 = ~\data<19>  & ~n504;
  assign n3490 = ~n2233 & n3489;
  assign n3491 = \inreg<28>  & n504;
  assign n3492 = ~n3490 & ~n3491;
  assign \data_new<51>  = n3488 | ~n3492;
  assign n3494 = \data<20>  & ~n504;
  assign n3495 = n1543 & n3494;
  assign n3496 = ~\data<20>  & ~n504;
  assign n3497 = ~n1543 & n3496;
  assign n3498 = \inreg<20>  & n504;
  assign n3499 = ~n3497 & ~n3498;
  assign \data_new<52>  = n3495 | ~n3499;
  assign n3501 = \data<18>  & ~n504;
  assign n3502 = n2450 & n3501;
  assign n3503 = ~\data<18>  & ~n504;
  assign n3504 = ~n2450 & n3503;
  assign n3505 = \inreg<36>  & n504;
  assign n3506 = ~n3504 & ~n3505;
  assign \data_new<50>  = n3502 | ~n3506;
  assign n3508 = ~\encrypt_mode<0>  & n3351;
  assign n3509 = n2528 & n3508;
  assign n3510 = n2523 & n3509;
  assign n3511 = ~\reset<0>  & n3510;
  assign n3512 = \D<1>  & ~n674;
  assign n3513 = \encrypt_mode<0>  & n3512;
  assign n3514 = n2528 & n3513;
  assign n3515 = n2523 & n3514;
  assign n3516 = ~\reset<0>  & n3515;
  assign n3517 = ~\encrypt_mode<0>  & n3382;
  assign n3518 = n2528 & n3517;
  assign n3519 = ~n2523 & n3518;
  assign n3520 = ~\reset<0>  & n3519;
  assign n3521 = \D<0>  & ~n674;
  assign n3522 = \encrypt_mode<0>  & n3521;
  assign n3523 = n2528 & n3522;
  assign n3524 = ~n2523 & n3523;
  assign n3525 = ~\reset<0>  & n3524;
  assign n3526 = \inreg<54>  & n2549;
  assign n3527 = ~\reset<0>  & n3526;
  assign n3528 = \D<27>  & ~n674;
  assign n3529 = ~n2528 & n3528;
  assign n3530 = ~\reset<0>  & n3529;
  assign n3531 = \data_in<3>  & n674;
  assign n3532 = ~\encrypt<0>  & n3531;
  assign n3533 = ~\reset<0>  & n3532;
  assign n3534 = ~n3530 & ~n3533;
  assign n3535 = ~n3527 & n3534;
  assign n3536 = ~n3525 & n3535;
  assign n3537 = ~n3520 & n3536;
  assign n3538 = ~n3516 & n3537;
  assign \D_new<27>  = n3511 | ~n3538;
  assign n3540 = n2523 & n3388;
  assign n3541 = ~\reset<0>  & n3540;
  assign n3542 = \encrypt_mode<0>  & n3528;
  assign n3543 = n2528 & n3542;
  assign n3544 = n2523 & n3543;
  assign n3545 = ~\reset<0>  & n3544;
  assign n3546 = ~\encrypt_mode<0>  & n3361;
  assign n3547 = n2528 & n3546;
  assign n3548 = ~n2523 & n3547;
  assign n3549 = ~\reset<0>  & n3548;
  assign n3550 = ~n2523 & n3384;
  assign n3551 = ~\reset<0>  & n3550;
  assign n3552 = \inreg<3>  & n2549;
  assign n3553 = ~\reset<0>  & n3552;
  assign n3554 = \inreg<11>  & n2577;
  assign n3555 = ~\reset<0>  & n3554;
  assign n3556 = ~n2528 & n3351;
  assign n3557 = ~\reset<0>  & n3556;
  assign n3558 = ~n3555 & ~n3557;
  assign n3559 = ~n3553 & n3558;
  assign n3560 = ~n3551 & n3559;
  assign n3561 = ~n3549 & n3560;
  assign n3562 = ~n3545 & n3561;
  assign \D_new<25>  = n3541 | ~n3562;
  assign n3564 = n2523 & n3547;
  assign n3565 = ~\reset<0>  & n3564;
  assign n3566 = n2523 & n3523;
  assign n3567 = ~\reset<0>  & n3566;
  assign n3568 = ~n2523 & n3509;
  assign n3569 = ~\reset<0>  & n3568;
  assign n3570 = ~n2523 & n3543;
  assign n3571 = ~\reset<0>  & n3570;
  assign n3572 = \inreg<3>  & n2577;
  assign n3573 = ~\reset<0>  & n3572;
  assign n3574 = ~n2528 & n3382;
  assign n3575 = ~\reset<0>  & n3574;
  assign n3576 = \encrypt<0>  & n3531;
  assign n3577 = ~\reset<0>  & n3576;
  assign n3578 = ~n3575 & ~n3577;
  assign n3579 = ~n3573 & n3578;
  assign n3580 = ~n3571 & n3579;
  assign n3581 = ~n3569 & n3580;
  assign n3582 = ~n3567 & n3581;
  assign \D_new<26>  = n3565 | ~n3582;
  assign n3584 = \data<27>  & ~n504;
  assign n3585 = n2027 & n3584;
  assign n3586 = ~\data<27>  & ~n504;
  assign n3587 = ~n2027 & n3586;
  assign n3588 = \inreg<30>  & n504;
  assign n3589 = ~n3587 & ~n3588;
  assign \data_new<59>  = n3585 | ~n3589;
  assign n3591 = ~n2104 & n2147;
  assign n3592 = ~n2104 & n2150;
  assign n3593 = ~n2104 & n2156;
  assign n3594 = ~n2107 & n2155;
  assign n3595 = n2104 & n3594;
  assign n3596 = n2107 & n2140;
  assign n3597 = n2104 & n3596;
  assign n3598 = n2107 & n2143;
  assign n3599 = n2104 & n3598;
  assign n3600 = ~n2104 & n2185;
  assign n3601 = ~n2104 & n2188;
  assign n3602 = ~n2104 & n2192;
  assign n3603 = n2107 & n2187;
  assign n3604 = n2104 & n3603;
  assign n3605 = ~n2110 & n2172;
  assign n3606 = ~n2107 & n3605;
  assign n3607 = n2104 & n3606;
  assign n3608 = n2107 & n3605;
  assign n3609 = n2104 & n3608;
  assign n3610 = n2107 & n2165;
  assign n3611 = n2104 & n3610;
  assign n3612 = n2107 & n2122;
  assign n3613 = n2104 & n3612;
  assign n3614 = ~n2104 & n2194;
  assign n3615 = ~n2193 & ~n2195;
  assign n3616 = ~n3609 & n3615;
  assign n3617 = ~n3607 & n3616;
  assign n3618 = ~n3604 & n3617;
  assign n3619 = ~n2189 & n3618;
  assign n3620 = ~n2186 & n3619;
  assign n3621 = ~n2184 & n3620;
  assign n3622 = ~n3602 & n3621;
  assign n3623 = ~n2175 & n3622;
  assign n3624 = ~n2167 & n3623;
  assign n3625 = ~n3601 & n3624;
  assign n3626 = ~n2163 & n3625;
  assign n3627 = ~n3600 & n3626;
  assign n3628 = ~n3599 & n3627;
  assign n3629 = ~n3597 & n3628;
  assign n3630 = ~n2157 & n3629;
  assign n3631 = ~n3595 & n3630;
  assign n3632 = ~n2153 & n3631;
  assign n3633 = ~n2151 & n3632;
  assign n3634 = ~n2148 & n3633;
  assign n3635 = ~n2145 & n3634;
  assign n3636 = ~n3593 & n3635;
  assign n3637 = ~n2138 & n3636;
  assign n3638 = ~n3592 & n3637;
  assign n3639 = ~n3591 & n3638;
  assign n3640 = ~n2129 & n3639;
  assign n3641 = ~n2124 & n3640;
  assign n3642 = ~n2104 & n2152;
  assign n3643 = n3641 & ~n3642;
  assign n3644 = ~n3614 & n3643;
  assign n3645 = ~n3613 & n3644;
  assign n3646 = ~n3611 & n3645;
  assign n3647 = \data<25>  & ~n504;
  assign n3648 = n3646 & n3647;
  assign n3649 = ~\data<25>  & ~n504;
  assign n3650 = ~n3646 & n3649;
  assign n3651 = \inreg<46>  & n504;
  assign n3652 = ~n3650 & ~n3651;
  assign \data_new<57>  = n3648 | ~n3652;
  assign n3654 = \data<26>  & ~n504;
  assign n3655 = n2499 & n3654;
  assign n3656 = ~\data<26>  & ~n504;
  assign n3657 = ~n2499 & n3656;
  assign n3658 = \inreg<38>  & n504;
  assign n3659 = ~n3657 & ~n3658;
  assign \data_new<58>  = n3655 | ~n3659;
  assign n3661 = ~n1117 & n1160;
  assign n3662 = n1117 & n1142;
  assign n3663 = ~n1117 & n1199;
  assign n3664 = n1117 & n1183;
  assign n3665 = n1117 & n1420;
  assign n3666 = n1117 & n1246;
  assign n3667 = ~n1117 & n1165;
  assign n3668 = ~n1214 & ~n1433;
  assign n3669 = ~n1432 & n3668;
  assign n3670 = ~n1210 & n3669;
  assign n3671 = ~n1205 & n3670;
  assign n3672 = ~n3664 & n3671;
  assign n3673 = ~n1200 & n3672;
  assign n3674 = ~n1198 & n3673;
  assign n3675 = ~n1193 & n3674;
  assign n3676 = ~n1429 & n3675;
  assign n3677 = ~n1428 & n3676;
  assign n3678 = ~n3663 & n3677;
  assign n3679 = ~n1180 & n3678;
  assign n3680 = ~n1177 & n3679;
  assign n3681 = ~n1172 & n3680;
  assign n3682 = ~n1169 & n3681;
  assign n3683 = ~n1167 & n3682;
  assign n3684 = ~n1164 & n3683;
  assign n3685 = ~n3662 & n3684;
  assign n3686 = ~n1426 & n3685;
  assign n3687 = ~n1425 & n3686;
  assign n3688 = ~n1423 & n3687;
  assign n3689 = ~n1158 & n3688;
  assign n3690 = ~n1154 & n3689;
  assign n3691 = ~n1146 & n3690;
  assign n3692 = ~n1419 & n3691;
  assign n3693 = ~n1139 & n3692;
  assign n3694 = ~n3661 & n3693;
  assign n3695 = ~n1117 & n1204;
  assign n3696 = n3694 & ~n3695;
  assign n3697 = ~n3667 & n3696;
  assign n3698 = ~n3666 & n3697;
  assign n3699 = ~n3665 & n3698;
  assign n3700 = \data<23>  & ~n504;
  assign n3701 = n3699 & n3700;
  assign n3702 = ~\data<23>  & ~n504;
  assign n3703 = ~n3699 & n3702;
  assign n3704 = \data_in<4>  & n504;
  assign n3705 = ~n3703 & ~n3704;
  assign \data_new<55>  = n3701 | ~n3705;
  assign n3707 = ~n880 & n924;
  assign n3708 = n880 & n2263;
  assign n3709 = ~n880 & n967;
  assign n3710 = n880 & n953;
  assign n3711 = n880 & n960;
  assign n3712 = ~n883 & n977;
  assign n3713 = n880 & n3712;
  assign n3714 = ~n880 & n980;
  assign n3715 = ~n880 & n932;
  assign n3716 = ~n974 & ~n3710;
  assign n3717 = ~n2260 & n3716;
  assign n3718 = ~n972 & n3717;
  assign n3719 = ~n2259 & n3718;
  assign n3720 = ~n968 & n3719;
  assign n3721 = ~n963 & n3720;
  assign n3722 = ~n961 & n3721;
  assign n3723 = ~n2257 & n3722;
  assign n3724 = ~n954 & n3723;
  assign n3725 = ~n943 & n3724;
  assign n3726 = ~n3709 & n3725;
  assign n3727 = ~n2256 & n3726;
  assign n3728 = ~n939 & n3727;
  assign n3729 = ~n2253 & n3728;
  assign n3730 = ~n3708 & n3729;
  assign n3731 = ~n933 & n3730;
  assign n3732 = ~n931 & n3731;
  assign n3733 = ~n925 & n3732;
  assign n3734 = ~n2251 & n3733;
  assign n3735 = ~n922 & n3734;
  assign n3736 = ~n2250 & n3735;
  assign n3737 = ~n918 & n3736;
  assign n3738 = ~n914 & n3737;
  assign n3739 = ~n906 & n3738;
  assign n3740 = ~n904 & n3739;
  assign n3741 = ~n3707 & n3740;
  assign n3742 = ~n2248 & n3741;
  assign n3743 = ~n3715 & n3742;
  assign n3744 = ~n3714 & n3743;
  assign n3745 = ~n3713 & n3744;
  assign n3746 = ~n3711 & n3745;
  assign n3747 = \data<24>  & ~n504;
  assign n3748 = n3746 & n3747;
  assign n3749 = ~\data<24>  & ~n504;
  assign n3750 = ~n3746 & n3749;
  assign n3751 = \inreg<54>  & n504;
  assign n3752 = ~n3750 & ~n3751;
  assign \data_new<56>  = n3748 | ~n3752;
  assign n3754 = \D<5>  & ~n674;
  assign n3755 = ~\encrypt_mode<0>  & n3754;
  assign n3756 = n2528 & n3755;
  assign n3757 = n2523 & n3756;
  assign n3758 = ~\reset<0>  & n3757;
  assign n3759 = \encrypt_mode<0>  & n3080;
  assign n3760 = n2528 & n3759;
  assign n3761 = n2523 & n3760;
  assign n3762 = ~\reset<0>  & n3761;
  assign n3763 = \D<6>  & ~n674;
  assign n3764 = ~\encrypt_mode<0>  & n3763;
  assign n3765 = n2528 & n3764;
  assign n3766 = ~n2523 & n3765;
  assign n3767 = ~\reset<0>  & n3766;
  assign n3768 = \encrypt_mode<0>  & n3130;
  assign n3769 = n2528 & n3768;
  assign n3770 = ~n2523 & n3769;
  assign n3771 = ~\reset<0>  & n3770;
  assign n3772 = \inreg<53>  & n2549;
  assign n3773 = ~\reset<0>  & n3772;
  assign n3774 = \D<7>  & ~n674;
  assign n3775 = ~n2528 & n3774;
  assign n3776 = ~\reset<0>  & n3775;
  assign n3777 = \data_in<6>  & n674;
  assign n3778 = ~\encrypt<0>  & n3777;
  assign n3779 = ~\reset<0>  & n3778;
  assign n3780 = ~n3776 & ~n3779;
  assign n3781 = ~n3773 & n3780;
  assign n3782 = ~n3771 & n3781;
  assign n3783 = ~n3767 & n3782;
  assign n3784 = ~n3762 & n3783;
  assign \D_new<7>  = n3758 | ~n3784;
  assign n3786 = \C<4>  & ~n674;
  assign n3787 = ~\encrypt_mode<0>  & n3786;
  assign n3788 = n2528 & n3787;
  assign n3789 = n2523 & n3788;
  assign n3790 = ~\reset<0>  & n3789;
  assign n3791 = \encrypt_mode<0>  & n2864;
  assign n3792 = n2528 & n3791;
  assign n3793 = n2523 & n3792;
  assign n3794 = ~\reset<0>  & n3793;
  assign n3795 = \C<5>  & ~n674;
  assign n3796 = ~\encrypt_mode<0>  & n3795;
  assign n3797 = n2528 & n3796;
  assign n3798 = ~n2523 & n3797;
  assign n3799 = ~\reset<0>  & n3798;
  assign n3800 = \C<7>  & ~n674;
  assign n3801 = \encrypt_mode<0>  & n3800;
  assign n3802 = n2528 & n3801;
  assign n3803 = ~n2523 & n3802;
  assign n3804 = ~\reset<0>  & n3803;
  assign n3805 = \inreg<0>  & n2577;
  assign n3806 = ~\reset<0>  & n3805;
  assign n3807 = \C<6>  & ~n674;
  assign n3808 = ~n2528 & n3807;
  assign n3809 = ~\reset<0>  & n3808;
  assign n3810 = \data_in<0>  & n674;
  assign n3811 = \encrypt<0>  & n3810;
  assign n3812 = ~\reset<0>  & n3811;
  assign n3813 = ~n3809 & ~n3812;
  assign n3814 = ~n3806 & n3813;
  assign n3815 = ~n3804 & n3814;
  assign n3816 = ~n3799 & n3815;
  assign n3817 = ~n3794 & n3816;
  assign \C_new<6>  = n3790 | ~n3817;
  assign n3819 = n2523 & n3765;
  assign n3820 = ~\reset<0>  & n3819;
  assign n3821 = \encrypt_mode<0>  & n3089;
  assign n3822 = n2528 & n3821;
  assign n3823 = n2523 & n3822;
  assign n3824 = ~\reset<0>  & n3823;
  assign n3825 = ~\encrypt_mode<0>  & n3774;
  assign n3826 = n2528 & n3825;
  assign n3827 = ~n2523 & n3826;
  assign n3828 = ~\reset<0>  & n3827;
  assign n3829 = ~n2523 & n3760;
  assign n3830 = ~\reset<0>  & n3829;
  assign n3831 = \inreg<53>  & n2577;
  assign n3832 = ~\reset<0>  & n3831;
  assign n3833 = ~n2528 & n3130;
  assign n3834 = ~\reset<0>  & n3833;
  assign n3835 = \inreg<45>  & n2549;
  assign n3836 = ~\reset<0>  & n3835;
  assign n3837 = ~n3834 & ~n3836;
  assign n3838 = ~n3832 & n3837;
  assign n3839 = ~n3830 & n3838;
  assign n3840 = ~n3828 & n3839;
  assign n3841 = ~n3824 & n3840;
  assign \D_new<8>  = n3820 | ~n3841;
  assign n3843 = \C<3>  & ~n674;
  assign n3844 = ~\encrypt_mode<0>  & n3843;
  assign n3845 = n2528 & n3844;
  assign n3846 = n2523 & n3845;
  assign n3847 = ~\reset<0>  & n3846;
  assign n3848 = n2523 & n3802;
  assign n3849 = ~\reset<0>  & n3848;
  assign n3850 = ~n2523 & n3788;
  assign n3851 = ~\reset<0>  & n3850;
  assign n3852 = \encrypt_mode<0>  & n3807;
  assign n3853 = n2528 & n3852;
  assign n3854 = ~n2523 & n3853;
  assign n3855 = ~\reset<0>  & n3854;
  assign n3856 = \inreg<8>  & n2577;
  assign n3857 = ~\reset<0>  & n3856;
  assign n3858 = ~n2528 & n3795;
  assign n3859 = ~\reset<0>  & n3858;
  assign n3860 = \inreg<0>  & n2549;
  assign n3861 = ~\reset<0>  & n3860;
  assign n3862 = ~n3859 & ~n3861;
  assign n3863 = ~n3857 & n3862;
  assign n3864 = ~n3855 & n3863;
  assign n3865 = ~n3851 & n3864;
  assign n3866 = ~n3849 & n3865;
  assign \C_new<5>  = n3847 | ~n3866;
  assign n3868 = \D<3>  & ~n674;
  assign n3869 = ~\encrypt_mode<0>  & n3868;
  assign n3870 = n2528 & n3869;
  assign n3871 = n2523 & n3870;
  assign n3872 = ~\reset<0>  & n3871;
  assign n3873 = \encrypt_mode<0>  & n3774;
  assign n3874 = n2528 & n3873;
  assign n3875 = n2523 & n3874;
  assign n3876 = ~\reset<0>  & n3875;
  assign n3877 = \D<4>  & ~n674;
  assign n3878 = ~\encrypt_mode<0>  & n3877;
  assign n3879 = n2528 & n3878;
  assign n3880 = ~n2523 & n3879;
  assign n3881 = ~\reset<0>  & n3880;
  assign n3882 = \encrypt_mode<0>  & n3763;
  assign n3883 = n2528 & n3882;
  assign n3884 = ~n2523 & n3883;
  assign n3885 = ~\reset<0>  & n3884;
  assign n3886 = \inreg<6>  & n2549;
  assign n3887 = ~\reset<0>  & n3886;
  assign n3888 = \inreg<14>  & n2577;
  assign n3889 = ~\reset<0>  & n3888;
  assign n3890 = ~n2528 & n3754;
  assign n3891 = ~\reset<0>  & n3890;
  assign n3892 = ~n3889 & ~n3891;
  assign n3893 = ~n3887 & n3892;
  assign n3894 = ~n3885 & n3893;
  assign n3895 = ~n3881 & n3894;
  assign n3896 = ~n3876 & n3895;
  assign \D_new<5>  = n3872 | ~n3896;
  assign n3898 = ~\encrypt_mode<0>  & n3807;
  assign n3899 = n2528 & n3898;
  assign n3900 = n2523 & n3899;
  assign n3901 = ~\reset<0>  & n3900;
  assign n3902 = \encrypt_mode<0>  & n2823;
  assign n3903 = n2528 & n3902;
  assign n3904 = n2523 & n3903;
  assign n3905 = ~\reset<0>  & n3904;
  assign n3906 = ~\encrypt_mode<0>  & n3800;
  assign n3907 = n2528 & n3906;
  assign n3908 = ~n2523 & n3907;
  assign n3909 = ~\reset<0>  & n3908;
  assign n3910 = \encrypt_mode<0>  & n2814;
  assign n3911 = n2528 & n3910;
  assign n3912 = ~n2523 & n3911;
  assign n3913 = ~\reset<0>  & n3912;
  assign n3914 = \inreg<49>  & n2577;
  assign n3915 = ~\reset<0>  & n3914;
  assign n3916 = ~n2528 & n2864;
  assign n3917 = ~\reset<0>  & n3916;
  assign n3918 = \inreg<41>  & n2549;
  assign n3919 = ~\reset<0>  & n3918;
  assign n3920 = ~n3917 & ~n3919;
  assign n3921 = ~n3915 & n3920;
  assign n3922 = ~n3913 & n3921;
  assign n3923 = ~n3909 & n3922;
  assign n3924 = ~n3905 & n3923;
  assign \C_new<8>  = n3901 | ~n3924;
  assign n3926 = n2523 & n3879;
  assign n3927 = ~\reset<0>  & n3926;
  assign n3928 = n2523 & n3769;
  assign n3929 = ~\reset<0>  & n3928;
  assign n3930 = ~n2523 & n3756;
  assign n3931 = ~\reset<0>  & n3930;
  assign n3932 = ~n2523 & n3874;
  assign n3933 = ~\reset<0>  & n3932;
  assign n3934 = \inreg<6>  & n2577;
  assign n3935 = ~\reset<0>  & n3934;
  assign n3936 = ~n2528 & n3763;
  assign n3937 = ~\reset<0>  & n3936;
  assign n3938 = \encrypt<0>  & n3777;
  assign n3939 = ~\reset<0>  & n3938;
  assign n3940 = ~n3937 & ~n3939;
  assign n3941 = ~n3935 & n3940;
  assign n3942 = ~n3933 & n3941;
  assign n3943 = ~n3931 & n3942;
  assign n3944 = ~n3929 & n3943;
  assign \D_new<6>  = n3927 | ~n3944;
  assign n3946 = n2523 & n3797;
  assign n3947 = ~\reset<0>  & n3946;
  assign n3948 = n2523 & n3911;
  assign n3949 = ~\reset<0>  & n3948;
  assign n3950 = ~n2523 & n3899;
  assign n3951 = ~\reset<0>  & n3950;
  assign n3952 = ~n2523 & n3792;
  assign n3953 = ~\reset<0>  & n3952;
  assign n3954 = \inreg<49>  & n2549;
  assign n3955 = ~\reset<0>  & n3954;
  assign n3956 = ~n2528 & n3800;
  assign n3957 = ~\reset<0>  & n3956;
  assign n3958 = ~\encrypt<0>  & n3810;
  assign n3959 = ~\reset<0>  & n3958;
  assign n3960 = ~n3957 & ~n3959;
  assign n3961 = ~n3955 & n3960;
  assign n3962 = ~n3953 & n3961;
  assign n3963 = ~n3951 & n3962;
  assign n3964 = ~n3949 & n3963;
  assign \C_new<7>  = n3947 | ~n3964;
  assign n3966 = n2523 & n3907;
  assign n3967 = ~\reset<0>  & n3966;
  assign n3968 = n2523 & n2874;
  assign n3969 = ~\reset<0>  & n3968;
  assign n3970 = ~n2523 & n2866;
  assign n3971 = ~\reset<0>  & n3970;
  assign n3972 = ~n2523 & n3903;
  assign n3973 = ~\reset<0>  & n3972;
  assign n3974 = \inreg<41>  & n2577;
  assign n3975 = ~\reset<0>  & n3974;
  assign n3976 = ~n2528 & n2814;
  assign n3977 = ~\reset<0>  & n3976;
  assign n3978 = \inreg<33>  & n2549;
  assign n3979 = ~\reset<0>  & n3978;
  assign n3980 = ~n3977 & ~n3979;
  assign n3981 = ~n3975 & n3980;
  assign n3982 = ~n3973 & n3981;
  assign n3983 = ~n3971 & n3982;
  assign n3984 = ~n3969 & n3983;
  assign \C_new<9>  = n3967 | ~n3984;
  assign n3986 = n2523 & n3826;
  assign n3987 = ~\reset<0>  & n3986;
  assign n3988 = n2523 & n3140;
  assign n3989 = ~\reset<0>  & n3988;
  assign n3990 = ~n2523 & n3132;
  assign n3991 = ~\reset<0>  & n3990;
  assign n3992 = ~n2523 & n3822;
  assign n3993 = ~\reset<0>  & n3992;
  assign n3994 = \inreg<45>  & n2577;
  assign n3995 = ~\reset<0>  & n3994;
  assign n3996 = ~n2528 & n3080;
  assign n3997 = ~\reset<0>  & n3996;
  assign n3998 = \inreg<37>  & n2549;
  assign n3999 = ~\reset<0>  & n3998;
  assign n4000 = ~n3997 & ~n3999;
  assign n4001 = ~n3995 & n4000;
  assign n4002 = ~n3993 & n4001;
  assign n4003 = ~n3991 & n4002;
  assign n4004 = ~n3989 & n4003;
  assign \D_new<9>  = n3987 | ~n4004;
  assign n4006 = n2523 & n3518;
  assign n4007 = ~\reset<0>  & n4006;
  assign n4008 = \D<2>  & ~n674;
  assign n4009 = \encrypt_mode<0>  & n4008;
  assign n4010 = n2528 & n4009;
  assign n4011 = n2523 & n4010;
  assign n4012 = ~\reset<0>  & n4011;
  assign n4013 = ~\encrypt_mode<0>  & n3528;
  assign n4014 = n2528 & n4013;
  assign n4015 = ~n2523 & n4014;
  assign n4016 = ~\reset<0>  & n4015;
  assign n4017 = ~n2523 & n3514;
  assign n4018 = ~\reset<0>  & n4017;
  assign n4019 = \inreg<54>  & n2577;
  assign n4020 = ~\reset<0>  & n4019;
  assign n4021 = ~n2528 & n3521;
  assign n4022 = ~\reset<0>  & n4021;
  assign n4023 = \inreg<46>  & n2549;
  assign n4024 = ~\reset<0>  & n4023;
  assign n4025 = ~n4022 & ~n4024;
  assign n4026 = ~n4020 & n4025;
  assign n4027 = ~n4018 & n4026;
  assign n4028 = ~n4016 & n4027;
  assign n4029 = ~n4012 & n4028;
  assign \D_new<0>  = n4007 | ~n4029;
  assign n4031 = n2523 & n2681;
  assign n4032 = ~\reset<0>  & n4031;
  assign n4033 = \C<2>  & ~n674;
  assign n4034 = \encrypt_mode<0>  & n4033;
  assign n4035 = n2528 & n4034;
  assign n4036 = n2523 & n4035;
  assign n4037 = ~\reset<0>  & n4036;
  assign n4038 = ~\encrypt_mode<0>  & n2693;
  assign n4039 = n2528 & n4038;
  assign n4040 = ~n2523 & n4039;
  assign n4041 = ~\reset<0>  & n4040;
  assign n4042 = ~n2523 & n2677;
  assign n4043 = ~\reset<0>  & n4042;
  assign n4044 = \inreg<48>  & n2577;
  assign n4045 = ~\reset<0>  & n4044;
  assign n4046 = ~n2528 & n2684;
  assign n4047 = ~\reset<0>  & n4046;
  assign n4048 = \inreg<40>  & n2549;
  assign n4049 = ~\reset<0>  & n4048;
  assign n4050 = ~n4047 & ~n4049;
  assign n4051 = ~n4045 & n4050;
  assign n4052 = ~n4043 & n4051;
  assign n4053 = ~n4041 & n4052;
  assign n4054 = ~n4037 & n4053;
  assign \C_new<0>  = n4032 | ~n4054;
  assign n4056 = ~\encrypt_mode<0>  & n3512;
  assign n4057 = n2528 & n4056;
  assign n4058 = n2523 & n4057;
  assign n4059 = ~\reset<0>  & n4058;
  assign n4060 = \encrypt_mode<0>  & n3754;
  assign n4061 = n2528 & n4060;
  assign n4062 = n2523 & n4061;
  assign n4063 = ~\reset<0>  & n4062;
  assign n4064 = ~\encrypt_mode<0>  & n4008;
  assign n4065 = n2528 & n4064;
  assign n4066 = ~n2523 & n4065;
  assign n4067 = ~\reset<0>  & n4066;
  assign n4068 = \encrypt_mode<0>  & n3877;
  assign n4069 = n2528 & n4068;
  assign n4070 = ~n2523 & n4069;
  assign n4071 = ~\reset<0>  & n4070;
  assign n4072 = \inreg<30>  & n2577;
  assign n4073 = ~\reset<0>  & n4072;
  assign n4074 = ~n2528 & n3868;
  assign n4075 = ~\reset<0>  & n4074;
  assign n4076 = \inreg<22>  & n2549;
  assign n4077 = ~\reset<0>  & n4076;
  assign n4078 = ~n4075 & ~n4077;
  assign n4079 = ~n4073 & n4078;
  assign n4080 = ~n4071 & n4079;
  assign n4081 = ~n4067 & n4080;
  assign n4082 = ~n4063 & n4081;
  assign \D_new<3>  = n4059 | ~n4082;
  assign n4084 = ~\encrypt_mode<0>  & n2684;
  assign n4085 = n2528 & n4084;
  assign n4086 = n2523 & n4085;
  assign n4087 = ~\reset<0>  & n4086;
  assign n4088 = \encrypt_mode<0>  & n3786;
  assign n4089 = n2528 & n4088;
  assign n4090 = n2523 & n4089;
  assign n4091 = ~\reset<0>  & n4090;
  assign n4092 = ~\encrypt_mode<0>  & n2675;
  assign n4093 = n2528 & n4092;
  assign n4094 = ~n2523 & n4093;
  assign n4095 = ~\reset<0>  & n4094;
  assign n4096 = \encrypt_mode<0>  & n3843;
  assign n4097 = n2528 & n4096;
  assign n4098 = ~n2523 & n4097;
  assign n4099 = ~\reset<0>  & n4098;
  assign n4100 = \inreg<32>  & n2577;
  assign n4101 = ~\reset<0>  & n4100;
  assign n4102 = ~n2528 & n4033;
  assign n4103 = ~\reset<0>  & n4102;
  assign n4104 = \inreg<24>  & n2549;
  assign n4105 = ~\reset<0>  & n4104;
  assign n4106 = ~n4103 & ~n4105;
  assign n4107 = ~n4101 & n4106;
  assign n4108 = ~n4099 & n4107;
  assign n4109 = ~n4095 & n4108;
  assign n4110 = ~n4091 & n4109;
  assign \C_new<2>  = n4087 | ~n4110;
  assign n4112 = n2523 & n4065;
  assign n4113 = ~\reset<0>  & n4112;
  assign n4114 = n2523 & n3883;
  assign n4115 = ~\reset<0>  & n4114;
  assign n4116 = ~n2523 & n3870;
  assign n4117 = ~\reset<0>  & n4116;
  assign n4118 = ~n2523 & n4061;
  assign n4119 = ~\reset<0>  & n4118;
  assign n4120 = \inreg<22>  & n2577;
  assign n4121 = ~\reset<0>  & n4120;
  assign n4122 = ~n2528 & n3877;
  assign n4123 = ~\reset<0>  & n4122;
  assign n4124 = \inreg<14>  & n2549;
  assign n4125 = ~\reset<0>  & n4124;
  assign n4126 = ~n4123 & ~n4125;
  assign n4127 = ~n4121 & n4126;
  assign n4128 = ~n4119 & n4127;
  assign n4129 = ~n4117 & n4128;
  assign n4130 = ~n4115 & n4129;
  assign \D_new<4>  = n4113 | ~n4130;
  assign n4132 = n2523 & n4039;
  assign n4133 = ~\reset<0>  & n4132;
  assign n4134 = n2523 & n4097;
  assign n4135 = ~\reset<0>  & n4134;
  assign n4136 = ~n2523 & n4085;
  assign n4137 = ~\reset<0>  & n4136;
  assign n4138 = ~n2523 & n4035;
  assign n4139 = ~\reset<0>  & n4138;
  assign n4140 = \inreg<40>  & n2577;
  assign n4141 = ~\reset<0>  & n4140;
  assign n4142 = ~n2528 & n2675;
  assign n4143 = ~\reset<0>  & n4142;
  assign n4144 = \inreg<32>  & n2549;
  assign n4145 = ~\reset<0>  & n4144;
  assign n4146 = ~n4143 & ~n4145;
  assign n4147 = ~n4141 & n4146;
  assign n4148 = ~n4139 & n4147;
  assign n4149 = ~n4137 & n4148;
  assign n4150 = ~n4135 & n4149;
  assign \C_new<1>  = n4133 | ~n4150;
  assign n4152 = n2523 & n4014;
  assign n4153 = ~\reset<0>  & n4152;
  assign n4154 = \encrypt_mode<0>  & n3868;
  assign n4155 = n2528 & n4154;
  assign n4156 = n2523 & n4155;
  assign n4157 = ~\reset<0>  & n4156;
  assign n4158 = ~\encrypt_mode<0>  & n3521;
  assign n4159 = n2528 & n4158;
  assign n4160 = ~n2523 & n4159;
  assign n4161 = ~\reset<0>  & n4160;
  assign n4162 = ~n2523 & n4010;
  assign n4163 = ~\reset<0>  & n4162;
  assign n4164 = \inreg<46>  & n2577;
  assign n4165 = ~\reset<0>  & n4164;
  assign n4166 = ~n2528 & n3512;
  assign n4167 = ~\reset<0>  & n4166;
  assign n4168 = \inreg<38>  & n2549;
  assign n4169 = ~\reset<0>  & n4168;
  assign n4170 = ~n4167 & ~n4169;
  assign n4171 = ~n4165 & n4170;
  assign n4172 = ~n4163 & n4171;
  assign n4173 = ~n4161 & n4172;
  assign n4174 = ~n4157 & n4173;
  assign \D_new<1>  = n4153 | ~n4174;
  assign n4176 = ~\encrypt_mode<0>  & n4033;
  assign n4177 = n2528 & n4176;
  assign n4178 = n2523 & n4177;
  assign n4179 = ~\reset<0>  & n4178;
  assign n4180 = n2523 & n3853;
  assign n4181 = ~\reset<0>  & n4180;
  assign n4182 = ~n2523 & n3845;
  assign n4183 = ~\reset<0>  & n4182;
  assign n4184 = \encrypt_mode<0>  & n3795;
  assign n4185 = n2528 & n4184;
  assign n4186 = ~n2523 & n4185;
  assign n4187 = ~\reset<0>  & n4186;
  assign n4188 = \inreg<8>  & n2549;
  assign n4189 = ~\reset<0>  & n4188;
  assign n4190 = \inreg<16>  & n2577;
  assign n4191 = ~\reset<0>  & n4190;
  assign n4192 = ~n2528 & n3786;
  assign n4193 = ~\reset<0>  & n4192;
  assign n4194 = ~n4191 & ~n4193;
  assign n4195 = ~n4189 & n4194;
  assign n4196 = ~n4187 & n4195;
  assign n4197 = ~n4183 & n4196;
  assign n4198 = ~n4181 & n4197;
  assign \C_new<4>  = n4179 | ~n4198;
  assign n4200 = n2523 & n4159;
  assign n4201 = ~\reset<0>  & n4200;
  assign n4202 = n2523 & n4069;
  assign n4203 = ~\reset<0>  & n4202;
  assign n4204 = ~n2523 & n4057;
  assign n4205 = ~\reset<0>  & n4204;
  assign n4206 = ~n2523 & n4155;
  assign n4207 = ~\reset<0>  & n4206;
  assign n4208 = \inreg<38>  & n2577;
  assign n4209 = ~\reset<0>  & n4208;
  assign n4210 = ~n2528 & n4008;
  assign n4211 = ~\reset<0>  & n4210;
  assign n4212 = \inreg<30>  & n2549;
  assign n4213 = ~\reset<0>  & n4212;
  assign n4214 = ~n4211 & ~n4213;
  assign n4215 = ~n4209 & n4214;
  assign n4216 = ~n4207 & n4215;
  assign n4217 = ~n4205 & n4216;
  assign n4218 = ~n4203 & n4217;
  assign \D_new<2>  = n4201 | ~n4218;
  assign n4220 = n2523 & n4093;
  assign n4221 = ~\reset<0>  & n4220;
  assign n4222 = n2523 & n4185;
  assign n4223 = ~\reset<0>  & n4222;
  assign n4224 = ~n2523 & n4177;
  assign n4225 = ~\reset<0>  & n4224;
  assign n4226 = ~n2523 & n4089;
  assign n4227 = ~\reset<0>  & n4226;
  assign n4228 = \inreg<24>  & n2577;
  assign n4229 = ~\reset<0>  & n4228;
  assign n4230 = ~n2528 & n3843;
  assign n4231 = ~\reset<0>  & n4230;
  assign n4232 = \inreg<16>  & n2549;
  assign n4233 = ~\reset<0>  & n4232;
  assign n4234 = ~n4231 & ~n4233;
  assign n4235 = ~n4229 & n4234;
  assign n4236 = ~n4227 & n4235;
  assign n4237 = ~n4225 & n4236;
  assign n4238 = ~n4223 & n4237;
  assign \C_new<3>  = n4221 | ~n4238;
  assign n4240 = \inreg<50>  & n508;
  assign n4241 = \inreg<42>  & n510;
  assign \inreg_new<50>  = n4240 | n4241;
  assign n4243 = \inreg<9>  & n508;
  assign n4244 = \inreg<1>  & n510;
  assign \inreg_new<9>  = n4243 | n4244;
  assign n4246 = \inreg<54>  & n508;
  assign n4247 = \inreg<46>  & n510;
  assign \inreg_new<54>  = n4246 | n4247;
  assign n4249 = \inreg<53>  & n508;
  assign n4250 = \inreg<45>  & n510;
  assign \inreg_new<53>  = n4249 | n4250;
  assign n4252 = \inreg<52>  & n508;
  assign n4253 = \inreg<44>  & n510;
  assign \inreg_new<52>  = n4252 | n4253;
  assign n4255 = \inreg<6>  & n508;
  assign n4256 = \data_in<6>  & n510;
  assign \inreg_new<6>  = n4255 | n4256;
  assign n4258 = \inreg<51>  & n508;
  assign n4259 = \inreg<43>  & n510;
  assign \inreg_new<51>  = n4258 | n4259;
  assign n4261 = \inreg<5>  & n508;
  assign n4262 = \data_in<5>  & n510;
  assign \inreg_new<5>  = n4261 | n4262;
  assign n4264 = \inreg<8>  & n508;
  assign n4265 = \inreg<0>  & n510;
  assign \inreg_new<8>  = n4264 | n4265;
  assign n4267 = \inreg<7>  & n508;
  assign n4268 = \data_in<7>  & n510;
  assign \inreg_new<7>  = n4267 | n4268;
  assign n4270 = \inreg<2>  & n508;
  assign n4271 = \data_in<2>  & n510;
  assign \inreg_new<2>  = n4270 | n4271;
  assign n4273 = \inreg<55>  & n508;
  assign n4274 = \inreg<47>  & n510;
  assign \inreg_new<55>  = n4273 | n4274;
  assign n4276 = \inreg<1>  & n508;
  assign n4277 = \data_in<1>  & n510;
  assign \inreg_new<1>  = n4276 | n4277;
  assign n4279 = \inreg<4>  & n508;
  assign n4280 = \data_in<4>  & n510;
  assign \inreg_new<4>  = n4279 | n4280;
  assign n4282 = \inreg<3>  & n508;
  assign n4283 = \data_in<3>  & n510;
  assign \inreg_new<3>  = n4282 | n4283;
  assign n4285 = \inreg<0>  & n508;
  assign n4286 = \data_in<0>  & n510;
  assign \inreg_new<0>  = n4285 | n4286;
  assign n4288 = \count<0>  & \encrypt<0> ;
  assign n4289 = \count<1>  & n4288;
  assign n4290 = \count<2>  & n4289;
  assign n4291 = \count<3>  & n4290;
  assign n4292 = ~\count<3>  & \encrypt_mode<0> ;
  assign n4293 = ~\count<2>  & \encrypt_mode<0> ;
  assign n4294 = ~\count<1>  & \encrypt_mode<0> ;
  assign n4295 = ~\count<0>  & \encrypt_mode<0> ;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = ~n4293 & n4296;
  assign n4298 = ~n4292 & n4297;
  assign \encrypt_mode_new<0>  = n4291 | ~n4298;
  assign n4300 = n1271 & n1310;
  assign n4301 = n1271 & n1330;
  assign n4302 = ~n1271 & n2041;
  assign n4303 = ~n1361 & ~n1365;
  assign n4304 = ~n2052 & n4303;
  assign n4305 = ~n1358 & n4304;
  assign n4306 = ~n3159 & n4305;
  assign n4307 = ~n1357 & n4306;
  assign n4308 = ~n2050 & n4307;
  assign n4309 = ~n2049 & n4308;
  assign n4310 = ~n1351 & n4309;
  assign n4311 = ~n1349 & n4310;
  assign n4312 = ~n3158 & n4311;
  assign n4313 = ~n1338 & n4312;
  assign n4314 = ~n2047 & n4313;
  assign n4315 = ~n1334 & n4314;
  assign n4316 = ~n1326 & n4315;
  assign n4317 = ~n2044 & n4316;
  assign n4318 = ~n1323 & n4317;
  assign n4319 = ~n1320 & n4318;
  assign n4320 = ~n1316 & n4319;
  assign n4321 = ~n2040 & n4320;
  assign n4322 = ~n3156 & n4321;
  assign n4323 = ~n1309 & n4322;
  assign n4324 = ~n2039 & n4323;
  assign n4325 = ~n1303 & n4324;
  assign n4326 = ~n3155 & n4325;
  assign n4327 = ~n2038 & n4326;
  assign n4328 = ~n1298 & n4327;
  assign n4329 = ~n1291 & n4328;
  assign n4330 = ~n1271 & n3160;
  assign n4331 = n4329 & ~n4330;
  assign n4332 = ~n4302 & n4331;
  assign n4333 = ~n4301 & n4332;
  assign n4334 = ~n4300 & n4333;
  assign n4335 = \data<6>  & n504;
  assign n4336 = n4334 & n4335;
  assign n4337 = ~\data<6>  & n504;
  assign n4338 = ~n4334 & n4337;
  assign n4339 = \outreg<9>  & n508;
  assign n4340 = \outreg<17>  & n510;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = ~n4338 & n4341;
  assign \outreg_new<9>  = n4336 | ~n4342;
  assign n4344 = ~n2104 & n3598;
  assign n4345 = n2104 & n2132;
  assign n4346 = ~n2104 & n3606;
  assign n4347 = n2104 & n2180;
  assign n4348 = n2104 & n2169;
  assign n4349 = n2104 & n2126;
  assign n4350 = ~n2193 & ~n2196;
  assign n4351 = ~n4347 & n4350;
  assign n4352 = ~n2191 & n4351;
  assign n4353 = ~n3607 & n4352;
  assign n4354 = ~n3604 & n4353;
  assign n4355 = ~n2186 & n4354;
  assign n4356 = ~n3602 & n4355;
  assign n4357 = ~n2177 & n4356;
  assign n4358 = ~n2175 & n4357;
  assign n4359 = ~n4346 & n4358;
  assign n4360 = ~n2170 & n4359;
  assign n4361 = ~n3601 & n4360;
  assign n4362 = ~n2163 & n4361;
  assign n4363 = ~n3599 & n4362;
  assign n4364 = ~n2158 & n4363;
  assign n4365 = ~n3595 & n4364;
  assign n4366 = ~n2154 & n4365;
  assign n4367 = ~n2151 & n4366;
  assign n4368 = ~n4345 & n4367;
  assign n4369 = ~n2148 & n4368;
  assign n4370 = ~n4344 & n4369;
  assign n4371 = ~n2145 & n4370;
  assign n4372 = ~n2142 & n4371;
  assign n4373 = ~n3593 & n4372;
  assign n4374 = ~n3591 & n4373;
  assign n4375 = ~n2127 & n4374;
  assign n4376 = ~n2124 & n4375;
  assign n4377 = ~n2104 & n3612;
  assign n4378 = n4376 & ~n4377;
  assign n4379 = ~n2104 & n3610;
  assign n4380 = n4378 & ~n4379;
  assign n4381 = ~n4349 & n4380;
  assign n4382 = ~n4348 & n4381;
  assign n4383 = \data<9>  & n504;
  assign n4384 = n4382 & n4383;
  assign n4385 = ~\data<9>  & n504;
  assign n4386 = ~n4382 & n4385;
  assign n4387 = \outreg<59>  & n510;
  assign n4388 = \outreg<51>  & n508;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390 = ~n4386 & n4389;
  assign \outreg_new<51>  = n4384 | ~n4390;
  assign n4392 = \outreg<60>  & n510;
  assign n4393 = \outreg<52>  & n508;
  assign n4394 = \data<49>  & n504;
  assign n4395 = ~n4393 & ~n4394;
  assign \outreg_new<52>  = n4392 | ~n4395;
  assign n4397 = n1607 & n1666;
  assign n4398 = ~n1607 & n1704;
  assign n4399 = ~n1607 & n1640;
  assign n4400 = ~n1701 & ~n1703;
  assign n4401 = ~n1989 & n4400;
  assign n4402 = ~n1696 & n4401;
  assign n4403 = ~n2372 & n4402;
  assign n4404 = ~n1692 & n4403;
  assign n4405 = ~n1689 & n4404;
  assign n4406 = ~n2371 & n4405;
  assign n4407 = ~n1685 & n4406;
  assign n4408 = ~n1682 & n4407;
  assign n4409 = ~n1986 & n4408;
  assign n4410 = ~n1985 & n4409;
  assign n4411 = ~n1674 & n4410;
  assign n4412 = ~n1670 & n4411;
  assign n4413 = ~n1665 & n4412;
  assign n4414 = ~n2370 & n4413;
  assign n4415 = ~n1662 & n4414;
  assign n4416 = ~n1982 & n4415;
  assign n4417 = ~n1660 & n4416;
  assign n4418 = ~n1981 & n4417;
  assign n4419 = ~n2369 & n4418;
  assign n4420 = ~n1649 & n4419;
  assign n4421 = ~n1980 & n4420;
  assign n4422 = ~n1647 & n4421;
  assign n4423 = ~n1637 & n4422;
  assign n4424 = ~n1632 & n4423;
  assign n4425 = ~n1978 & n4424;
  assign n4426 = ~n1977 & n4425;
  assign n4427 = ~n1607 & n1990;
  assign n4428 = n4426 & ~n4427;
  assign n4429 = ~n4399 & n4428;
  assign n4430 = ~n4398 & n4429;
  assign n4431 = ~n4397 & n4430;
  assign n4432 = \data<17>  & n504;
  assign n4433 = n4431 & n4432;
  assign n4434 = ~\data<17>  & n504;
  assign n4435 = ~n4431 & n4434;
  assign n4436 = \outreg<61>  & n510;
  assign n4437 = \outreg<53>  & n508;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = ~n4435 & n4438;
  assign \outreg_new<53>  = n4433 | ~n4439;
  assign n4441 = \data<23>  & n504;
  assign n4442 = n3699 & n4441;
  assign n4443 = ~\data<23>  & n504;
  assign n4444 = ~n3699 & n4443;
  assign n4445 = \outreg<5>  & n508;
  assign n4446 = \outreg<13>  & n510;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = ~n4444 & n4447;
  assign \outreg_new<5>  = n4442 | ~n4448;
  assign n4450 = \outreg<62>  & n510;
  assign n4451 = \outreg<54>  & n508;
  assign n4452 = \data<57>  & n504;
  assign n4453 = ~n4451 & ~n4452;
  assign \outreg_new<54>  = n4450 | ~n4453;
  assign n4455 = \outreg<6>  & n508;
  assign n4456 = \outreg<14>  & n510;
  assign n4457 = \data<63>  & n504;
  assign n4458 = ~n4456 & ~n4457;
  assign \outreg_new<6>  = n4455 | ~n4458;
  assign n4460 = \data<31>  & n504;
  assign n4461 = n3193 & n4460;
  assign n4462 = ~\data<31>  & n504;
  assign n4463 = ~n3193 & n4462;
  assign n4464 = \outreg<7>  & n508;
  assign n4465 = \outreg<15>  & n510;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~n4463 & n4466;
  assign \outreg_new<7>  = n4461 | ~n4467;
  assign n4469 = \outreg<8>  & n508;
  assign n4470 = \outreg<16>  & n510;
  assign n4471 = \data<38>  & n504;
  assign n4472 = ~n4470 & ~n4471;
  assign \outreg_new<8>  = n4469 | ~n4472;
  assign n4474 = n880 & n945;
  assign n4475 = n880 & n910;
  assign n4476 = ~n880 & n962;
  assign n4477 = ~n976 & ~n3710;
  assign n4478 = ~n2260 & n4477;
  assign n4479 = ~n968 & n4478;
  assign n4480 = ~n966 & n4479;
  assign n4481 = ~n963 & n4480;
  assign n4482 = ~n2258 & n4481;
  assign n4483 = ~n961 & n4482;
  assign n4484 = ~n2257 & n4483;
  assign n4485 = ~n958 & n4484;
  assign n4486 = ~n951 & n4485;
  assign n4487 = ~n943 & n4486;
  assign n4488 = ~n3709 & n4487;
  assign n4489 = ~n2255 & n4488;
  assign n4490 = ~n2253 & n4489;
  assign n4491 = ~n3708 & n4490;
  assign n4492 = ~n934 & n4491;
  assign n4493 = ~n931 & n4492;
  assign n4494 = ~n2252 & n4493;
  assign n4495 = ~n930 & n4494;
  assign n4496 = ~n922 & n4495;
  assign n4497 = ~n2250 & n4496;
  assign n4498 = ~n920 & n4497;
  assign n4499 = ~n914 & n4498;
  assign n4500 = ~n911 & n4499;
  assign n4501 = ~n904 & n4500;
  assign n4502 = ~n2249 & n4501;
  assign n4503 = ~n3707 & n4502;
  assign n4504 = ~n880 & n3712;
  assign n4505 = n4503 & ~n4504;
  assign n4506 = ~n4476 & n4505;
  assign n4507 = ~n4475 & n4506;
  assign n4508 = ~n4474 & n4507;
  assign n4509 = \data<7>  & n504;
  assign n4510 = n4508 & n4509;
  assign n4511 = ~\data<7>  & n504;
  assign n4512 = ~n4508 & n4511;
  assign n4513 = \outreg<9>  & n510;
  assign n4514 = \outreg<1>  & n508;
  assign n4515 = ~n4513 & ~n4514;
  assign n4516 = ~n4512 & n4515;
  assign \outreg_new<1>  = n4510 | ~n4516;
  assign n4518 = \outreg<58>  & n510;
  assign n4519 = \outreg<50>  & n508;
  assign n4520 = \data<41>  & n504;
  assign n4521 = ~n4519 & ~n4520;
  assign \outreg_new<50>  = n4518 | ~n4521;
  assign n4523 = \outreg<2>  & n508;
  assign n4524 = \outreg<10>  & n510;
  assign n4525 = \data<47>  & n504;
  assign n4526 = ~n4524 & ~n4525;
  assign \outreg_new<2>  = n4523 | ~n4526;
  assign n4528 = ~n687 & n1063;
  assign n4529 = n687 & n733;
  assign n4530 = ~n687 & n777;
  assign n4531 = n687 & n762;
  assign n4532 = n687 & n812;
  assign n4533 = n687 & n1068;
  assign n4534 = ~n687 & n755;
  assign n4535 = ~n780 & ~n4531;
  assign n4536 = ~n1061 & n4535;
  assign n4537 = ~n774 & n4536;
  assign n4538 = ~n767 & n4537;
  assign n4539 = ~n1060 & n4538;
  assign n4540 = ~n765 & n4539;
  assign n4541 = ~n4530 & n4540;
  assign n4542 = ~n763 & n4541;
  assign n4543 = ~n1059 & n4542;
  assign n4544 = ~n1054 & n4543;
  assign n4545 = ~n756 & n4544;
  assign n4546 = ~n1053 & n4545;
  assign n4547 = ~n750 & n4546;
  assign n4548 = ~n749 & n4547;
  assign n4549 = ~n4529 & n4548;
  assign n4550 = ~n1051 & n4549;
  assign n4551 = ~n745 & n4550;
  assign n4552 = ~n743 & n4551;
  assign n4553 = ~n4528 & n4552;
  assign n4554 = ~n1049 & n4553;
  assign n4555 = ~n734 & n4554;
  assign n4556 = ~n729 & n4555;
  assign n4557 = ~n725 & n4556;
  assign n4558 = ~n722 & n4557;
  assign n4559 = ~n1047 & n4558;
  assign n4560 = ~n714 & n4559;
  assign n4561 = ~n707 & n4560;
  assign n4562 = ~n687 & n775;
  assign n4563 = n4561 & ~n4562;
  assign n4564 = ~n4534 & n4563;
  assign n4565 = ~n4533 & n4564;
  assign n4566 = ~n4532 & n4565;
  assign n4567 = \data<8>  & n504;
  assign n4568 = n4566 & n4567;
  assign n4569 = ~\data<8>  & n504;
  assign n4570 = ~n4566 & n4569;
  assign n4571 = \outreg<59>  & n508;
  assign n4572 = ~n4570 & ~n4571;
  assign \outreg_new<59>  = n4568 | ~n4572;
  assign n4574 = n1117 & n1157;
  assign n4575 = n1117 & n1179;
  assign n4576 = ~n1117 & n1163;
  assign n4577 = ~n1117 & n1211;
  assign n4578 = ~n1431 & ~n1432;
  assign n4579 = ~n1210 & n4578;
  assign n4580 = ~n1208 & n4579;
  assign n4581 = ~n1205 & n4580;
  assign n4582 = ~n3664 & n4581;
  assign n4583 = ~n1202 & n4582;
  assign n4584 = ~n1198 & n4583;
  assign n4585 = ~n1196 & n4584;
  assign n4586 = ~n1430 & n4585;
  assign n4587 = ~n1184 & n4586;
  assign n4588 = ~n1428 & n4587;
  assign n4589 = ~n3663 & n4588;
  assign n4590 = ~n1177 & n4589;
  assign n4591 = ~n1172 & n4590;
  assign n4592 = ~n1427 & n4591;
  assign n4593 = ~n1167 & n4592;
  assign n4594 = ~n3662 & n4593;
  assign n4595 = ~n1162 & n4594;
  assign n4596 = ~n1425 & n4595;
  assign n4597 = ~n1161 & n4596;
  assign n4598 = ~n1158 & n4597;
  assign n4599 = ~n1421 & n4598;
  assign n4600 = ~n1151 & n4599;
  assign n4601 = ~n1146 & n4600;
  assign n4602 = ~n1419 & n4601;
  assign n4603 = ~n1137 & n4602;
  assign n4604 = ~n3661 & n4603;
  assign n4605 = ~n4577 & n4604;
  assign n4606 = ~n4576 & n4605;
  assign n4607 = ~n4575 & n4606;
  assign n4608 = ~n4574 & n4607;
  assign n4609 = \data<15>  & n504;
  assign n4610 = n4608 & n4609;
  assign n4611 = ~\data<15>  & n504;
  assign n4612 = ~n4608 & n4611;
  assign n4613 = \outreg<3>  & n508;
  assign n4614 = \outreg<11>  & n510;
  assign n4615 = ~n4613 & ~n4614;
  assign n4616 = ~n4612 & n4615;
  assign \outreg_new<3>  = n4610 | ~n4616;
  assign n4618 = \outreg<4>  & n508;
  assign n4619 = \outreg<12>  & n510;
  assign n4620 = \data<55>  & n504;
  assign n4621 = ~n4619 & ~n4620;
  assign \outreg_new<4>  = n4618 | ~n4621;
  assign n4623 = \data<25>  & n504;
  assign n4624 = n3646 & n4623;
  assign n4625 = ~\data<25>  & n504;
  assign n4626 = ~n3646 & n4625;
  assign n4627 = \outreg<63>  & n510;
  assign n4628 = \outreg<55>  & n508;
  assign n4629 = ~n4627 & ~n4628;
  assign n4630 = ~n4626 & n4629;
  assign \outreg_new<55>  = n4624 | ~n4630;
  assign n4632 = \data<11>  & ~n504;
  assign n4633 = n2087 & n4632;
  assign n4634 = ~\data<11>  & ~n504;
  assign n4635 = ~n2087 & n4634;
  assign n4636 = \inreg<26>  & n504;
  assign n4637 = ~n4635 & ~n4636;
  assign \data_new<43>  = n4633 | ~n4637;
  assign n4639 = \outreg<56>  & n508;
  assign n4640 = \data<32>  & n504;
  assign \outreg_new<56>  = n4639 | n4640;
  assign n4642 = \data<12>  & ~n504;
  assign n4643 = n1740 & n4642;
  assign n4644 = ~\data<12>  & ~n504;
  assign n4645 = ~n1740 & n4644;
  assign n4646 = \inreg<18>  & n504;
  assign n4647 = ~n4645 & ~n4646;
  assign \data_new<44>  = n4643 | ~n4647;
  assign n4649 = \outreg<8>  & n510;
  assign n4650 = \outreg<0>  & n508;
  assign n4651 = \data<39>  & n504;
  assign n4652 = ~n4650 & ~n4651;
  assign \outreg_new<0>  = n4649 | ~n4652;
  assign n4654 = n2104 & n2199;
  assign n4655 = n2104 & n2228;
  assign n4656 = ~n2104 & n3603;
  assign n4657 = n2201 & ~n4347;
  assign n4658 = ~n3609 & n4657;
  assign n4659 = ~n2190 & n4658;
  assign n4660 = ~n3604 & n4659;
  assign n4661 = ~n2186 & n4660;
  assign n4662 = ~n2184 & n4661;
  assign n4663 = ~n3602 & n4662;
  assign n4664 = ~n2181 & n4663;
  assign n4665 = ~n2175 & n4664;
  assign n4666 = ~n4346 & n4665;
  assign n4667 = ~n2170 & n4666;
  assign n4668 = ~n3600 & n4667;
  assign n4669 = ~n3597 & n4668;
  assign n4670 = ~n3595 & n4669;
  assign n4671 = ~n2154 & n4670;
  assign n4672 = ~n2153 & n4671;
  assign n4673 = ~n2151 & n4672;
  assign n4674 = ~n4345 & n4673;
  assign n4675 = ~n2146 & n4674;
  assign n4676 = ~n4344 & n4675;
  assign n4677 = ~n2145 & n4676;
  assign n4678 = ~n2138 & n4677;
  assign n4679 = ~n3592 & n4678;
  assign n4680 = ~n2133 & n4679;
  assign n4681 = ~n3591 & n4680;
  assign n4682 = ~n2127 & n4681;
  assign n4683 = ~n2104 & n3594;
  assign n4684 = n4682 & ~n4683;
  assign n4685 = ~n4656 & n4684;
  assign n4686 = ~n4655 & n4685;
  assign n4687 = ~n4654 & n4686;
  assign n4688 = \data<0>  & n504;
  assign n4689 = n4687 & n4688;
  assign n4690 = ~\data<0>  & n504;
  assign n4691 = ~n4687 & n4690;
  assign n4692 = \outreg<57>  & n508;
  assign n4693 = ~n4691 & ~n4692;
  assign \outreg_new<57>  = n4689 | ~n4693;
  assign n4695 = \data<9>  & ~n504;
  assign n4696 = n4382 & n4695;
  assign n4697 = ~\data<9>  & ~n504;
  assign n4698 = ~n4382 & n4697;
  assign n4699 = \inreg<42>  & n504;
  assign n4700 = ~n4698 & ~n4699;
  assign \data_new<41>  = n4696 | ~n4700;
  assign n4702 = \outreg<58>  & n508;
  assign n4703 = \data<40>  & n504;
  assign \outreg_new<58>  = n4702 | n4703;
  assign n4705 = \data<10>  & ~n504;
  assign n4706 = n2349 & n4705;
  assign n4707 = ~\data<10>  & ~n504;
  assign n4708 = ~n2349 & n4707;
  assign n4709 = \inreg<34>  & n504;
  assign n4710 = ~n4708 & ~n4709;
  assign \data_new<42>  = n4706 | ~n4710;
  assign n4712 = \inreg<20>  & n508;
  assign n4713 = \inreg<12>  & n510;
  assign \inreg_new<20>  = n4712 | n4713;
  assign n4715 = n687 & n742;
  assign n4716 = n687 & n773;
  assign n4717 = ~n687 & n1065;
  assign n4718 = n785 & ~n4531;
  assign n4719 = ~n1062 & n4718;
  assign n4720 = ~n776 & n4719;
  assign n4721 = ~n774 & n4720;
  assign n4722 = ~n771 & n4721;
  assign n4723 = ~n767 & n4722;
  assign n4724 = ~n1060 & n4723;
  assign n4725 = ~n764 & n4724;
  assign n4726 = ~n4530 & n4725;
  assign n4727 = ~n1057 & n4726;
  assign n4728 = ~n1054 & n4727;
  assign n4729 = ~n756 & n4728;
  assign n4730 = ~n1053 & n4729;
  assign n4731 = ~n753 & n4730;
  assign n4732 = ~n749 & n4731;
  assign n4733 = ~n4529 & n4732;
  assign n4734 = ~n747 & n4733;
  assign n4735 = ~n1050 & n4734;
  assign n4736 = ~n743 & n4735;
  assign n4737 = ~n4528 & n4736;
  assign n4738 = ~n739 & n4737;
  assign n4739 = ~n1048 & n4738;
  assign n4740 = ~n729 & n4739;
  assign n4741 = ~n725 & n4740;
  assign n4742 = ~n719 & n4741;
  assign n4743 = ~n1047 & n4742;
  assign n4744 = ~n4717 & n4743;
  assign n4745 = ~n687 & n1052;
  assign n4746 = n4744 & ~n4745;
  assign n4747 = ~n4716 & n4746;
  assign n4748 = ~n4715 & n4747;
  assign n4749 = \data<16>  & n504;
  assign n4750 = n4748 & n4749;
  assign n4751 = ~\data<16>  & n504;
  assign n4752 = ~n4748 & n4751;
  assign n4753 = \outreg<61>  & n508;
  assign n4754 = ~n4752 & ~n4753;
  assign \outreg_new<61>  = n4750 | ~n4754;
  assign n4756 = \outreg<62>  & n508;
  assign n4757 = \data<56>  & n504;
  assign \outreg_new<62>  = n4756 | n4757;
  assign n4759 = \data<8>  & ~n504;
  assign n4760 = n4566 & n4759;
  assign n4761 = ~\data<8>  & ~n504;
  assign n4762 = ~n4566 & n4761;
  assign n4763 = \inreg<50>  & n504;
  assign n4764 = ~n4762 & ~n4763;
  assign \data_new<40>  = n4760 | ~n4764;
  assign n4766 = \data<24>  & n504;
  assign n4767 = n3746 & n4766;
  assign n4768 = ~\data<24>  & n504;
  assign n4769 = ~n3746 & n4768;
  assign n4770 = \outreg<63>  & n508;
  assign n4771 = ~n4769 & ~n4770;
  assign \outreg_new<63>  = n4767 | ~n4771;
  assign n4773 = \inreg<24>  & n508;
  assign n4774 = \inreg<16>  & n510;
  assign \inreg_new<24>  = n4773 | n4774;
  assign n4776 = \inreg<23>  & n508;
  assign n4777 = \inreg<15>  & n510;
  assign \inreg_new<23>  = n4776 | n4777;
  assign n4779 = \inreg<22>  & n508;
  assign n4780 = \inreg<14>  & n510;
  assign \inreg_new<22>  = n4779 | n4780;
  assign n4782 = \data<17>  & ~n504;
  assign n4783 = n4431 & n4782;
  assign n4784 = ~\data<17>  & ~n504;
  assign n4785 = ~n4431 & n4784;
  assign n4786 = \inreg<44>  & n504;
  assign n4787 = ~n4785 & ~n4786;
  assign \data_new<49>  = n4783 | ~n4787;
  assign n4789 = \inreg<21>  & n508;
  assign n4790 = \inreg<13>  & n510;
  assign \inreg_new<21>  = n4789 | n4790;
  assign n4792 = \outreg<60>  & n508;
  assign n4793 = \data<48>  & n504;
  assign \outreg_new<60>  = n4792 | n4793;
  assign n4795 = \inreg<28>  & n508;
  assign n4796 = \inreg<20>  & n510;
  assign \inreg_new<28>  = n4795 | n4796;
  assign n4798 = \data<15>  & ~n504;
  assign n4799 = n4608 & n4798;
  assign n4800 = ~\data<15>  & ~n504;
  assign n4801 = ~n4608 & n4800;
  assign n4802 = \data_in<2>  & n504;
  assign n4803 = ~n4801 & ~n4802;
  assign \data_new<47>  = n4799 | ~n4803;
  assign n4805 = \inreg<27>  & n508;
  assign n4806 = \inreg<19>  & n510;
  assign \inreg_new<27>  = n4805 | n4806;
  assign n4808 = \data<16>  & ~n504;
  assign n4809 = n4748 & n4808;
  assign n4810 = ~\data<16>  & ~n504;
  assign n4811 = ~n4748 & n4810;
  assign n4812 = \inreg<52>  & n504;
  assign n4813 = ~n4811 & ~n4812;
  assign \data_new<48>  = n4809 | ~n4813;
  assign n4815 = \inreg<26>  & n508;
  assign n4816 = \inreg<18>  & n510;
  assign \inreg_new<26>  = n4815 | n4816;
  assign n4818 = \data<13>  & ~n504;
  assign n4819 = n1015 & n4818;
  assign n4820 = ~\data<13>  & ~n504;
  assign n4821 = ~n1015 & n4820;
  assign n4822 = \inreg<10>  & n504;
  assign n4823 = ~n4821 & ~n4822;
  assign \data_new<45>  = n4819 | ~n4823;
  assign n4825 = \inreg<25>  & n508;
  assign n4826 = \inreg<17>  & n510;
  assign \inreg_new<25>  = n4825 | n4826;
  assign n4828 = \data<14>  & ~n504;
  assign n4829 = n664 & n4828;
  assign n4830 = ~\data<14>  & ~n504;
  assign n4831 = ~n664 & n4830;
  assign n4832 = \inreg<2>  & n504;
  assign n4833 = ~n4831 & ~n4832;
  assign \data_new<46>  = n4829 | ~n4833;
  assign n4835 = \data<1>  & ~n504;
  assign n4836 = n2406 & n4835;
  assign n4837 = ~\data<1>  & ~n504;
  assign n4838 = ~n2406 & n4837;
  assign n4839 = \inreg<40>  & n504;
  assign n4840 = ~n4838 & ~n4839;
  assign \data_new<33>  = n4836 | ~n4840;
  assign n4842 = \data<2>  & ~n504;
  assign n4843 = n2296 & n4842;
  assign n4844 = ~\data<2>  & ~n504;
  assign n4845 = ~n2296 & n4844;
  assign n4846 = \inreg<32>  & n504;
  assign n4847 = ~n4845 & ~n4846;
  assign \data_new<34>  = n4843 | ~n4847;
  assign n4849 = \data<63>  & ~n504;
  assign n4850 = \data_in<7>  & n504;
  assign \data_new<31>  = n4849 | n4850;
  assign n4852 = \inreg<29>  & n508;
  assign n4853 = \inreg<21>  & n510;
  assign \inreg_new<29>  = n4852 | n4853;
  assign n4855 = \data<0>  & ~n504;
  assign n4856 = n4687 & n4855;
  assign n4857 = ~\data<0>  & ~n504;
  assign n4858 = ~n4687 & n4857;
  assign n4859 = \inreg<48>  & n504;
  assign n4860 = ~n4858 & ~n4859;
  assign \data_new<32>  = n4856 | ~n4860;
  assign n4862 = \inreg<2>  & n510;
  assign n4863 = \inreg<10>  & n508;
  assign \inreg_new<10>  = n4862 | n4863;
  assign n4865 = \data<62>  & ~n504;
  assign n4866 = \inreg<7>  & n504;
  assign \data_new<30>  = n4865 | n4866;
  assign n4868 = \inreg<6>  & n510;
  assign n4869 = \inreg<14>  & n508;
  assign \inreg_new<14>  = n4868 | n4869;
  assign n4871 = \inreg<5>  & n510;
  assign n4872 = \inreg<13>  & n508;
  assign \inreg_new<13>  = n4871 | n4872;
  assign n4874 = \inreg<4>  & n510;
  assign n4875 = \inreg<12>  & n508;
  assign \inreg_new<12>  = n4874 | n4875;
  assign n4877 = \data<7>  & ~n504;
  assign n4878 = n4508 & n4877;
  assign n4879 = ~\data<7>  & ~n504;
  assign n4880 = ~n4508 & n4879;
  assign n4881 = \data_in<0>  & n504;
  assign n4882 = ~n4880 & ~n4881;
  assign \data_new<39>  = n4878 | ~n4882;
  assign n4884 = \inreg<3>  & n510;
  assign n4885 = \inreg<11>  & n508;
  assign \inreg_new<11>  = n4884 | n4885;
  assign n4887 = \inreg<18>  & n508;
  assign n4888 = \inreg<10>  & n510;
  assign \inreg_new<18>  = n4887 | n4888;
  assign n4890 = \data<5>  & ~n504;
  assign n4891 = n1251 & n4890;
  assign n4892 = ~\data<5>  & ~n504;
  assign n4893 = ~n1251 & n4892;
  assign n4894 = \inreg<8>  & n504;
  assign n4895 = ~n4893 & ~n4894;
  assign \data_new<37>  = n4891 | ~n4895;
  assign n4897 = \inreg<9>  & n510;
  assign n4898 = \inreg<17>  & n508;
  assign \inreg_new<17>  = n4897 | n4898;
  assign n4900 = \data<6>  & ~n504;
  assign n4901 = n4334 & n4900;
  assign n4902 = ~\data<6>  & ~n504;
  assign n4903 = ~n4334 & n4902;
  assign n4904 = \inreg<0>  & n504;
  assign n4905 = ~n4903 & ~n4904;
  assign \data_new<38>  = n4901 | ~n4905;
  assign n4907 = \inreg<8>  & n510;
  assign n4908 = \inreg<16>  & n508;
  assign \inreg_new<16>  = n4907 | n4908;
  assign n4910 = \data<3>  & ~n504;
  assign n4911 = n1956 & n4910;
  assign n4912 = ~\data<3>  & ~n504;
  assign n4913 = ~n1956 & n4912;
  assign n4914 = \inreg<24>  & n504;
  assign n4915 = ~n4913 & ~n4914;
  assign \data_new<35>  = n4911 | ~n4915;
  assign n4917 = \inreg<7>  & n510;
  assign n4918 = \inreg<15>  & n508;
  assign \inreg_new<15>  = n4917 | n4918;
  assign n4920 = \data<4>  & ~n504;
  assign n4921 = n1590 & n4920;
  assign n4922 = ~\data<4>  & ~n504;
  assign n4923 = ~n1590 & n4922;
  assign n4924 = \inreg<16>  & n504;
  assign n4925 = ~n4923 & ~n4924;
  assign \data_new<36>  = n4921 | ~n4925;
  assign n4927 = \data<55>  & ~n504;
  assign n4928 = \data_in<5>  & n504;
  assign \data_new<23>  = n4927 | n4928;
  assign n4930 = \data<56>  & ~n504;
  assign n4931 = \inreg<55>  & n504;
  assign \data_new<24>  = n4930 | n4931;
  assign n4933 = \data<53>  & ~n504;
  assign n4934 = \inreg<13>  & n504;
  assign \data_new<21>  = n4933 | n4934;
  assign n4936 = \inreg<19>  & n508;
  assign n4937 = \inreg<11>  & n510;
  assign \inreg_new<19>  = n4936 | n4937;
  assign n4939 = \data<54>  & ~n504;
  assign n4940 = \inreg<5>  & n504;
  assign \data_new<22>  = n4939 | n4940;
  assign n4942 = \inreg<40>  & n508;
  assign n4943 = \inreg<32>  & n510;
  assign \inreg_new<40>  = n4942 | n4943;
  assign n4945 = \data<52>  & ~n504;
  assign n4946 = \inreg<21>  & n504;
  assign \data_new<20>  = n4945 | n4946;
  assign n4948 = \inreg<44>  & n508;
  assign n4949 = \inreg<36>  & n510;
  assign \inreg_new<44>  = n4948 | n4949;
  assign n4951 = \inreg<43>  & n508;
  assign n4952 = \inreg<35>  & n510;
  assign \inreg_new<43>  = n4951 | n4952;
  assign n4954 = \inreg<42>  & n508;
  assign n4955 = \inreg<34>  & n510;
  assign \inreg_new<42>  = n4954 | n4955;
  assign n4957 = \data<61>  & ~n504;
  assign n4958 = \inreg<15>  & n504;
  assign \data_new<29>  = n4957 | n4958;
  assign n4960 = \inreg<41>  & n508;
  assign n4961 = \inreg<33>  & n510;
  assign \inreg_new<41>  = n4960 | n4961;
  assign n4963 = \inreg<48>  & n508;
  assign n4964 = \inreg<40>  & n510;
  assign \inreg_new<48>  = n4963 | n4964;
  assign n4966 = \data<59>  & ~n504;
  assign n4967 = \inreg<31>  & n504;
  assign \data_new<27>  = n4966 | n4967;
  assign n4969 = \inreg<47>  & n508;
  assign n4970 = \inreg<39>  & n510;
  assign \inreg_new<47>  = n4969 | n4970;
  assign n4972 = \data<60>  & ~n504;
  assign n4973 = \inreg<23>  & n504;
  assign \data_new<28>  = n4972 | n4973;
  assign n4975 = \inreg<46>  & n508;
  assign n4976 = \inreg<38>  & n510;
  assign \inreg_new<46>  = n4975 | n4976;
endmodule


