// Benchmark "vda" written by ABC on Tue May 16 16:07:53 2017

module vda ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q,
    r, s, t, u, v, w, x, y, z, a0, a1, b0, b1, c0, c1, d0, d1, e0, f0, g0,
    h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0,
    z0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q;
  output r, s, t, u, v, w, x, y, z, a0, a1, b0, b1, c0, c1, d0, d1, e0, f0,
    g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0,
    y0, z0;
  wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n411, n412, n415, n416, n418, n419, n420, n421,
    n422, n423, n425, n426, n427, n428, n429, n431, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n794, n795, n796, n797, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1080, n1081, n1082, n1083, n1084, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112;
  assign n57 = l & m;
  assign n58 = ~n & n57;
  assign n59 = o & n58;
  assign n60 = ~p & n59;
  assign n61 = ~q & n60;
  assign n62 = ~o & n58;
  assign n63 = p & n62;
  assign n64 = q & n63;
  assign n65 = ~g & ~l;
  assign n66 = m & n65;
  assign n67 = ~n & n66;
  assign n68 = o & n67;
  assign n69 = p & n68;
  assign n70 = ~q & n69;
  assign n71 = n & n57;
  assign n72 = ~o & n71;
  assign n73 = ~p & n72;
  assign n74 = ~q & n73;
  assign n75 = l & ~m;
  assign n76 = ~n & n75;
  assign n77 = o & n76;
  assign n78 = ~p & n77;
  assign n79 = q & n78;
  assign n80 = p & n72;
  assign n81 = q & n80;
  assign n82 = n & n66;
  assign n83 = ~o & n82;
  assign n84 = p & n83;
  assign n85 = q & n84;
  assign n86 = ~l & ~m;
  assign n87 = n & n86;
  assign n88 = o & n87;
  assign n89 = ~p & n88;
  assign n90 = q & n89;
  assign n91 = ~l & m;
  assign n92 = ~n & n91;
  assign n93 = o & n92;
  assign n94 = p & n93;
  assign n95 = q & n94;
  assign n96 = p & n77;
  assign n97 = ~q & n96;
  assign n98 = ~o & n92;
  assign n99 = ~p & n98;
  assign n100 = ~q & n99;
  assign n101 = i & ~l;
  assign n102 = ~m & n101;
  assign n103 = n & n102;
  assign n104 = ~o & n103;
  assign n105 = p & n104;
  assign n106 = q & n105;
  assign n107 = ~q & n89;
  assign n108 = ~n & n86;
  assign n109 = o & n108;
  assign n110 = ~p & n109;
  assign n111 = ~q & n110;
  assign n112 = p & n109;
  assign n113 = ~q & n112;
  assign n114 = ~g & l;
  assign n115 = ~m & n114;
  assign n116 = ~n & n115;
  assign n117 = o & n116;
  assign n118 = p & n117;
  assign n119 = q & n118;
  assign n120 = g & ~l;
  assign n121 = ~m & n120;
  assign n122 = n & n121;
  assign n123 = o & n122;
  assign n124 = p & n123;
  assign n125 = q & n124;
  assign n126 = ~b & f;
  assign n127 = ~l & n126;
  assign n128 = ~m & n127;
  assign n129 = ~n & n128;
  assign n130 = ~o & n129;
  assign n131 = p & n130;
  assign n132 = q & n131;
  assign n133 = ~o & n76;
  assign n134 = p & n133;
  assign n135 = ~q & n134;
  assign n136 = m & n120;
  assign n137 = ~n & n136;
  assign n138 = o & n137;
  assign n139 = ~p & n138;
  assign n140 = ~q & n139;
  assign n141 = ~o & n87;
  assign n142 = ~p & n141;
  assign n143 = ~q & n142;
  assign n144 = ~o & n108;
  assign n145 = p & n144;
  assign n146 = ~q & n145;
  assign n147 = q & n110;
  assign n148 = ~f & ~l;
  assign n149 = ~m & n148;
  assign n150 = n & n149;
  assign n151 = ~o & n150;
  assign n152 = p & n151;
  assign n153 = ~q & n152;
  assign n154 = g & l;
  assign n155 = ~m & n154;
  assign n156 = ~n & n155;
  assign n157 = o & n156;
  assign n158 = p & n157;
  assign n159 = q & n158;
  assign n160 = f & ~l;
  assign n161 = ~m & n160;
  assign n162 = n & n161;
  assign n163 = ~o & n162;
  assign n164 = p & n163;
  assign n165 = ~q & n164;
  assign n166 = c & ~l;
  assign n167 = ~m & n166;
  assign n168 = ~n & n167;
  assign n169 = ~o & n168;
  assign n170 = ~p & n169;
  assign n171 = q & n170;
  assign n172 = e & ~f;
  assign n173 = ~l & n172;
  assign n174 = ~m & n173;
  assign n175 = ~n & n174;
  assign n176 = ~o & n175;
  assign n177 = p & n176;
  assign n178 = q & n177;
  assign n179 = b & e;
  assign n180 = ~l & n179;
  assign n181 = ~m & n180;
  assign n182 = ~n & n181;
  assign n183 = ~o & n182;
  assign n184 = p & n183;
  assign n185 = q & n184;
  assign n186 = a & e;
  assign n187 = l & n186;
  assign n188 = ~m & n187;
  assign n189 = ~n & n188;
  assign n190 = o & n189;
  assign n191 = ~p & n190;
  assign n192 = ~q & n191;
  assign n193 = h & n172;
  assign n194 = ~i & n193;
  assign n195 = j & n194;
  assign n196 = ~l & n195;
  assign n197 = m & n196;
  assign n198 = n & n197;
  assign n199 = o & n198;
  assign n200 = p & n199;
  assign n201 = ~q & n200;
  assign n202 = ~c & e;
  assign n203 = h & n202;
  assign n204 = ~i & n203;
  assign n205 = j & n204;
  assign n206 = ~l & n205;
  assign n207 = m & n206;
  assign n208 = n & n207;
  assign n209 = o & n208;
  assign n210 = p & n209;
  assign n211 = ~q & n210;
  assign n212 = h & n179;
  assign n213 = ~i & n212;
  assign n214 = j & n213;
  assign n215 = ~l & n214;
  assign n216 = m & n215;
  assign n217 = n & n216;
  assign n218 = o & n217;
  assign n219 = p & n218;
  assign n220 = ~q & n219;
  assign n221 = ~n211 & ~n220;
  assign n222 = ~n201 & n221;
  assign n223 = ~n192 & n222;
  assign n224 = ~n185 & n223;
  assign n225 = ~n178 & n224;
  assign n226 = ~n171 & n225;
  assign n227 = ~n165 & n226;
  assign n228 = ~n159 & n227;
  assign n229 = ~n153 & n228;
  assign n230 = ~n147 & n229;
  assign n231 = ~n146 & n230;
  assign n232 = ~n143 & n231;
  assign n233 = ~n140 & n232;
  assign n234 = ~n135 & n233;
  assign n235 = ~n132 & n234;
  assign n236 = ~n125 & n235;
  assign n237 = ~n119 & n236;
  assign n238 = ~n113 & n237;
  assign n239 = ~n111 & n238;
  assign n240 = ~n107 & n239;
  assign n241 = ~n106 & n240;
  assign n242 = ~n100 & n241;
  assign n243 = ~n97 & n242;
  assign n244 = ~n95 & n243;
  assign n245 = ~n90 & n244;
  assign n246 = ~n85 & n245;
  assign n247 = ~n81 & n246;
  assign n248 = ~n79 & n247;
  assign n249 = ~n74 & n248;
  assign n250 = ~n70 & n249;
  assign n251 = ~n64 & n250;
  assign r = n61 | ~n251;
  assign a1 = q & n134;
  assign n254 = n & n75;
  assign n255 = o & n254;
  assign n256 = p & n255;
  assign n257 = ~q & n256;
  assign n258 = ~p & n144;
  assign n259 = ~q & n258;
  assign n260 = ~h & ~l;
  assign n261 = m & n260;
  assign n262 = n & n261;
  assign n263 = o & n262;
  assign n264 = ~p & n263;
  assign n265 = ~q & n264;
  assign n266 = ~h & ~i;
  assign n267 = ~l & n266;
  assign n268 = m & n267;
  assign n269 = n & n268;
  assign n270 = o & n269;
  assign n271 = ~q & n270;
  assign n272 = ~e & ~f;
  assign n273 = ~m & n272;
  assign n274 = ~n & n273;
  assign n275 = ~o & n274;
  assign n276 = p & n275;
  assign n277 = q & n276;
  assign n278 = ~i & n272;
  assign n279 = ~l & n278;
  assign n280 = m & n279;
  assign n281 = n & n280;
  assign n282 = o & n281;
  assign n283 = p & n282;
  assign n284 = ~q & n283;
  assign n285 = ~c & ~e;
  assign n286 = ~i & n285;
  assign n287 = ~l & n286;
  assign n288 = m & n287;
  assign n289 = n & n288;
  assign n290 = o & n289;
  assign n291 = p & n290;
  assign n292 = ~q & n291;
  assign n293 = b & ~e;
  assign n294 = ~i & n293;
  assign n295 = ~l & n294;
  assign n296 = m & n295;
  assign n297 = n & n296;
  assign n298 = o & n297;
  assign n299 = p & n298;
  assign n300 = ~q & n299;
  assign n301 = a & ~e;
  assign n302 = ~f & n301;
  assign n303 = l & n302;
  assign n304 = ~m & n303;
  assign n305 = ~n & n304;
  assign n306 = o & n305;
  assign n307 = ~p & n306;
  assign n308 = ~q & n307;
  assign n309 = ~n300 & ~n308;
  assign n310 = ~n292 & n309;
  assign n311 = ~n284 & n310;
  assign n312 = ~n277 & n311;
  assign n313 = ~n271 & n312;
  assign n314 = ~n265 & n313;
  assign n315 = ~n259 & n314;
  assign n316 = ~n257 & n315;
  assign s = a1 | ~n316;
  assign n318 = ~n147 & n226;
  assign n319 = ~n146 & n318;
  assign n320 = ~n135 & n319;
  assign n321 = ~n132 & n320;
  assign n322 = ~n119 & n321;
  assign n323 = ~n113 & n322;
  assign n324 = ~n111 & n323;
  assign n325 = ~n107 & n324;
  assign n326 = ~n106 & n325;
  assign n327 = ~n100 & n326;
  assign n328 = ~n97 & n327;
  assign n329 = ~n95 & n328;
  assign n330 = ~n90 & n329;
  assign n331 = ~n85 & n330;
  assign n332 = ~n81 & n331;
  assign n333 = ~n79 & n332;
  assign n334 = ~n74 & n333;
  assign n335 = ~n70 & n334;
  assign n336 = ~n64 & n335;
  assign t = n61 | ~n336;
  assign n338 = p & n98;
  assign n339 = ~q & n338;
  assign n340 = q & n60;
  assign c0 = q & n142;
  assign n342 = n & n91;
  assign n343 = ~o & n342;
  assign n344 = ~p & n343;
  assign n345 = q & n344;
  assign n346 = q & n256;
  assign n347 = ~o & n254;
  assign n348 = ~p & n347;
  assign n349 = q & n348;
  assign n350 = ~n346 & ~n349;
  assign n351 = ~n345 & n350;
  assign n352 = ~c0 & n351;
  assign n353 = ~n340 & n352;
  assign u = n339 | ~n353;
  assign n355 = c & g;
  assign n356 = ~l & n355;
  assign n357 = m & n356;
  assign n358 = ~n & n357;
  assign n359 = o & n358;
  assign n360 = p & n359;
  assign n361 = ~q & n360;
  assign n362 = g & i;
  assign n363 = ~l & n362;
  assign n364 = m & n363;
  assign n365 = ~n & n364;
  assign n366 = o & n365;
  assign n367 = p & n366;
  assign n368 = ~q & n367;
  assign n369 = g & k;
  assign n370 = ~l & n369;
  assign n371 = m & n370;
  assign n372 = ~n & n371;
  assign n373 = o & n372;
  assign n374 = p & n373;
  assign n375 = ~q & n374;
  assign n376 = d & ~i;
  assign n377 = ~l & n376;
  assign n378 = ~m & n377;
  assign n379 = n & n378;
  assign n380 = ~o & n379;
  assign n381 = p & n380;
  assign n382 = q & n381;
  assign n383 = ~k & ~l;
  assign n384 = ~m & n383;
  assign n385 = ~n & n384;
  assign n386 = o & n385;
  assign n387 = p & n386;
  assign b0 = q & n387;
  assign n389 = ~d & ~i;
  assign n390 = ~l & n389;
  assign n391 = ~m & n390;
  assign n392 = n & n391;
  assign n393 = ~o & n392;
  assign n394 = p & n393;
  assign n395 = q & n394;
  assign n396 = ~b0 & ~n395;
  assign n397 = ~n382 & n396;
  assign n398 = ~n375 & n397;
  assign n399 = ~n368 & n398;
  assign n400 = ~n361 & n399;
  assign n401 = ~n349 & n400;
  assign n402 = ~n346 & n401;
  assign n403 = ~n159 & n402;
  assign n404 = ~n345 & n403;
  assign n405 = ~c0 & n404;
  assign n406 = ~n340 & n405;
  assign n407 = ~n143 & n406;
  assign n408 = ~n140 & n407;
  assign n409 = ~n125 & n408;
  assign v = n339 | ~n409;
  assign n411 = ~n140 & n406;
  assign n412 = ~n125 & n411;
  assign y = n339 | ~n412;
  assign z = n111 | n113;
  assign n415 = ~c0 & ~b0;
  assign n416 = ~n140 & n415;
  assign a0 = n125 | ~n416;
  assign n418 = h & j;
  assign n419 = ~l & n418;
  assign n420 = m & n419;
  assign n421 = n & n420;
  assign n422 = o & n421;
  assign n423 = ~p & n422;
  assign b1 = ~q & n423;
  assign n425 = ~p & n133;
  assign n426 = ~q & n425;
  assign n427 = o & n342;
  assign n428 = p & n427;
  assign n429 = q & n428;
  assign c1 = n426 | n429;
  assign n431 = ~q & n88;
  assign d1 = q & n73;
  assign n433 = q & n338;
  assign n434 = p & n58;
  assign n435 = ~q & n434;
  assign n436 = o & n71;
  assign n437 = ~p & n436;
  assign n438 = ~q & n437;
  assign n439 = ~q & n62;
  assign n440 = ~p & n62;
  assign n441 = q & n440;
  assign n442 = ~p & n93;
  assign n443 = q & n442;
  assign z0 = q & n425;
  assign n445 = ~q & n348;
  assign n446 = ~a & l;
  assign n447 = ~n & n446;
  assign n448 = o & n447;
  assign n449 = ~p & n448;
  assign n450 = k & ~l;
  assign n451 = ~m & n450;
  assign n452 = ~n & n451;
  assign n453 = o & n452;
  assign n454 = p & n453;
  assign n455 = q & n454;
  assign n456 = ~b & c;
  assign n457 = f & n456;
  assign n458 = h & n457;
  assign n459 = ~i & n458;
  assign n460 = ~l & n459;
  assign n461 = m & n460;
  assign n462 = n & n461;
  assign n463 = o & n462;
  assign n464 = p & n463;
  assign n465 = ~q & n464;
  assign n466 = m & n;
  assign n467 = ~o & n466;
  assign n468 = p & n467;
  assign n469 = ~q & n468;
  assign n470 = ~n308 & ~n465;
  assign n471 = ~n220 & n470;
  assign n472 = ~n211 & n471;
  assign n473 = ~n201 & n472;
  assign n474 = ~n300 & n473;
  assign n475 = ~n292 & n474;
  assign n476 = ~n284 & n475;
  assign n477 = ~n277 & n476;
  assign n478 = ~n455 & n477;
  assign n479 = ~n271 & n478;
  assign n480 = ~n449 & n479;
  assign n481 = ~n445 & n480;
  assign n482 = ~n265 & n481;
  assign n483 = ~z0 & n482;
  assign n484 = ~n443 & n483;
  assign n485 = ~n441 & n484;
  assign n486 = ~n439 & n485;
  assign n487 = ~n438 & n486;
  assign n488 = ~n435 & n487;
  assign n489 = ~n257 & n488;
  assign n490 = ~n433 & n489;
  assign n491 = ~d1 & n490;
  assign n492 = ~a1 & n491;
  assign n493 = ~n426 & n492;
  assign n494 = ~n346 & n493;
  assign n495 = ~n431 & n494;
  assign n496 = ~n159 & n495;
  assign n497 = ~n340 & n496;
  assign n498 = ~n135 & n497;
  assign n499 = ~n132 & n498;
  assign n500 = ~n119 & n499;
  assign n501 = ~n97 & n500;
  assign n502 = ~n79 & n501;
  assign n503 = ~n74 & n502;
  assign n504 = ~n64 & n503;
  assign n505 = ~n61 & n504;
  assign d0 = n469 | ~n505;
  assign n507 = ~m & n;
  assign n508 = o & n507;
  assign n509 = ~p & n508;
  assign n510 = ~q & n509;
  assign n511 = m & n101;
  assign n512 = n & n511;
  assign n513 = o & n512;
  assign n514 = p & n513;
  assign n515 = ~q & n514;
  assign n516 = p & n347;
  assign n517 = ~q & n516;
  assign n518 = ~o & n91;
  assign n519 = ~p & n518;
  assign n520 = q & n519;
  assign n521 = ~q & n344;
  assign n522 = n & n65;
  assign n523 = o & n522;
  assign n524 = p & n523;
  assign n525 = q & n524;
  assign n526 = n & n136;
  assign n527 = p & n526;
  assign n528 = q & n527;
  assign n529 = ~p & n254;
  assign n530 = q & n529;
  assign n531 = h & ~l;
  assign n532 = m & n531;
  assign n533 = n & n532;
  assign n534 = o & n533;
  assign n535 = ~p & n534;
  assign n536 = ~q & n535;
  assign n537 = ~p & n68;
  assign n538 = ~q & n537;
  assign n539 = ~j & n193;
  assign n540 = ~l & n539;
  assign n541 = m & n540;
  assign n542 = n & n541;
  assign n543 = o & n542;
  assign n544 = p & n543;
  assign n545 = ~j & n203;
  assign n546 = ~l & n545;
  assign n547 = m & n546;
  assign n548 = n & n547;
  assign n549 = o & n548;
  assign n550 = p & n549;
  assign n551 = ~j & n212;
  assign n552 = ~l & n551;
  assign n553 = m & n552;
  assign n554 = n & n553;
  assign n555 = o & n554;
  assign n556 = p & n555;
  assign n557 = ~c & g;
  assign n558 = ~i & n557;
  assign n559 = ~k & n558;
  assign n560 = ~l & n559;
  assign n561 = m & n560;
  assign n562 = ~n & n561;
  assign n563 = o & n562;
  assign n564 = p & n563;
  assign n565 = ~q & n564;
  assign n566 = ~n465 & ~n565;
  assign n567 = ~n556 & n566;
  assign n568 = ~n550 & n567;
  assign n569 = ~n544 & n568;
  assign n570 = ~n455 & n569;
  assign n571 = ~n538 & n570;
  assign n572 = ~n536 & n571;
  assign n573 = ~n530 & n572;
  assign n574 = ~n528 & n573;
  assign n575 = ~n525 & n574;
  assign n576 = ~n521 & n575;
  assign n577 = ~n520 & n576;
  assign n578 = ~n517 & n577;
  assign n579 = ~n439 & n578;
  assign n580 = ~n515 & n579;
  assign n581 = ~n395 & n580;
  assign n582 = ~n435 & n581;
  assign n583 = ~n510 & n582;
  assign n584 = ~d1 & n583;
  assign n585 = ~a1 & n584;
  assign n586 = ~n346 & n585;
  assign n587 = ~n153 & n586;
  assign n588 = ~n340 & n587;
  assign n589 = ~n140 & n588;
  assign n590 = ~n125 & n589;
  assign n591 = ~n339 & n590;
  assign n592 = ~n119 & n591;
  assign n593 = ~n100 & n592;
  assign n594 = ~n95 & n593;
  assign n595 = ~n85 & n594;
  assign n596 = ~n74 & n595;
  assign n597 = ~n70 & n596;
  assign e0 = n64 | ~n597;
  assign n599 = q & n516;
  assign n600 = p & n343;
  assign n601 = ~q & n600;
  assign n602 = f & n301;
  assign n603 = l & n602;
  assign n604 = ~m & n603;
  assign n605 = ~n & n604;
  assign n606 = o & n605;
  assign n607 = ~q & n606;
  assign n608 = f & n293;
  assign n609 = ~l & n608;
  assign n610 = ~m & n609;
  assign n611 = ~n & n610;
  assign n612 = ~o & n611;
  assign n613 = p & n612;
  assign n614 = q & n613;
  assign n615 = n566 & ~n614;
  assign n616 = ~n607 & n615;
  assign n617 = ~n556 & n616;
  assign n618 = ~n550 & n617;
  assign n619 = ~n544 & n618;
  assign n620 = ~n538 & n619;
  assign n621 = ~n536 & n620;
  assign n622 = ~n445 & n621;
  assign n623 = ~n528 & n622;
  assign n624 = ~n525 & n623;
  assign n625 = ~n601 & n624;
  assign n626 = ~n521 & n625;
  assign n627 = ~n443 & n626;
  assign n628 = ~n515 & n627;
  assign n629 = ~n599 & n628;
  assign n630 = ~b0 & n629;
  assign n631 = ~n433 & n630;
  assign n632 = ~n382 & n631;
  assign n633 = ~n375 & n632;
  assign n634 = ~n368 & n633;
  assign n635 = ~n361 & n634;
  assign n636 = ~n510 & n635;
  assign n637 = ~d1 & n636;
  assign n638 = ~a1 & n637;
  assign n639 = ~n165 & n638;
  assign n640 = ~n426 & n639;
  assign n641 = ~n431 & n640;
  assign n642 = ~n159 & n641;
  assign n643 = ~n345 & n642;
  assign n644 = ~c0 & n643;
  assign n645 = ~n153 & n644;
  assign n646 = ~n143 & n645;
  assign n647 = ~n119 & n646;
  assign n648 = ~n106 & n647;
  assign n649 = ~n97 & n648;
  assign n650 = ~n95 & n649;
  assign n651 = ~n90 & n650;
  assign n652 = ~n81 & n651;
  assign f0 = n61 | ~n652;
  assign n654 = p & n59;
  assign n655 = ~n308 & ~n565;
  assign n656 = ~n556 & n655;
  assign n657 = ~n550 & n656;
  assign n658 = ~n544 & n657;
  assign n659 = ~n300 & n658;
  assign n660 = ~n292 & n659;
  assign n661 = ~n284 & n660;
  assign n662 = ~n277 & n661;
  assign n663 = ~n538 & n662;
  assign n664 = ~n536 & n663;
  assign n665 = ~n271 & n664;
  assign n666 = ~n449 & n665;
  assign n667 = ~n265 & n666;
  assign n668 = ~n530 & n667;
  assign n669 = ~n528 & n668;
  assign n670 = ~n525 & n669;
  assign n671 = ~n601 & n670;
  assign n672 = ~n192 & n671;
  assign n673 = ~n517 & n672;
  assign n674 = ~n441 & n673;
  assign n675 = ~n438 & n674;
  assign n676 = ~n185 & n675;
  assign n677 = ~n178 & n676;
  assign n678 = ~n515 & n677;
  assign n679 = ~n599 & n678;
  assign n680 = ~n395 & n679;
  assign n681 = ~n435 & n680;
  assign n682 = ~n257 & n681;
  assign n683 = ~n433 & n682;
  assign n684 = ~n654 & n683;
  assign n685 = ~n382 & n684;
  assign n686 = ~n375 & n685;
  assign n687 = ~n368 & n686;
  assign n688 = ~n361 & n687;
  assign n689 = ~a1 & n688;
  assign n690 = ~n426 & n689;
  assign n691 = ~n153 & n690;
  assign n692 = ~n147 & n691;
  assign n693 = ~n340 & n692;
  assign n694 = ~n132 & n693;
  assign n695 = ~n113 & n694;
  assign n696 = ~n111 & n695;
  assign n697 = ~n106 & n696;
  assign n698 = ~n97 & n697;
  assign n699 = ~n85 & n698;
  assign n700 = ~n81 & n699;
  assign n701 = ~n79 & n700;
  assign n702 = ~n70 & n701;
  assign n703 = ~n64 & n702;
  assign g0 = n61 | ~n703;
  assign n705 = ~c & ~g;
  assign n706 = ~i & n705;
  assign n707 = ~l & n706;
  assign n708 = n & n707;
  assign n709 = o & n708;
  assign n710 = p & n709;
  assign n711 = q & n710;
  assign n712 = ~n565 & ~n614;
  assign n713 = ~n607 & n712;
  assign n714 = ~n556 & n713;
  assign n715 = ~n550 & n714;
  assign n716 = ~n544 & n715;
  assign n717 = ~b1 & n716;
  assign n718 = ~n455 & n717;
  assign n719 = ~n520 & n718;
  assign n720 = ~n517 & n719;
  assign n721 = ~z0 & n720;
  assign n722 = ~n443 & n721;
  assign n723 = ~n441 & n722;
  assign n724 = ~n515 & n723;
  assign n725 = ~n429 & n724;
  assign n726 = ~n599 & n725;
  assign n727 = ~n654 & n726;
  assign n728 = ~n171 & n727;
  assign n729 = ~n382 & n728;
  assign n730 = ~n375 & n729;
  assign n731 = ~n368 & n730;
  assign n732 = ~n361 & n731;
  assign n733 = ~n510 & n732;
  assign n734 = ~d1 & n733;
  assign n735 = ~n165 & n734;
  assign n736 = ~n426 & n735;
  assign n737 = ~n431 & n736;
  assign n738 = ~c0 & n737;
  assign n739 = ~n153 & n738;
  assign n740 = ~n147 & n739;
  assign n741 = ~n146 & n740;
  assign n742 = ~n340 & n741;
  assign n743 = ~n135 & n742;
  assign n744 = ~n339 & n743;
  assign n745 = ~n113 & n744;
  assign n746 = ~n97 & n745;
  assign n747 = ~n90 & n746;
  assign n748 = ~n85 & n747;
  assign n749 = ~n79 & n748;
  assign n750 = ~n74 & n749;
  assign n751 = ~n70 & n750;
  assign n752 = ~n61 & n751;
  assign h0 = n711 | ~n752;
  assign n754 = ~c & ~l;
  assign n755 = ~m & n754;
  assign n756 = ~n & n755;
  assign n757 = ~o & n756;
  assign n758 = ~p & n757;
  assign n759 = ~n465 & ~n614;
  assign n760 = ~n607 & n759;
  assign n761 = ~n220 & n760;
  assign n762 = ~n211 & n761;
  assign n763 = ~n201 & n762;
  assign n764 = ~n445 & n763;
  assign n765 = ~n259 & n764;
  assign n766 = ~n521 & n765;
  assign n767 = ~n441 & n766;
  assign n768 = ~n439 & n767;
  assign n769 = ~n515 & n768;
  assign n770 = ~n599 & n769;
  assign n771 = ~n395 & n770;
  assign n772 = ~n433 & n771;
  assign n773 = ~n654 & n772;
  assign n774 = ~n510 & n773;
  assign n775 = ~n349 & n774;
  assign n776 = ~n165 & n775;
  assign n777 = ~n431 & n776;
  assign n778 = ~n146 & n777;
  assign n779 = ~n143 & n778;
  assign n780 = ~n135 & n779;
  assign n781 = ~n132 & n780;
  assign n782 = ~n339 & n781;
  assign n783 = ~n113 & n782;
  assign n784 = ~n111 & n783;
  assign n785 = ~n100 & n784;
  assign n786 = ~n97 & n785;
  assign n787 = ~n90 & n786;
  assign n788 = ~n85 & n787;
  assign n789 = ~n81 & n788;
  assign n790 = ~n74 & n789;
  assign n791 = ~n70 & n790;
  assign n792 = ~n61 & n791;
  assign i0 = n758 | ~n792;
  assign n794 = ~n271 & n311;
  assign n795 = ~n265 & n794;
  assign n796 = ~n259 & n795;
  assign n797 = ~n438 & n796;
  assign j0 = n257 | ~n797;
  assign n799 = n311 & ~b1;
  assign n800 = ~n271 & n799;
  assign n801 = ~n265 & n800;
  assign n802 = ~n259 & n801;
  assign n803 = ~n438 & n802;
  assign n804 = ~n429 & n803;
  assign n805 = ~n257 & n804;
  assign n806 = ~d1 & n805;
  assign n807 = ~n426 & n806;
  assign n808 = ~n159 & n807;
  assign n809 = ~n140 & n808;
  assign n810 = ~n132 & n809;
  assign n811 = ~n125 & n810;
  assign n812 = ~n119 & n811;
  assign n813 = ~n107 & n812;
  assign n814 = ~n106 & n813;
  assign n815 = ~n100 & n814;
  assign n816 = ~n95 & n815;
  assign n817 = ~n90 & n816;
  assign n818 = ~n85 & n817;
  assign n819 = ~n81 & n818;
  assign n820 = ~n79 & n819;
  assign n821 = ~n74 & n820;
  assign n822 = ~n70 & n821;
  assign n823 = ~n64 & n822;
  assign k0 = n61 | ~n823;
  assign n825 = ~b1 & ~z0;
  assign n826 = ~b0 & n825;
  assign n827 = ~n171 & n826;
  assign n828 = ~d1 & n827;
  assign n829 = ~a1 & n828;
  assign n830 = ~n165 & n829;
  assign n831 = ~c0 & n830;
  assign n832 = ~n153 & n831;
  assign n833 = ~n146 & n832;
  assign n834 = ~n143 & n833;
  assign n835 = ~n140 & n834;
  assign n836 = ~n125 & n835;
  assign n837 = ~n113 & n836;
  assign n838 = ~n111 & n837;
  assign n839 = ~n107 & n838;
  assign n840 = ~n106 & n839;
  assign n841 = ~n100 & n840;
  assign n842 = ~n97 & n841;
  assign n843 = ~n95 & n842;
  assign n844 = ~n85 & n843;
  assign n845 = ~n81 & n844;
  assign n846 = ~n79 & n845;
  assign n847 = ~n74 & n846;
  assign n848 = ~n70 & n847;
  assign n849 = ~n64 & n848;
  assign l0 = n61 | ~n849;
  assign n851 = ~n185 & ~n192;
  assign n852 = ~n178 & n851;
  assign n853 = ~n429 & n852;
  assign n854 = ~n171 & n853;
  assign n855 = ~n426 & n854;
  assign n856 = ~n159 & n855;
  assign n857 = ~n147 & n856;
  assign n858 = ~n146 & n857;
  assign n859 = ~n132 & n858;
  assign n860 = ~n119 & n859;
  assign n861 = ~n113 & n860;
  assign n862 = ~n111 & n861;
  assign n863 = ~n107 & n862;
  assign n864 = ~n100 & n863;
  assign n865 = ~n90 & n864;
  assign n866 = ~n85 & n865;
  assign n867 = ~n79 & n866;
  assign n868 = ~n70 & n867;
  assign m0 = n61 | ~n868;
  assign n870 = ~n429 & n825;
  assign n871 = ~b0 & n870;
  assign n872 = ~d1 & n871;
  assign n873 = ~a1 & n872;
  assign n874 = ~n165 & n873;
  assign n875 = ~n426 & n874;
  assign n876 = ~n159 & n875;
  assign n877 = ~c0 & n876;
  assign n878 = ~n153 & n877;
  assign n879 = ~n143 & n878;
  assign n880 = ~n140 & n879;
  assign n881 = ~n132 & n880;
  assign n882 = ~n125 & n881;
  assign n883 = ~n119 & n882;
  assign n884 = ~n107 & n883;
  assign n885 = ~n106 & n884;
  assign n886 = ~n100 & n885;
  assign n887 = ~n97 & n886;
  assign n888 = ~n95 & n887;
  assign n889 = ~n90 & n888;
  assign n890 = ~n85 & n889;
  assign n891 = ~n81 & n890;
  assign n892 = ~n79 & n891;
  assign n893 = ~n74 & n892;
  assign n894 = ~n70 & n893;
  assign n895 = ~n64 & n894;
  assign n0 = n61 | ~n895;
  assign n897 = ~n220 & ~n308;
  assign n898 = ~n211 & n897;
  assign n899 = ~n201 & n898;
  assign n900 = ~n300 & n899;
  assign n901 = ~n292 & n900;
  assign n902 = ~n284 & n901;
  assign n903 = ~b1 & n902;
  assign n904 = ~n271 & n903;
  assign n905 = ~n265 & n904;
  assign n906 = ~n259 & n905;
  assign n907 = ~n192 & n906;
  assign n908 = ~z0 & n907;
  assign n909 = ~n438 & n908;
  assign n910 = ~n185 & n909;
  assign n911 = ~n178 & n910;
  assign n912 = ~n257 & n911;
  assign n913 = ~b0 & n912;
  assign n914 = ~n171 & n913;
  assign n915 = ~n143 & n914;
  assign n916 = ~n140 & n915;
  assign n917 = ~n125 & n916;
  assign n918 = ~n111 & n917;
  assign n919 = ~n106 & n918;
  assign n920 = ~n97 & n919;
  assign n921 = ~n95 & n920;
  assign o0 = n64 | ~n921;
  assign n923 = ~n382 & ~n395;
  assign n924 = ~n375 & n923;
  assign n925 = ~n368 & n924;
  assign n926 = ~n361 & n925;
  assign n927 = ~n349 & n926;
  assign n928 = ~n346 & n927;
  assign n929 = ~n159 & n928;
  assign n930 = ~n345 & n929;
  assign n931 = ~n140 & n930;
  assign n932 = ~n132 & n931;
  assign n933 = ~n125 & n932;
  assign n934 = ~n339 & n933;
  assign n935 = ~n119 & n934;
  assign n936 = ~n107 & n935;
  assign n937 = ~n106 & n936;
  assign n938 = ~n100 & n937;
  assign n939 = ~n95 & n938;
  assign n940 = ~n90 & n939;
  assign n941 = ~n85 & n940;
  assign n942 = ~n81 & n941;
  assign n943 = ~n79 & n942;
  assign n944 = ~n74 & n943;
  assign n945 = ~n70 & n944;
  assign n946 = ~n64 & n945;
  assign p0 = n61 | ~n946;
  assign n948 = n222 & ~n395;
  assign n949 = ~b0 & n948;
  assign n950 = ~n382 & n949;
  assign n951 = ~n375 & n950;
  assign n952 = ~n368 & n951;
  assign n953 = ~n361 & n952;
  assign n954 = ~n349 & n953;
  assign n955 = ~n165 & n954;
  assign n956 = ~n345 & n955;
  assign n957 = ~c0 & n956;
  assign n958 = ~n153 & n957;
  assign n959 = ~n340 & n958;
  assign n960 = ~n143 & n959;
  assign n961 = ~n140 & n960;
  assign n962 = ~n135 & n961;
  assign n963 = ~n132 & n962;
  assign n964 = ~n125 & n963;
  assign n965 = ~n339 & n964;
  assign n966 = ~n113 & n965;
  assign n967 = ~n111 & n966;
  assign n968 = ~n107 & n967;
  assign n969 = ~n106 & n968;
  assign n970 = ~n100 & n969;
  assign n971 = ~n95 & n970;
  assign n972 = ~n85 & n971;
  assign n973 = ~n81 & n972;
  assign n974 = ~n79 & n973;
  assign n975 = ~n74 & n974;
  assign n976 = ~n70 & n975;
  assign n977 = ~n64 & n976;
  assign q0 = n61 | ~n977;
  assign n979 = ~n395 & n852;
  assign n980 = ~b0 & n979;
  assign n981 = ~n349 & n980;
  assign n982 = ~n165 & n981;
  assign n983 = ~n346 & n982;
  assign n984 = ~n159 & n983;
  assign n985 = ~n345 & n984;
  assign n986 = ~c0 & n985;
  assign n987 = ~n153 & n986;
  assign n988 = ~n147 & n987;
  assign n989 = ~n340 & n988;
  assign n990 = ~n143 & n989;
  assign n991 = ~n119 & n990;
  assign n992 = ~n113 & n991;
  assign n993 = ~n111 & n992;
  assign n994 = ~n107 & n993;
  assign n995 = ~n95 & n994;
  assign n996 = ~n90 & n995;
  assign n997 = ~n85 & n996;
  assign n998 = ~n70 & n997;
  assign r0 = n61 | ~n998;
  assign n1000 = ~n382 & n948;
  assign n1001 = ~n375 & n1000;
  assign n1002 = ~n368 & n1001;
  assign n1003 = ~n361 & n1002;
  assign n1004 = ~n349 & n1003;
  assign n1005 = ~n346 & n1004;
  assign n1006 = ~n159 & n1005;
  assign n1007 = ~n345 & n1006;
  assign n1008 = ~n140 & n1007;
  assign n1009 = ~n135 & n1008;
  assign n1010 = ~n132 & n1009;
  assign n1011 = ~n125 & n1010;
  assign n1012 = ~n339 & n1011;
  assign n1013 = ~n119 & n1012;
  assign n1014 = ~n107 & n1013;
  assign n1015 = ~n106 & n1014;
  assign n1016 = ~n100 & n1015;
  assign n1017 = ~n95 & n1016;
  assign n1018 = ~n90 & n1017;
  assign n1019 = ~n85 & n1018;
  assign n1020 = ~n81 & n1019;
  assign n1021 = ~n79 & n1020;
  assign n1022 = ~n74 & n1021;
  assign n1023 = ~n70 & n1022;
  assign n1024 = ~n64 & n1023;
  assign s0 = n61 | ~n1024;
  assign n1026 = n225 & ~b0;
  assign n1027 = ~n171 & n1026;
  assign n1028 = ~n382 & n1027;
  assign n1029 = ~n375 & n1028;
  assign n1030 = ~n368 & n1029;
  assign n1031 = ~n361 & n1030;
  assign n1032 = ~n340 & n1031;
  assign n1033 = ~n143 & n1032;
  assign n1034 = ~n140 & n1033;
  assign n1035 = ~n125 & n1034;
  assign n1036 = ~n339 & n1035;
  assign n1037 = ~n111 & n1036;
  assign n1038 = ~n106 & n1037;
  assign n1039 = ~n100 & n1038;
  assign n1040 = ~n97 & n1039;
  assign n1041 = ~n79 & n1040;
  assign t0 = n64 | ~n1041;
  assign n1043 = ~n171 & n222;
  assign n1044 = ~n346 & n1043;
  assign n1045 = ~n159 & n1044;
  assign n1046 = ~n146 & n1045;
  assign n1047 = ~n140 & n1046;
  assign n1048 = ~n135 & n1047;
  assign n1049 = ~n132 & n1048;
  assign n1050 = ~n125 & n1049;
  assign n1051 = ~n119 & n1050;
  assign n1052 = ~n107 & n1051;
  assign n1053 = ~n106 & n1052;
  assign n1054 = ~n100 & n1053;
  assign n1055 = ~n97 & n1054;
  assign n1056 = ~n95 & n1055;
  assign n1057 = ~n90 & n1056;
  assign n1058 = ~n85 & n1057;
  assign n1059 = ~n81 & n1058;
  assign n1060 = ~n79 & n1059;
  assign n1061 = ~n74 & n1060;
  assign n1062 = ~n70 & n1061;
  assign n1063 = ~n64 & n1062;
  assign u0 = n61 | ~n1063;
  assign n1065 = ~n345 & n927;
  assign n1066 = ~n340 & n1065;
  assign n1067 = ~n140 & n1066;
  assign n1068 = ~n132 & n1067;
  assign n1069 = ~n125 & n1068;
  assign n1070 = ~n339 & n1069;
  assign n1071 = ~n119 & n1070;
  assign n1072 = ~n113 & n1071;
  assign n1073 = ~n111 & n1072;
  assign n1074 = ~n90 & n1073;
  assign n1075 = ~n85 & n1074;
  assign n1076 = ~n81 & n1075;
  assign n1077 = ~n79 & n1076;
  assign n1078 = ~n74 & n1077;
  assign v0 = n70 | ~n1078;
  assign n1080 = ~n147 & n852;
  assign n1081 = ~n340 & n1080;
  assign n1082 = ~n107 & n1081;
  assign n1083 = ~n106 & n1082;
  assign n1084 = ~n64 & n1083;
  assign w0 = n61 | ~n1084;
  assign n1086 = ~n382 & n979;
  assign n1087 = ~n375 & n1086;
  assign n1088 = ~n368 & n1087;
  assign n1089 = ~n361 & n1088;
  assign n1090 = ~n349 & n1089;
  assign n1091 = ~n346 & n1090;
  assign n1092 = ~n345 & n1091;
  assign n1093 = ~n147 & n1092;
  assign n1094 = ~n339 & n1093;
  assign n1095 = ~n107 & n1094;
  assign n1096 = ~n106 & n1095;
  assign n1097 = ~n64 & n1096;
  assign x0 = n61 | ~n1097;
  assign n1099 = ~n165 & n1090;
  assign n1100 = ~n345 & n1099;
  assign n1101 = ~c0 & n1100;
  assign n1102 = ~n153 & n1101;
  assign n1103 = ~n132 & n1102;
  assign n1104 = ~n339 & n1103;
  assign n1105 = ~n119 & n1104;
  assign n1106 = ~n111 & n1105;
  assign n1107 = ~n107 & n1106;
  assign n1108 = ~n106 & n1107;
  assign n1109 = ~n90 & n1108;
  assign n1110 = ~n81 & n1109;
  assign n1111 = ~n74 & n1110;
  assign n1112 = ~n64 & n1111;
  assign y0 = n61 | ~n1112;
  assign w = t;
  assign x = t;
endmodule


