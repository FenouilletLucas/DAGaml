// Benchmark "x1" written by ABC on Tue May 16 16:07:53 2017

module x1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0,
    a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2, i1, i2,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0;
  output a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2, i1,
    i2, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1;
  wire n87, n88, n89, n91, n92, n93, n94, n95, n96, n97, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n133, n135, n136, n137, n138, n139, n140,
    n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n186, n187, n188, n189, n190, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n231,
    n232, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n250, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n329, n330, n331, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n357, n358,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n388, n389, n391, n392, n393;
  assign n87 = ~j & ~v;
  assign n88 = b & l;
  assign n89 = ~n & n88;
  assign a2 = f0 | r0;
  assign n91 = ~r & a0;
  assign n92 = n87 & n91;
  assign n93 = a0 & ~n89;
  assign n94 = ~b & a2;
  assign n95 = m & a0;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~n93 & n96;
  assign a1 = n92 | ~n97;
  assign n99 = ~a & ~m;
  assign n100 = ~j & v;
  assign n101 = k0 & n99;
  assign n102 = n100 & n101;
  assign n103 = j & g0;
  assign n104 = ~k & a0;
  assign n105 = n99 & n104;
  assign n106 = ~n87 & n105;
  assign n107 = n89 & n106;
  assign n108 = b & ~n;
  assign n109 = n102 & n108;
  assign n110 = o0 & t0;
  assign n111 = c & ~w;
  assign n112 = n103 & n111;
  assign n113 = ~n110 & ~n112;
  assign n114 = ~n109 & n113;
  assign b1 = n107 | ~n114;
  assign n116 = ~p & ~v;
  assign n117 = ~e & ~u;
  assign n118 = ~w & n117;
  assign n119 = n99 & n118;
  assign n120 = o & n119;
  assign n121 = ~g & ~v;
  assign n122 = p0 & n120;
  assign n123 = n116 & n122;
  assign n124 = e0 & n120;
  assign n125 = n116 & n124;
  assign n126 = p0 & n121;
  assign n127 = n120 & n126;
  assign n128 = e0 & n121;
  assign n129 = n120 & n128;
  assign n130 = ~n127 & ~n129;
  assign n131 = ~n125 & n130;
  assign b2 = n123 | ~n131;
  assign n133 = m & ~v;
  assign c1 = b0 & ~n133;
  assign n135 = ~h & n99;
  assign n136 = o & p;
  assign n137 = c0 & ~n133;
  assign n138 = ~d & ~v;
  assign n139 = d0 & n138;
  assign n140 = ~n136 & n139;
  assign n141 = n135 & n140;
  assign d1 = n137 | n141;
  assign n143 = q & n136;
  assign n144 = g & ~v;
  assign n145 = q0 & n144;
  assign n146 = ~n143 & n145;
  assign n147 = g & p0;
  assign n148 = ~n143 & n147;
  assign n149 = v & p0;
  assign n150 = ~n148 & ~n149;
  assign n151 = ~n146 & n150;
  assign n152 = ~z & ~h0;
  assign n153 = ~a & i;
  assign n154 = ~n151 & n153;
  assign n155 = ~y & ~i0;
  assign n156 = n152 & n155;
  assign e2 = ~n154 & n156;
  assign n158 = d & d0;
  assign n159 = g & ~m;
  assign n160 = ~o & n159;
  assign n161 = ~n117 & n160;
  assign n162 = n158 & n161;
  assign n163 = ~m & ~o;
  assign n164 = n118 & n163;
  assign n165 = n158 & n164;
  assign n166 = o0 & u0;
  assign n167 = ~o & e0;
  assign n168 = n135 & n167;
  assign n169 = ~n166 & ~n168;
  assign n170 = ~n165 & n169;
  assign e1 = n162 | ~n170;
  assign n172 = e0 & n136;
  assign n173 = n135 & n172;
  assign n174 = ~i & ~q;
  assign n175 = q0 & n174;
  assign n176 = ~g & ~q;
  assign n177 = q0 & n176;
  assign n178 = ~i & ~o;
  assign n179 = q0 & n178;
  assign n180 = ~g & ~o;
  assign n181 = q0 & n180;
  assign n182 = ~n179 & ~n181;
  assign n183 = ~n177 & n182;
  assign n184 = ~n175 & n183;
  assign f1 = n173 | ~n184;
  assign n186 = ~p0 & ~s0;
  assign n187 = ~d & d0;
  assign n188 = n186 & ~n187;
  assign n189 = ~n167 & n188;
  assign n190 = h & t;
  assign s1 = i0 & n190;
  assign n192 = ~z0 & n91;
  assign n193 = ~z0 & n95;
  assign n194 = j & a0;
  assign n195 = ~z0 & n194;
  assign n196 = h & ~n189;
  assign n197 = a0 & ~n88;
  assign n198 = ~m0 & ~x0;
  assign n199 = ~s1 & n198;
  assign n200 = ~a2 & n199;
  assign n201 = ~n197 & n200;
  assign n202 = ~n196 & n201;
  assign n203 = ~n195 & n202;
  assign n204 = ~n193 & n203;
  assign f2 = ~n192 & n204;
  assign n206 = r & s;
  assign n207 = c & d;
  assign n208 = ~a & ~h;
  assign n209 = ~i & n208;
  assign n210 = p0 & n209;
  assign n211 = ~n143 & n210;
  assign n212 = ~n206 & n211;
  assign n213 = ~n121 & n212;
  assign n214 = p0 & ~n143;
  assign n215 = ~n206 & n214;
  assign n216 = n121 & n215;
  assign n217 = ~n207 & n216;
  assign n218 = n135 & n217;
  assign n219 = d0 & n136;
  assign n220 = ~n121 & n219;
  assign n221 = ~n133 & n220;
  assign n222 = n117 & n219;
  assign n223 = ~n133 & n222;
  assign n224 = o0 & v0;
  assign n225 = v & d0;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n223 & n226;
  assign n228 = ~n221 & n227;
  assign n229 = ~n218 & n228;
  assign g1 = n213 | ~n229;
  assign n231 = ~a & h;
  assign n232 = n118 & n231;
  assign h1 = ~n189 & n232;
  assign n234 = a0 & n99;
  assign n235 = ~n87 & n234;
  assign n236 = n89 & n235;
  assign n237 = n89 & n102;
  assign n238 = c & n103;
  assign n239 = i & i0;
  assign n240 = ~h & d0;
  assign n241 = ~y & ~b0;
  assign n242 = ~c0 & n241;
  assign n243 = ~n158 & n242;
  assign n244 = n152 & n243;
  assign n245 = ~n240 & n244;
  assign n246 = ~n239 & n245;
  assign n247 = ~n238 & n246;
  assign n248 = ~n237 & n247;
  assign h2 = ~n236 & n248;
  assign n250 = a & t;
  assign z1 = c0 | d0;
  assign n252 = ~v & w;
  assign n253 = n158 & n252;
  assign n254 = a & ~j;
  assign n255 = g0 & n254;
  assign n256 = i0 & n250;
  assign n257 = n133 & z1;
  assign n258 = p0 & n133;
  assign n259 = p0 & n206;
  assign n260 = l0 & n206;
  assign n261 = s0 & ~n99;
  assign n262 = q0 & ~n99;
  assign n263 = k0 & ~n99;
  assign n264 = h0 & ~n99;
  assign n265 = e0 & ~n99;
  assign n266 = b0 & ~c1;
  assign n267 = b & r0;
  assign n268 = a & p0;
  assign n269 = a & j0;
  assign n270 = m & g0;
  assign n271 = a & d0;
  assign n272 = a & a0;
  assign n273 = ~n271 & ~n272;
  assign n274 = ~n270 & n273;
  assign n275 = ~n269 & n274;
  assign n276 = ~n268 & n275;
  assign n277 = ~n267 & n276;
  assign n278 = ~n266 & n277;
  assign n279 = ~n265 & n278;
  assign n280 = ~n264 & n279;
  assign n281 = ~n263 & n280;
  assign n282 = ~n262 & n281;
  assign n283 = ~n261 & n282;
  assign n284 = ~n260 & n283;
  assign n285 = ~n259 & n284;
  assign n286 = ~n258 & n285;
  assign n287 = ~n257 & n286;
  assign n288 = ~n256 & n287;
  assign n289 = ~n255 & n288;
  assign k1 = n253 | ~n289;
  assign n291 = ~a & o;
  assign n292 = ~n117 & n291;
  assign n293 = n158 & n292;
  assign n294 = n116 & n293;
  assign n295 = e0 & n291;
  assign n296 = ~n117 & n295;
  assign n297 = n116 & n296;
  assign n298 = ~a & d0;
  assign n299 = n136 & n298;
  assign n300 = ~n117 & n299;
  assign n301 = n121 & n300;
  assign n302 = ~a & ~n117;
  assign n303 = n121 & n302;
  assign n304 = n158 & n303;
  assign n305 = ~a & e0;
  assign n306 = ~n117 & n305;
  assign n307 = n121 & n306;
  assign n308 = h & e0;
  assign n309 = ~n117 & n308;
  assign n310 = h & d0;
  assign n311 = ~n117 & n310;
  assign n312 = b & k;
  assign n313 = a0 & n312;
  assign n314 = h0 & ~n118;
  assign n315 = q0 & n143;
  assign n316 = p0 & n143;
  assign n317 = b & f0;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n315 & n318;
  assign n320 = ~n314 & n319;
  assign n321 = ~n313 & n320;
  assign n322 = ~n311 & n321;
  assign n323 = ~n309 & n322;
  assign n324 = ~n307 & n323;
  assign n325 = ~n304 & n324;
  assign n326 = ~n301 & n325;
  assign n327 = ~n297 & n326;
  assign l1 = n294 | ~n327;
  assign n329 = j & h0;
  assign n330 = n120 & n158;
  assign n331 = n116 & n330;
  assign m1 = n329 | n331;
  assign n333 = n136 & n177;
  assign n334 = n119 & n333;
  assign n335 = ~a & f;
  assign n336 = g0 & n335;
  assign n337 = n100 & n336;
  assign n338 = n119 & n126;
  assign n339 = n207 & n338;
  assign n340 = ~c & n135;
  assign n341 = n103 & n340;
  assign n342 = ~p & e0;
  assign n343 = n120 & n342;
  assign n344 = o0 & w0;
  assign n345 = n119 & n344;
  assign n346 = ~h & s0;
  assign n347 = n119 & n346;
  assign n348 = ~j & h0;
  assign n349 = n119 & n348;
  assign n350 = ~n347 & ~n349;
  assign n351 = ~n345 & n350;
  assign n352 = ~n343 & n351;
  assign n353 = ~n341 & n352;
  assign n354 = ~n339 & n353;
  assign n355 = ~n337 & n354;
  assign n1 = n334 | ~n355;
  assign n357 = i & n208;
  assign n358 = i0 & n357;
  assign o1 = n154 | n358;
  assign n360 = ~k & r;
  assign n361 = a0 & n360;
  assign n362 = n99 & n361;
  assign n363 = ~n206 & n362;
  assign n364 = n87 & n363;
  assign n365 = n88 & n364;
  assign n366 = b & r;
  assign n367 = ~n206 & n366;
  assign n368 = n87 & n367;
  assign n369 = n101 & n368;
  assign n370 = ~a & j0;
  assign n371 = ~h & ~i;
  assign n372 = i0 & n371;
  assign n373 = ~n250 & n372;
  assign n374 = ~n370 & ~n373;
  assign n375 = ~n369 & n374;
  assign r1 = n365 | ~n375;
  assign n377 = ~f & ~j;
  assign n378 = g0 & n377;
  assign n379 = n99 & n378;
  assign n380 = ~r & n87;
  assign n381 = n101 & n380;
  assign n382 = g0 & n99;
  assign n383 = n87 & n382;
  assign n384 = n & n102;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n381 & n385;
  assign v1 = n379 | ~n386;
  assign n388 = k0 & n206;
  assign n389 = a0 & n206;
  assign w1 = n388 | n389;
  assign n391 = ~g0 & ~a2;
  assign n392 = n152 & n391;
  assign n393 = j & n152;
  assign x1 = ~n392 & ~n393;
  assign d2 = ~e2;
  assign g2 = ~f2;
  assign i2 = ~h2;
  assign y1 = ~x1;
  assign c2 = h0;
  assign i1 = m0;
  assign j1 = n0;
  assign p1 = y;
  assign q1 = z;
  assign t1 = x0;
  assign u1 = y0;
endmodule


