// Benchmark "DES" written by ABC on Tue May 16 16:07:49 2017

module DES ( 
    \data<63> , \data<61> , \data<62> , \reset<0> , \outreg<58> ,
    \inreg<0> , \outreg<57> , \inreg<1> , \outreg<56> , \inreg<2> ,
    \outreg<55> , \inreg<3> , \inreg<4> , \inreg<5> , \inreg<6> ,
    \outreg<59> , \inreg<7> , \outreg<50> , \inreg<8> , \inreg<9> ,
    \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \load_key<0> ,
    \outreg<60> , \outreg<63> , \outreg<62> , \outreg<61> , \D<0> , \D<1> ,
    \D<2> , \D<3> , \D<4> , \D<5> , \D<6> , \C<10> , \D<7> , \C<11> ,
    \D<8> , \C<12> , \D<9> , \C<13> , \C<14> , \C<15> , \C<16> , \C<17> ,
    \C<18> , \C<19> , \outreg<18> , \outreg<17> , \outreg<16> ,
    \outreg<15> , \C<20> , \outreg<19> , \C<21> , \outreg<10> , \C<22> ,
    \C<23> , \C<24> , \C<25> , \outreg<14> , \C<26> , \outreg<13> ,
    \C<27> , \outreg<12> , \outreg<11> , \outreg<28> , \outreg<27> ,
    \outreg<26> , \outreg<25> , \outreg<29> , \outreg<20> , \data<3> ,
    \data<4> , \data<1> , \outreg<24> , \data<2> , \outreg<23> ,
    \outreg<22> , \data<0> , \outreg<21> , \outreg<38> , \outreg<37> ,
    \outreg<36> , \outreg<35> , \data<9> , \data<7> , \data<8> ,
    \outreg<39> , \data<5> , \outreg<30> , \data<6> , \outreg<34> ,
    \outreg<33> , \outreg<32> , \outreg<31> , \outreg<48> , \outreg<47> ,
    \outreg<46> , \outreg<45> , \outreg<49> , \outreg<40> , \outreg<44> ,
    \outreg<43> , \outreg<42> , \outreg<41> , \D<10> , \D<11> , \D<12> ,
    \D<13> , \D<14> , \D<15> , \D<16> , \D<17> , \D<18> , \D<19> , \D<20> ,
    \D<21> , \data_in<7> , \D<22> , \D<23> , \data_in<5> , \D<24> ,
    \data_in<6> , \D<25> , \D<26> , \D<27> , \data_in<0> , \data_in<3> ,
    \data_in<4> , \data_in<1> , \data_in<2> , \data<37> , \data<38> ,
    \data<35> , \data<36> , \data<39> , \data<30> , \data<33> , \data<34> ,
    \data<31> , \data<32> , \data<47> , \data<48> , \data<45> , \data<46> ,
    \data<49> , \data<40> , \data<43> , \data<44> , \data<41> , \data<42> ,
    \data<17> , \data<18> , \data<15> , \count<0> , \data<16> , \count<3> ,
    \data<19> , \count<1> , \count<2> , \data<10> , \data<13> , \data<14> ,
    \data<11> , \data<12> , \data<27> , \data<28> , \data<25> , \data<26> ,
    \data<29> , \data<20> , \data<23> , \data<24> , \data<21> , \data<22> ,
    \C<0> , \C<1> , \C<2> , \C<3> , \C<4> , \C<5> , \C<6> , \C<7> , \C<8> ,
    \C<9> , \inreg<12> , \inreg<11> , \inreg<14> , \inreg<13> ,
    \inreg<10> , \inreg<19> , \inreg<16> , \inreg<15> , \inreg<18> ,
    \inreg<17> , \inreg<22> , \inreg<21> , \inreg<24> , \inreg<23> ,
    \inreg<20> , \inreg<29> , \inreg<26> , \inreg<25> , \outreg<9> ,
    \inreg<28> , \inreg<27> , \inreg<32> , \inreg<31> , \outreg<5> ,
    \inreg<34> , \outreg<6> , \inreg<33> , \outreg<7> , \outreg<8> ,
    \outreg<1> , \inreg<30> , \outreg<2> , \outreg<3> , \outreg<4> ,
    \inreg<39> , \inreg<36> , \outreg<0> , \inreg<35> , \inreg<38> ,
    \inreg<37> , \inreg<42> , \inreg<41> , \inreg<44> , \inreg<43> ,
    \inreg<40> , \inreg<49> , \inreg<46> , \inreg<45> , \encrypt_mode<0> ,
    \inreg<48> , \inreg<47> , \inreg<52> , \inreg<51> , \inreg<54> ,
    \inreg<53> , \inreg<50> , \inreg<55> , \data<57> , \data<58> ,
    \data<55> , \data<56> , \encrypt<0> , \data<59> , \data<50> ,
    \data<53> , \data<54> , \data<51> , \data<52> , \data<60> ,
    \data_new<25> , \inreg_new<45> , \data_new<26> , \data_new<13> ,
    \data_new<14> , \data_new<11> , \inreg_new<49> , \data_new<12> ,
    \inreg_new<30> , \outreg_new<11> , \count_new<0> , \outreg_new<12> ,
    \data_new<10> , \outreg_new<13> , \outreg_new<14> , \inreg_new<34> ,
    \count_new<3> , \inreg_new<33> , \inreg_new<32> , \count_new<1> ,
    \data_new<19> , \inreg_new<31> , \count_new<2> , \outreg_new<10> ,
    \inreg_new<38> , \outreg_new<19> , \data_new<17> , \inreg_new<37> ,
    \data_new<18> , \inreg_new<36> , \data_new<15> , \inreg_new<35> ,
    \data_new<16> , \outreg_new<15> , \outreg_new<16> , \outreg_new<17> ,
    \inreg_new<39> , \outreg_new<18> , \outreg_new<21> , \outreg_new<22> ,
    \outreg_new<23> , \outreg_new<24> , \outreg_new<20> , \outreg_new<29> ,
    \outreg_new<25> , \outreg_new<26> , \outreg_new<27> , \outreg_new<28> ,
    \outreg_new<31> , \outreg_new<32> , \outreg_new<33> , \outreg_new<34> ,
    \outreg_new<30> , \outreg_new<39> , \outreg_new<35> , \outreg_new<36> ,
    \outreg_new<37> , \outreg_new<38> , \outreg_new<41> , \outreg_new<42> ,
    \outreg_new<43> , \outreg_new<44> , \outreg_new<40> , \outreg_new<49> ,
    \outreg_new<45> , \outreg_new<46> , \outreg_new<47> , \outreg_new<48> ,
    \C_new<23> , \C_new<24> , \C_new<21> , \C_new<22> , \C_new<20> ,
    \data_new<4> , \data_new<3> , \C_new<27> , \data_new<2> ,
    \data_new<1> , \C_new<25> , \data_new<0> , \C_new<26> , \C_new<13> ,
    \C_new<14> , \C_new<11> , \C_new<12> , \C_new<10> , \data_new<9> ,
    \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> ,
    \C_new<19> , \C_new<17> , \C_new<18> , \C_new<15> , \C_new<16> ,
    \D_new<13> , \D_new<14> , \D_new<11> , \D_new<12> , \D_new<10> ,
    \data_new<63> , \data_new<61> , \data_new<62> , \D_new<19> ,
    \data_new<60> , \D_new<17> , \D_new<18> , \D_new<15> , \D_new<16> ,
    \D_new<23> , \D_new<24> , \D_new<21> , \D_new<22> , \D_new<20> ,
    \data_new<53> , \data_new<54> , \data_new<51> , \data_new<52> ,
    \data_new<50> , \D_new<27> , \D_new<25> , \D_new<26> , \data_new<59> ,
    \data_new<57> , \data_new<58> , \data_new<55> , \data_new<56> ,
    \D_new<7> , \C_new<6> , \D_new<8> , \C_new<5> , \D_new<5> , \C_new<8> ,
    \D_new<6> , \C_new<7> , \C_new<9> , \D_new<9> , \D_new<0> , \C_new<0> ,
    \D_new<3> , \C_new<2> , \D_new<4> , \C_new<1> , \D_new<1> , \C_new<4> ,
    \D_new<2> , \C_new<3> , \inreg_new<50> , \inreg_new<9> ,
    \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<6> ,
    \inreg_new<51> , \inreg_new<5> , \inreg_new<8> , \inreg_new<7> ,
    \inreg_new<2> , \inreg_new<55> , \inreg_new<1> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<0> , \encrypt_mode_new<0> , \outreg_new<9> ,
    \outreg_new<51> , \outreg_new<52> , \outreg_new<53> , \outreg_new<5> ,
    \outreg_new<54> , \outreg_new<6> , \outreg_new<7> , \outreg_new<8> ,
    \outreg_new<1> , \outreg_new<50> , \outreg_new<2> , \outreg_new<59> ,
    \outreg_new<3> , \outreg_new<4> , \outreg_new<55> , \data_new<43> ,
    \outreg_new<56> , \data_new<44> , \outreg_new<0> , \outreg_new<57> ,
    \data_new<41> , \outreg_new<58> , \data_new<42> , \inreg_new<20> ,
    \outreg_new<61> , \outreg_new<62> , \data_new<40> , \outreg_new<63> ,
    \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \data_new<49> ,
    \inreg_new<21> , \outreg_new<60> , \inreg_new<28> , \data_new<47> ,
    \inreg_new<27> , \data_new<48> , \inreg_new<26> , \data_new<45> ,
    \inreg_new<25> , \data_new<46> , \data_new<33> , \data_new<34> ,
    \data_new<31> , \inreg_new<29> , \data_new<32> , \inreg_new<10> ,
    \data_new<30> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \data_new<39> , \inreg_new<11> , \inreg_new<18> , \data_new<37> ,
    \inreg_new<17> , \data_new<38> , \inreg_new<16> , \data_new<35> ,
    \inreg_new<15> , \data_new<36> , \data_new<23> , \data_new<24> ,
    \data_new<21> , \inreg_new<19> , \data_new<22> , \inreg_new<40> ,
    \data_new<20> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> ,
    \data_new<29> , \inreg_new<41> , \inreg_new<48> , \data_new<27> ,
    \inreg_new<47> , \data_new<28> , \inreg_new<46>   );
  input  \data<63> , \data<61> , \data<62> , \reset<0> , \outreg<58> ,
    \inreg<0> , \outreg<57> , \inreg<1> , \outreg<56> , \inreg<2> ,
    \outreg<55> , \inreg<3> , \inreg<4> , \inreg<5> , \inreg<6> ,
    \outreg<59> , \inreg<7> , \outreg<50> , \inreg<8> , \inreg<9> ,
    \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \load_key<0> ,
    \outreg<60> , \outreg<63> , \outreg<62> , \outreg<61> , \D<0> , \D<1> ,
    \D<2> , \D<3> , \D<4> , \D<5> , \D<6> , \C<10> , \D<7> , \C<11> ,
    \D<8> , \C<12> , \D<9> , \C<13> , \C<14> , \C<15> , \C<16> , \C<17> ,
    \C<18> , \C<19> , \outreg<18> , \outreg<17> , \outreg<16> ,
    \outreg<15> , \C<20> , \outreg<19> , \C<21> , \outreg<10> , \C<22> ,
    \C<23> , \C<24> , \C<25> , \outreg<14> , \C<26> , \outreg<13> ,
    \C<27> , \outreg<12> , \outreg<11> , \outreg<28> , \outreg<27> ,
    \outreg<26> , \outreg<25> , \outreg<29> , \outreg<20> , \data<3> ,
    \data<4> , \data<1> , \outreg<24> , \data<2> , \outreg<23> ,
    \outreg<22> , \data<0> , \outreg<21> , \outreg<38> , \outreg<37> ,
    \outreg<36> , \outreg<35> , \data<9> , \data<7> , \data<8> ,
    \outreg<39> , \data<5> , \outreg<30> , \data<6> , \outreg<34> ,
    \outreg<33> , \outreg<32> , \outreg<31> , \outreg<48> , \outreg<47> ,
    \outreg<46> , \outreg<45> , \outreg<49> , \outreg<40> , \outreg<44> ,
    \outreg<43> , \outreg<42> , \outreg<41> , \D<10> , \D<11> , \D<12> ,
    \D<13> , \D<14> , \D<15> , \D<16> , \D<17> , \D<18> , \D<19> , \D<20> ,
    \D<21> , \data_in<7> , \D<22> , \D<23> , \data_in<5> , \D<24> ,
    \data_in<6> , \D<25> , \D<26> , \D<27> , \data_in<0> , \data_in<3> ,
    \data_in<4> , \data_in<1> , \data_in<2> , \data<37> , \data<38> ,
    \data<35> , \data<36> , \data<39> , \data<30> , \data<33> , \data<34> ,
    \data<31> , \data<32> , \data<47> , \data<48> , \data<45> , \data<46> ,
    \data<49> , \data<40> , \data<43> , \data<44> , \data<41> , \data<42> ,
    \data<17> , \data<18> , \data<15> , \count<0> , \data<16> , \count<3> ,
    \data<19> , \count<1> , \count<2> , \data<10> , \data<13> , \data<14> ,
    \data<11> , \data<12> , \data<27> , \data<28> , \data<25> , \data<26> ,
    \data<29> , \data<20> , \data<23> , \data<24> , \data<21> , \data<22> ,
    \C<0> , \C<1> , \C<2> , \C<3> , \C<4> , \C<5> , \C<6> , \C<7> , \C<8> ,
    \C<9> , \inreg<12> , \inreg<11> , \inreg<14> , \inreg<13> ,
    \inreg<10> , \inreg<19> , \inreg<16> , \inreg<15> , \inreg<18> ,
    \inreg<17> , \inreg<22> , \inreg<21> , \inreg<24> , \inreg<23> ,
    \inreg<20> , \inreg<29> , \inreg<26> , \inreg<25> , \outreg<9> ,
    \inreg<28> , \inreg<27> , \inreg<32> , \inreg<31> , \outreg<5> ,
    \inreg<34> , \outreg<6> , \inreg<33> , \outreg<7> , \outreg<8> ,
    \outreg<1> , \inreg<30> , \outreg<2> , \outreg<3> , \outreg<4> ,
    \inreg<39> , \inreg<36> , \outreg<0> , \inreg<35> , \inreg<38> ,
    \inreg<37> , \inreg<42> , \inreg<41> , \inreg<44> , \inreg<43> ,
    \inreg<40> , \inreg<49> , \inreg<46> , \inreg<45> , \encrypt_mode<0> ,
    \inreg<48> , \inreg<47> , \inreg<52> , \inreg<51> , \inreg<54> ,
    \inreg<53> , \inreg<50> , \inreg<55> , \data<57> , \data<58> ,
    \data<55> , \data<56> , \encrypt<0> , \data<59> , \data<50> ,
    \data<53> , \data<54> , \data<51> , \data<52> , \data<60> ;
  output \data_new<25> , \inreg_new<45> , \data_new<26> , \data_new<13> ,
    \data_new<14> , \data_new<11> , \inreg_new<49> , \data_new<12> ,
    \inreg_new<30> , \outreg_new<11> , \count_new<0> , \outreg_new<12> ,
    \data_new<10> , \outreg_new<13> , \outreg_new<14> , \inreg_new<34> ,
    \count_new<3> , \inreg_new<33> , \inreg_new<32> , \count_new<1> ,
    \data_new<19> , \inreg_new<31> , \count_new<2> , \outreg_new<10> ,
    \inreg_new<38> , \outreg_new<19> , \data_new<17> , \inreg_new<37> ,
    \data_new<18> , \inreg_new<36> , \data_new<15> , \inreg_new<35> ,
    \data_new<16> , \outreg_new<15> , \outreg_new<16> , \outreg_new<17> ,
    \inreg_new<39> , \outreg_new<18> , \outreg_new<21> , \outreg_new<22> ,
    \outreg_new<23> , \outreg_new<24> , \outreg_new<20> , \outreg_new<29> ,
    \outreg_new<25> , \outreg_new<26> , \outreg_new<27> , \outreg_new<28> ,
    \outreg_new<31> , \outreg_new<32> , \outreg_new<33> , \outreg_new<34> ,
    \outreg_new<30> , \outreg_new<39> , \outreg_new<35> , \outreg_new<36> ,
    \outreg_new<37> , \outreg_new<38> , \outreg_new<41> , \outreg_new<42> ,
    \outreg_new<43> , \outreg_new<44> , \outreg_new<40> , \outreg_new<49> ,
    \outreg_new<45> , \outreg_new<46> , \outreg_new<47> , \outreg_new<48> ,
    \C_new<23> , \C_new<24> , \C_new<21> , \C_new<22> , \C_new<20> ,
    \data_new<4> , \data_new<3> , \C_new<27> , \data_new<2> ,
    \data_new<1> , \C_new<25> , \data_new<0> , \C_new<26> , \C_new<13> ,
    \C_new<14> , \C_new<11> , \C_new<12> , \C_new<10> , \data_new<9> ,
    \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> ,
    \C_new<19> , \C_new<17> , \C_new<18> , \C_new<15> , \C_new<16> ,
    \D_new<13> , \D_new<14> , \D_new<11> , \D_new<12> , \D_new<10> ,
    \data_new<63> , \data_new<61> , \data_new<62> , \D_new<19> ,
    \data_new<60> , \D_new<17> , \D_new<18> , \D_new<15> , \D_new<16> ,
    \D_new<23> , \D_new<24> , \D_new<21> , \D_new<22> , \D_new<20> ,
    \data_new<53> , \data_new<54> , \data_new<51> , \data_new<52> ,
    \data_new<50> , \D_new<27> , \D_new<25> , \D_new<26> , \data_new<59> ,
    \data_new<57> , \data_new<58> , \data_new<55> , \data_new<56> ,
    \D_new<7> , \C_new<6> , \D_new<8> , \C_new<5> , \D_new<5> , \C_new<8> ,
    \D_new<6> , \C_new<7> , \C_new<9> , \D_new<9> , \D_new<0> , \C_new<0> ,
    \D_new<3> , \C_new<2> , \D_new<4> , \C_new<1> , \D_new<1> , \C_new<4> ,
    \D_new<2> , \C_new<3> , \inreg_new<50> , \inreg_new<9> ,
    \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<6> ,
    \inreg_new<51> , \inreg_new<5> , \inreg_new<8> , \inreg_new<7> ,
    \inreg_new<2> , \inreg_new<55> , \inreg_new<1> , \inreg_new<4> ,
    \inreg_new<3> , \inreg_new<0> , \encrypt_mode_new<0> , \outreg_new<9> ,
    \outreg_new<51> , \outreg_new<52> , \outreg_new<53> , \outreg_new<5> ,
    \outreg_new<54> , \outreg_new<6> , \outreg_new<7> , \outreg_new<8> ,
    \outreg_new<1> , \outreg_new<50> , \outreg_new<2> , \outreg_new<59> ,
    \outreg_new<3> , \outreg_new<4> , \outreg_new<55> , \data_new<43> ,
    \outreg_new<56> , \data_new<44> , \outreg_new<0> , \outreg_new<57> ,
    \data_new<41> , \outreg_new<58> , \data_new<42> , \inreg_new<20> ,
    \outreg_new<61> , \outreg_new<62> , \data_new<40> , \outreg_new<63> ,
    \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \data_new<49> ,
    \inreg_new<21> , \outreg_new<60> , \inreg_new<28> , \data_new<47> ,
    \inreg_new<27> , \data_new<48> , \inreg_new<26> , \data_new<45> ,
    \inreg_new<25> , \data_new<46> , \data_new<33> , \data_new<34> ,
    \data_new<31> , \inreg_new<29> , \data_new<32> , \inreg_new<10> ,
    \data_new<30> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> ,
    \data_new<39> , \inreg_new<11> , \inreg_new<18> , \data_new<37> ,
    \inreg_new<17> , \data_new<38> , \inreg_new<16> , \data_new<35> ,
    \inreg_new<15> , \data_new<36> , \data_new<23> , \data_new<24> ,
    \data_new<21> , \inreg_new<19> , \data_new<22> , \inreg_new<40> ,
    \data_new<20> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> ,
    \data_new<29> , \inreg_new<41> , \inreg_new<48> , \data_new<27> ,
    \inreg_new<47> , \data_new<28> , \inreg_new<46> ;
  wire n502, n503, n504, n505, n506, n508, n509, n510, n512, n513, n515,
    n516, n518, n519, n521, n522, n524, n525, n527, n528, n530, n531, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n644, n645, n647, n648, n649, n650, n652, n653, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n732, n733, n734, n735, n737, n738, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n752, n753, n755, n756, n758, n759,
    n760, n762, n763, n765, n766, n768, n769, n770, n771, n772, n773, n775,
    n776, n777, n778, n780, n781, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n862,
    n863, n865, n866, n868, n869, n871, n872, n874, n875, n877, n878, n880,
    n881, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n963, n964, n965, n966,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1088, n1089, n1091, n1092, n1093, n1094,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1236, n1237, n1238,
    n1239, n1241, n1242, n1243, n1244, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
    n1353, n1354, n1355, n1356, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1446, n1447, n1448, n1449, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1578, n1579, n1580, n1581, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1591, n1592, n1593, n1594, n1596, n1597, n1598, n1599,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1658, n1659, n1660, n1661, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1759, n1760, n1761, n1762, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1808, n1809, n1810, n1811, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1869, n1870, n1871, n1872, n1874, n1875, n1876, n1877, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1961, n1962,
    n1963, n1964, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1974,
    n1975, n1976, n1977, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2060,
    n2061, n2063, n2064, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2079, n2080, n2082, n2083, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2098, n2099, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2179, n2180, n2182, n2183, n2185,
    n2186, n2188, n2189, n2191, n2192, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2362, n2363, n2365, n2366, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2381, n2382,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2501, n2502,
    n2504, n2505, n2507, n2508, n2510, n2511, n2513, n2514, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2555, n2556, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2601, n2602,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2944, n2945,
    n2947, n2948, n2950, n2951, n2953, n2954, n2956, n2957, n2959, n2960,
    n2962, n2963, n2965, n2966, n2968, n2969, n2971, n2972, n2974, n2975,
    n2977, n2978, n2980, n2981, n2983, n2984, n2986, n2987, n2989, n2990,
    n2992, n2993, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3090, n3091, n3092, n3093, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3135, n3136,
    n3137, n3138, n3140, n3141, n3142, n3143, n3145, n3146, n3147, n3148,
    n3150, n3151, n3152, n3153, n3155, n3156, n3157, n3158, n3160, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3204, n3205, n3206, n3207, n3209, n3210, n3211, n3212, n3214,
    n3215, n3216, n3217, n3218, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3255, n3256,
    n3257, n3258, n3260, n3261, n3262, n3263, n3265, n3266, n3268, n3269,
    n3271, n3272, n3274, n3275, n3276, n3277, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3322, n3323,
    n3325, n3326, n3328, n3329, n3331, n3332, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3378,
    n3379, n3381, n3382, n3384, n3385, n3387, n3388, n3390, n3391, n3393,
    n3394, n3396, n3397, n3399, n3400, n3402, n3403, n3405, n3406, n3408,
    n3409, n3411, n3412, n3414, n3415, n3417, n3418, n3420, n3421, n3423,
    n3424, n3426, n3427, n3429, n3430, n3432, n3433, n3435, n3436, n3438,
    n3439, n3441, n3442, n3444, n3445, n3447, n3448, n3450, n3451, n3453,
    n3454, n3456, n3457, n3459, n3460, n3462, n3463, n3465, n3466, n3468,
    n3469, n3471, n3472, n3474, n3475, n3477, n3478, n3480, n3481, n3483,
    n3484, n3486, n3487, n3489, n3490, n3492, n3493, n3495, n3496, n3498,
    n3499, n3501, n3502, n3504, n3505, n3507, n3508, n3510, n3511, n3513,
    n3514, n3516, n3517, n3519, n3520, n3522, n3523, n3525, n3526, n3528,
    n3529, n3531, n3532, n3534, n3535, n3537, n3538;
  assign n502 = \count<0>  & \count<1> ;
  assign n503 = \count<2>  & n502;
  assign n504 = \count<3>  & n503;
  assign n505 = \inreg<47>  & n504;
  assign n506 = \data<57>  & ~n504;
  assign \data_new<25>  = n505 | n506;
  assign n508 = \count<0>  & ~n504;
  assign n509 = \inreg<37>  & n508;
  assign n510 = ~\count<0>  & \inreg<45> ;
  assign \inreg_new<45>  = n509 | n510;
  assign n512 = \inreg<39>  & n504;
  assign n513 = \data<58>  & ~n504;
  assign \data_new<26>  = n512 | n513;
  assign n515 = \inreg<11>  & n504;
  assign n516 = \data<45>  & ~n504;
  assign \data_new<13>  = n515 | n516;
  assign n518 = \inreg<3>  & n504;
  assign n519 = \data<46>  & ~n504;
  assign \data_new<14>  = n518 | n519;
  assign n521 = \inreg<27>  & n504;
  assign n522 = \data<43>  & ~n504;
  assign \data_new<11>  = n521 | n522;
  assign n524 = \inreg<41>  & n508;
  assign n525 = ~\count<0>  & \inreg<49> ;
  assign \inreg_new<49>  = n524 | n525;
  assign n527 = \inreg<19>  & n504;
  assign n528 = \data<44>  & ~n504;
  assign \data_new<12>  = n527 | n528;
  assign n530 = \inreg<22>  & n508;
  assign n531 = ~\count<0>  & \inreg<30> ;
  assign \inreg_new<30>  = n530 | n531;
  assign n533 = ~\D<3>  & \data<32> ;
  assign n534 = \D<3>  & ~\data<32> ;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~\D<13>  & \data<60> ;
  assign n537 = \D<13>  & ~\data<60> ;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n535 & ~n538;
  assign n540 = \data<62>  & ~\D<7> ;
  assign n541 = ~\data<62>  & \D<7> ;
  assign n542 = ~n540 & ~n541;
  assign n543 = n535 & n538;
  assign n544 = ~\D<17>  & \data<59> ;
  assign n545 = \D<17>  & ~\data<59> ;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n542 & ~n546;
  assign n548 = n543 & n547;
  assign n549 = ~n542 & n546;
  assign n550 = \data<63>  & ~\D<0> ;
  assign n551 = ~\data<63>  & \D<0> ;
  assign n552 = ~n550 & ~n551;
  assign n553 = \data<61>  & ~\D<21> ;
  assign n554 = ~\data<61>  & \D<21> ;
  assign n555 = ~n553 & ~n554;
  assign n556 = n552 & ~n555;
  assign n557 = n549 & n556;
  assign n558 = n552 & n555;
  assign n559 = ~n535 & n538;
  assign n560 = ~n552 & ~n555;
  assign n561 = ~n535 & n555;
  assign n562 = n542 & ~n546;
  assign n563 = n556 & n562;
  assign n564 = n535 & ~n538;
  assign n565 = n546 & ~n552;
  assign n566 = n538 & n561;
  assign n567 = n552 & n561;
  assign n568 = ~n542 & ~n561;
  assign n569 = ~n560 & n568;
  assign n570 = ~n559 & n569;
  assign n571 = ~n558 & n570;
  assign n572 = ~n557 & n571;
  assign n573 = ~n548 & n572;
  assign n574 = ~n543 & ~n555;
  assign n575 = n549 & n574;
  assign n576 = ~n539 & n575;
  assign n577 = n543 & n552;
  assign n578 = ~n549 & n577;
  assign n579 = ~n563 & n578;
  assign n580 = n564 & ~n565;
  assign n581 = ~n560 & n580;
  assign n582 = ~n558 & n581;
  assign n583 = n542 & ~n556;
  assign n584 = n539 & n583;
  assign n585 = n542 & n565;
  assign n586 = n566 & n585;
  assign n587 = n547 & ~n556;
  assign n588 = n559 & n587;
  assign n589 = n542 & n543;
  assign n590 = n560 & n589;
  assign n591 = n559 & n563;
  assign n592 = n549 & n567;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n590 & n593;
  assign n595 = ~n588 & n594;
  assign n596 = ~n586 & n595;
  assign n597 = ~n584 & n596;
  assign n598 = ~n582 & n597;
  assign n599 = ~n579 & n598;
  assign n600 = ~n576 & n599;
  assign n601 = ~n573 & n600;
  assign n602 = n543 & n562;
  assign n603 = ~n552 & n564;
  assign n604 = ~n538 & n565;
  assign n605 = n547 & n566;
  assign n606 = ~n535 & ~n555;
  assign n607 = n604 & n606;
  assign n608 = ~n542 & ~n601;
  assign n609 = n539 & n608;
  assign n610 = ~n562 & n564;
  assign n611 = n558 & n610;
  assign n612 = ~n535 & n601;
  assign n613 = n560 & n612;
  assign n614 = n538 & n542;
  assign n615 = n565 & n614;
  assign n616 = n538 & n546;
  assign n617 = n556 & n616;
  assign n618 = n555 & n602;
  assign n619 = n548 & ~n555;
  assign n620 = ~n538 & n563;
  assign n621 = n562 & n603;
  assign n622 = ~n542 & n604;
  assign n623 = n562 & n567;
  assign n624 = ~n605 & ~n607;
  assign n625 = ~n623 & n624;
  assign n626 = ~n622 & n625;
  assign n627 = ~n621 & n626;
  assign n628 = ~n620 & n627;
  assign n629 = ~n619 & n628;
  assign n630 = ~n618 & n629;
  assign n631 = ~n617 & n630;
  assign n632 = ~n615 & n631;
  assign n633 = ~n613 & n632;
  assign n634 = ~n611 & n633;
  assign n635 = ~n609 & n634;
  assign n636 = ~\data<14>  & ~n635;
  assign n637 = \data<14>  & n635;
  assign n638 = ~n636 & ~n637;
  assign n639 = n504 & ~n638;
  assign n640 = \outreg<19>  & n508;
  assign n641 = \outreg<11>  & ~\count<0> ;
  assign n642 = ~n640 & ~n641;
  assign \outreg_new<11>  = n639 | ~n642;
  assign n644 = \load_key<0>  & n504;
  assign n645 = ~\reset<0>  & ~n644;
  assign \count_new<0>  = ~\count<0>  & n645;
  assign n647 = \outreg<20>  & n508;
  assign n648 = \outreg<12>  & ~\count<0> ;
  assign n649 = \data<54>  & n504;
  assign n650 = ~n648 & ~n649;
  assign \outreg_new<12>  = n647 | ~n650;
  assign n652 = \inreg<35>  & n504;
  assign n653 = \data<42>  & ~n504;
  assign \data_new<10>  = n652 | n653;
  assign n655 = ~\C<23>  & \data<34> ;
  assign n656 = \C<23>  & ~\data<34> ;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~\C<16>  & \data<32> ;
  assign n659 = \C<16>  & ~\data<32> ;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n657 & ~n660;
  assign n662 = \data<36>  & ~\C<4> ;
  assign n663 = ~\data<36>  & \C<4> ;
  assign n664 = ~n662 & ~n663;
  assign n665 = \data<35>  & ~\C<0> ;
  assign n666 = ~\data<35>  & \C<0> ;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n664 & n667;
  assign n669 = n657 & n660;
  assign n670 = n664 & ~n667;
  assign n671 = ~\C<10>  & \data<33> ;
  assign n672 = \C<10>  & ~\data<33> ;
  assign n673 = ~n671 & ~n672;
  assign n674 = \data<63>  & ~\C<13> ;
  assign n675 = ~\data<63>  & \C<13> ;
  assign n676 = ~n674 & ~n675;
  assign n677 = n673 & ~n676;
  assign n678 = n657 & ~n660;
  assign n679 = ~n673 & n676;
  assign n680 = ~n664 & ~n667;
  assign n681 = n673 & n676;
  assign n682 = ~n657 & n660;
  assign n683 = n661 & n670;
  assign n684 = ~n673 & ~n676;
  assign n685 = n682 & n684;
  assign n686 = ~n673 & n682;
  assign n687 = n664 & n667;
  assign n688 = n673 & n680;
  assign n689 = ~n670 & n677;
  assign n690 = ~n669 & n689;
  assign n691 = ~n668 & n690;
  assign n692 = ~n661 & n691;
  assign n693 = ~n677 & ~n680;
  assign n694 = ~n679 & n693;
  assign n695 = n678 & n694;
  assign n696 = n681 & ~n682;
  assign n697 = ~n670 & n696;
  assign n698 = ~n668 & n697;
  assign n699 = ~n681 & ~n684;
  assign n700 = n683 & n699;
  assign n701 = n668 & ~n681;
  assign n702 = n661 & n701;
  assign n703 = n669 & n670;
  assign n704 = n684 & n703;
  assign n705 = n669 & n677;
  assign n706 = n668 & n705;
  assign n707 = n681 & n682;
  assign n708 = n668 & n707;
  assign n709 = ~n667 & n685;
  assign n710 = n686 & n687;
  assign n711 = n661 & n688;
  assign n712 = n669 & n679;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n710 & n713;
  assign n715 = ~n709 & n714;
  assign n716 = ~n708 & n715;
  assign n717 = ~n706 & n716;
  assign n718 = ~n704 & n717;
  assign n719 = ~n702 & n718;
  assign n720 = ~n700 & n719;
  assign n721 = ~n698 & n720;
  assign n722 = ~n695 & n721;
  assign n723 = ~n692 & n722;
  assign n724 = ~\data<22>  & ~n723;
  assign n725 = \data<22>  & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = n504 & ~n726;
  assign n728 = \outreg<21>  & n508;
  assign n729 = \outreg<13>  & ~\count<0> ;
  assign n730 = ~n728 & ~n729;
  assign \outreg_new<13>  = n727 | ~n730;
  assign n732 = \outreg<22>  & n508;
  assign n733 = \outreg<14>  & ~\count<0> ;
  assign n734 = \data<62>  & n504;
  assign n735 = ~n733 & ~n734;
  assign \outreg_new<14>  = n732 | ~n735;
  assign n737 = \inreg<26>  & n508;
  assign n738 = ~\count<0>  & \inreg<34> ;
  assign \inreg_new<34>  = n737 | n738;
  assign n740 = ~\count<0>  & ~\count<3> ;
  assign n741 = \count<1>  & \count<2> ;
  assign n742 = ~n740 & n741;
  assign n743 = ~\count<1>  & ~\count<2> ;
  assign n744 = n740 & n743;
  assign n745 = ~n742 & ~n744;
  assign n746 = \count<1>  & ~n504;
  assign n747 = ~n745 & n746;
  assign n748 = n645 & n747;
  assign n749 = \count<3>  & n745;
  assign n750 = n645 & n749;
  assign \count_new<3>  = n748 | n750;
  assign n752 = \inreg<25>  & n508;
  assign n753 = ~\count<0>  & \inreg<33> ;
  assign \inreg_new<33>  = n752 | n753;
  assign n755 = \inreg<24>  & n508;
  assign n756 = ~\count<0>  & \inreg<32> ;
  assign \inreg_new<32>  = n755 | n756;
  assign n758 = \count<1>  & \count_new<0> ;
  assign n759 = ~\count<1>  & ~\count_new<0> ;
  assign n760 = n645 & n759;
  assign \count_new<1>  = n758 | n760;
  assign n762 = \inreg<29>  & n504;
  assign n763 = \data<51>  & ~n504;
  assign \data_new<19>  = n762 | n763;
  assign n765 = \inreg<23>  & n508;
  assign n766 = ~\count<0>  & \inreg<31> ;
  assign \inreg_new<31>  = n765 | n766;
  assign n768 = \count<1>  & ~\count<2> ;
  assign n769 = ~\count_new<0>  & n768;
  assign n770 = n645 & n769;
  assign n771 = \count<2>  & \count_new<1> ;
  assign n772 = \count<2>  & \count_new<0> ;
  assign n773 = ~n771 & ~n772;
  assign \count_new<2>  = n770 | ~n773;
  assign n775 = \outreg<18>  & n508;
  assign n776 = \outreg<10>  & ~\count<0> ;
  assign n777 = \data<46>  & n504;
  assign n778 = ~n776 & ~n777;
  assign \outreg_new<10>  = n775 | ~n778;
  assign n780 = \inreg<30>  & n508;
  assign n781 = ~\count<0>  & \inreg<38> ;
  assign \inreg_new<38>  = n780 | n781;
  assign n783 = ~\D<2>  & \data<49> ;
  assign n784 = \D<2>  & ~\data<49> ;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~\D<23>  & \data<48> ;
  assign n787 = \D<23>  & ~\data<48> ;
  assign n788 = ~n786 & ~n787;
  assign n789 = n785 & n788;
  assign n790 = ~\D<26>  & \data<52> ;
  assign n791 = \D<26>  & ~\data<52> ;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~\D<8>  & \data<50> ;
  assign n794 = \D<8>  & ~\data<50> ;
  assign n795 = ~n793 & ~n794;
  assign n796 = n792 & n795;
  assign n797 = ~n792 & ~n795;
  assign n798 = ~\D<18>  & \data<51> ;
  assign n799 = \D<18>  & ~\data<51> ;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~\D<12>  & \data<47> ;
  assign n802 = \D<12>  & ~\data<47> ;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n800 & ~n803;
  assign n805 = ~n785 & n788;
  assign n806 = ~n785 & ~n788;
  assign n807 = n785 & ~n788;
  assign n808 = n800 & n803;
  assign n809 = n800 & ~n803;
  assign n810 = ~n792 & n795;
  assign n811 = ~n800 & n803;
  assign n812 = ~n809 & ~n811;
  assign n813 = ~n789 & ~n806;
  assign n814 = n792 & ~n795;
  assign n815 = n804 & ~n805;
  assign n816 = ~n797 & n815;
  assign n817 = ~n796 & n816;
  assign n818 = ~n789 & n817;
  assign n819 = n797 & n804;
  assign n820 = ~n807 & n819;
  assign n821 = ~n806 & n820;
  assign n822 = ~n797 & n808;
  assign n823 = ~n796 & n822;
  assign n824 = n789 & n823;
  assign n825 = n796 & n809;
  assign n826 = n806 & n825;
  assign n827 = n792 & n808;
  assign n828 = n806 & n827;
  assign n829 = n809 & n810;
  assign n830 = n807 & n829;
  assign n831 = n805 & n812;
  assign n832 = n796 & n831;
  assign n833 = n785 & ~n812;
  assign n834 = n796 & n833;
  assign n835 = ~n812 & ~n813;
  assign n836 = n797 & n835;
  assign n837 = ~n800 & n805;
  assign n838 = n810 & n837;
  assign n839 = ~n812 & n813;
  assign n840 = n814 & n839;
  assign n841 = ~n792 & n813;
  assign n842 = n808 & n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = ~n838 & n843;
  assign n845 = ~n836 & n844;
  assign n846 = ~n834 & n845;
  assign n847 = ~n832 & n846;
  assign n848 = ~n830 & n847;
  assign n849 = ~n828 & n848;
  assign n850 = ~n826 & n849;
  assign n851 = ~n824 & n850;
  assign n852 = ~n821 & n851;
  assign n853 = ~n818 & n852;
  assign n854 = ~\data<13>  & ~n853;
  assign n855 = \data<13>  & n853;
  assign n856 = ~n854 & ~n855;
  assign n857 = n504 & ~n856;
  assign n858 = \outreg<27>  & n508;
  assign n859 = \outreg<19>  & ~\count<0> ;
  assign n860 = ~n858 & ~n859;
  assign \outreg_new<19>  = n857 | ~n860;
  assign n862 = \inreg<45>  & n504;
  assign n863 = \data<49>  & ~n504;
  assign \data_new<17>  = n862 | n863;
  assign n865 = \inreg<29>  & n508;
  assign n866 = ~\count<0>  & \inreg<37> ;
  assign \inreg_new<37>  = n865 | n866;
  assign n868 = \inreg<37>  & n504;
  assign n869 = \data<50>  & ~n504;
  assign \data_new<18>  = n868 | n869;
  assign n871 = \inreg<28>  & n508;
  assign n872 = ~\count<0>  & \inreg<36> ;
  assign \inreg_new<36>  = n871 | n872;
  assign n874 = \data_in<3>  & n504;
  assign n875 = \data<47>  & ~n504;
  assign \data_new<15>  = n874 | n875;
  assign n877 = \inreg<27>  & n508;
  assign n878 = ~\count<0>  & \inreg<35> ;
  assign \inreg_new<35>  = n877 | n878;
  assign n880 = \inreg<53>  & n504;
  assign n881 = \data<48>  & ~n504;
  assign \data_new<16>  = n880 | n881;
  assign n883 = n661 & n680;
  assign n884 = n660 & ~n677;
  assign n885 = n687 & n884;
  assign n886 = ~n679 & n885;
  assign n887 = ~n685 & n886;
  assign n888 = n670 & ~n681;
  assign n889 = ~n669 & n888;
  assign n890 = ~n661 & n889;
  assign n891 = n660 & ~n680;
  assign n892 = ~n687 & n891;
  assign n893 = n679 & n892;
  assign n894 = ~n660 & ~n680;
  assign n895 = n681 & n894;
  assign n896 = ~n687 & n895;
  assign n897 = n679 & n687;
  assign n898 = n686 & n897;
  assign n899 = ~n668 & n677;
  assign n900 = n678 & n899;
  assign n901 = n668 & ~n673;
  assign n902 = n678 & n901;
  assign n903 = n669 & n680;
  assign n904 = ~n679 & n903;
  assign n905 = n660 & n677;
  assign n906 = n668 & n905;
  assign n907 = ~n657 & n677;
  assign n908 = n687 & n907;
  assign n909 = ~n883 & ~n908;
  assign n910 = ~n906 & n909;
  assign n911 = ~n904 & n910;
  assign n912 = ~n902 & n911;
  assign n913 = ~n900 & n912;
  assign n914 = ~n898 & n913;
  assign n915 = ~n896 & n914;
  assign n916 = ~n893 & n915;
  assign n917 = ~n890 & n916;
  assign n918 = ~n887 & n917;
  assign n919 = n676 & n918;
  assign n920 = ~n657 & n919;
  assign n921 = ~n680 & n920;
  assign n922 = ~n687 & n921;
  assign n923 = ~n660 & ~n664;
  assign n924 = n677 & n923;
  assign n925 = ~n883 & n924;
  assign n926 = n680 & ~n918;
  assign n927 = ~n677 & n926;
  assign n928 = ~n679 & n927;
  assign n929 = ~n676 & ~n918;
  assign n930 = n667 & n929;
  assign n931 = n669 & n930;
  assign n932 = n670 & n684;
  assign n933 = n686 & n932;
  assign n934 = n679 & n703;
  assign n935 = ~n660 & ~n676;
  assign n936 = n687 & n935;
  assign n937 = n677 & n918;
  assign n938 = n670 & n937;
  assign n939 = n667 & n676;
  assign n940 = n682 & n939;
  assign n941 = ~n664 & n686;
  assign n942 = n678 & n679;
  assign n943 = n678 & n687;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n941 & n944;
  assign n946 = ~n940 & n945;
  assign n947 = ~n938 & n946;
  assign n948 = ~n936 & n947;
  assign n949 = ~n934 & n948;
  assign n950 = ~n933 & n949;
  assign n951 = ~n931 & n950;
  assign n952 = ~n928 & n951;
  assign n953 = ~n925 & n952;
  assign n954 = ~n922 & n953;
  assign n955 = ~\data<30>  & ~n954;
  assign n956 = \data<30>  & n954;
  assign n957 = ~n955 & ~n956;
  assign n958 = n504 & ~n957;
  assign n959 = \outreg<23>  & n508;
  assign n960 = \outreg<15>  & ~\count<0> ;
  assign n961 = ~n959 & ~n960;
  assign \outreg_new<15>  = n958 | ~n961;
  assign n963 = \outreg<24>  & n508;
  assign n964 = \outreg<16>  & ~\count<0> ;
  assign n965 = \data<37>  & n504;
  assign n966 = ~n964 & ~n965;
  assign \outreg_new<16>  = n963 | ~n966;
  assign n968 = \data<42>  & ~\C<3> ;
  assign n969 = ~\data<42>  & \C<3> ;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~\C<18>  & \data<40> ;
  assign n972 = \C<18>  & ~\data<40> ;
  assign n973 = ~n971 & ~n972;
  assign n974 = n970 & ~n973;
  assign n975 = ~\C<11>  & \data<41> ;
  assign n976 = \C<11>  & ~\data<41> ;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n973 & n977;
  assign n979 = n973 & ~n977;
  assign n980 = ~n978 & ~n979;
  assign n981 = \data<44>  & ~\C<7> ;
  assign n982 = ~\data<44>  & \C<7> ;
  assign n983 = ~n981 & ~n982;
  assign n984 = ~\C<25>  & \data<43> ;
  assign n985 = \C<25>  & ~\data<43> ;
  assign n986 = ~n984 & ~n985;
  assign n987 = n977 & n986;
  assign n988 = ~\C<22>  & \data<39> ;
  assign n989 = \C<22>  & ~\data<39> ;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n983 & ~n990;
  assign n992 = n987 & n991;
  assign n993 = n974 & ~n986;
  assign n994 = ~n970 & ~n986;
  assign n995 = n970 & n973;
  assign n996 = n977 & n994;
  assign n997 = n986 & n995;
  assign n998 = ~n996 & ~n997;
  assign n999 = n983 & n990;
  assign n1000 = ~n973 & ~n977;
  assign n1001 = ~n977 & n986;
  assign n1002 = n983 & ~n990;
  assign n1003 = ~n983 & n990;
  assign n1004 = ~n986 & n995;
  assign n1005 = ~n970 & ~n973;
  assign n1006 = n1002 & n1004;
  assign n1007 = n977 & n991;
  assign n1008 = n993 & n1007;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = n970 & n977;
  assign n1011 = ~n999 & n1010;
  assign n1012 = n998 & n1011;
  assign n1013 = ~n993 & n1012;
  assign n1014 = ~n992 & n1013;
  assign n1015 = ~n1002 & ~n1003;
  assign n1016 = n1001 & n1015;
  assign n1017 = n1000 & n1016;
  assign n1018 = n993 & n1003;
  assign n1019 = n1000 & n1018;
  assign n1020 = ~n986 & n1002;
  assign n1021 = n1000 & n1020;
  assign n1022 = ~n980 & n983;
  assign n1023 = n1004 & n1022;
  assign n1024 = ~n983 & n1001;
  assign n1025 = ~n998 & n1024;
  assign n1026 = ~n990 & n1005;
  assign n1027 = n987 & n1026;
  assign n1028 = ~n980 & ~n983;
  assign n1029 = n994 & n1028;
  assign n1030 = ~n970 & ~n991;
  assign n1031 = n1001 & n1030;
  assign n1032 = ~n998 & n999;
  assign n1033 = n1009 & ~n1032;
  assign n1034 = ~n1031 & n1033;
  assign n1035 = ~n1029 & n1034;
  assign n1036 = ~n1027 & n1035;
  assign n1037 = ~n1025 & n1036;
  assign n1038 = ~n1023 & n1037;
  assign n1039 = ~n1021 & n1038;
  assign n1040 = ~n1019 & n1039;
  assign n1041 = ~n1017 & n1040;
  assign n1042 = ~n1014 & n1041;
  assign n1043 = ~n970 & n973;
  assign n1044 = n992 & n1043;
  assign n1045 = ~n983 & ~n1042;
  assign n1046 = n980 & n1045;
  assign n1047 = n974 & n1046;
  assign n1048 = ~n990 & n1042;
  assign n1049 = ~n986 & n1048;
  assign n1050 = n974 & n1049;
  assign n1051 = n980 & ~n991;
  assign n1052 = n994 & n1051;
  assign n1053 = ~n999 & n1052;
  assign n1054 = ~n980 & ~n986;
  assign n1055 = ~n1003 & n1054;
  assign n1056 = ~n1002 & n1055;
  assign n1057 = ~n977 & ~n1042;
  assign n1058 = ~n980 & n1057;
  assign n1059 = n1002 & n1058;
  assign n1060 = n986 & n999;
  assign n1061 = n1043 & n1060;
  assign n1062 = n995 & ~n999;
  assign n1063 = n987 & n1062;
  assign n1064 = n986 & n1003;
  assign n1065 = n1005 & n1064;
  assign n1066 = n983 & n986;
  assign n1067 = n974 & n1066;
  assign n1068 = n995 & ~n1042;
  assign n1069 = n1003 & n1068;
  assign n1070 = ~n1044 & ~n1069;
  assign n1071 = ~n1067 & n1070;
  assign n1072 = ~n1065 & n1071;
  assign n1073 = ~n1063 & n1072;
  assign n1074 = ~n1061 & n1073;
  assign n1075 = ~n1059 & n1074;
  assign n1076 = ~n1056 & n1075;
  assign n1077 = ~n1053 & n1076;
  assign n1078 = ~n1050 & n1077;
  assign n1079 = ~n1047 & n1078;
  assign n1080 = ~\data<5>  & ~n1079;
  assign n1081 = \data<5>  & n1079;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n504 & ~n1082;
  assign n1084 = \outreg<25>  & n508;
  assign n1085 = \outreg<17>  & ~\count<0> ;
  assign n1086 = ~n1084 & ~n1085;
  assign \outreg_new<17>  = n1083 | ~n1086;
  assign n1088 = \inreg<31>  & n508;
  assign n1089 = ~\count<0>  & \inreg<39> ;
  assign \inreg_new<39>  = n1088 | n1089;
  assign n1091 = \outreg<26>  & n508;
  assign n1092 = \outreg<18>  & ~\count<0> ;
  assign n1093 = \data<45>  & n504;
  assign n1094 = ~n1092 & ~n1093;
  assign \outreg_new<18>  = n1091 | ~n1094;
  assign n1096 = ~\D<24>  & \data<60> ;
  assign n1097 = \D<24>  & ~\data<60> ;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~\D<27>  & \data<58> ;
  assign n1100 = \D<27>  & ~\data<58> ;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = ~\D<20>  & \data<56> ;
  assign n1103 = \D<20>  & ~\data<56> ;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~\D<10>  & \data<57> ;
  assign n1106 = \D<10>  & ~\data<57> ;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = n1104 & ~n1107;
  assign n1109 = ~\D<5>  & \data<59> ;
  assign n1110 = \D<5>  & ~\data<59> ;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n1101 & ~n1111;
  assign n1113 = n1098 & n1112;
  assign n1114 = ~n1098 & n1111;
  assign n1115 = n1104 & n1107;
  assign n1116 = ~n1098 & ~n1111;
  assign n1117 = n1108 & n1116;
  assign n1118 = ~n1104 & n1113;
  assign n1119 = n1114 & n1115;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~n1117 & n1120;
  assign n1122 = n1098 & n1111;
  assign n1123 = ~\D<15>  & \data<55> ;
  assign n1124 = \D<15>  & ~\data<55> ;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = n1101 & ~n1125;
  assign n1127 = ~n1098 & ~n1104;
  assign n1128 = n1115 & n1125;
  assign n1129 = n1111 & n1125;
  assign n1130 = n1107 & n1127;
  assign n1131 = ~n1107 & n1125;
  assign n1132 = n1108 & n1122;
  assign n1133 = ~n1101 & ~n1111;
  assign n1134 = n1098 & n1133;
  assign n1135 = ~n1104 & n1107;
  assign n1136 = ~n1101 & ~n1125;
  assign n1137 = n1122 & n1136;
  assign n1138 = n1107 & n1125;
  assign n1139 = ~n1112 & n1138;
  assign n1140 = ~n1122 & n1139;
  assign n1141 = n1121 & n1140;
  assign n1142 = ~n1107 & ~n1111;
  assign n1143 = n1127 & n1142;
  assign n1144 = ~n1126 & n1143;
  assign n1145 = ~n1107 & n1111;
  assign n1146 = n1127 & n1145;
  assign n1147 = n1126 & n1146;
  assign n1148 = n1107 & n1113;
  assign n1149 = ~n1128 & n1148;
  assign n1150 = n1101 & n1104;
  assign n1151 = n1129 & n1150;
  assign n1152 = ~n1111 & ~n1125;
  assign n1153 = n1130 & n1152;
  assign n1154 = ~n1104 & n1122;
  assign n1155 = n1131 & n1154;
  assign n1156 = ~n1125 & n1132;
  assign n1157 = n1104 & n1134;
  assign n1158 = n1135 & n1137;
  assign n1159 = ~n1121 & ~n1125;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1157 & n1160;
  assign n1162 = ~n1156 & n1161;
  assign n1163 = ~n1155 & n1162;
  assign n1164 = ~n1153 & n1163;
  assign n1165 = ~n1151 & n1164;
  assign n1166 = ~n1149 & n1165;
  assign n1167 = ~n1147 & n1166;
  assign n1168 = ~n1144 & n1167;
  assign n1169 = ~n1141 & n1168;
  assign n1170 = n1112 & n1131;
  assign n1171 = ~n1111 & n1136;
  assign n1172 = n1098 & n1171;
  assign n1173 = n1114 & n1136;
  assign n1174 = n1113 & n1128;
  assign n1175 = n1113 & ~n1125;
  assign n1176 = n1135 & n1175;
  assign n1177 = ~n1174 & ~n1176;
  assign n1178 = ~n1098 & n1108;
  assign n1179 = n1171 & n1178;
  assign n1180 = ~n1104 & ~n1169;
  assign n1181 = ~n1101 & n1180;
  assign n1182 = n1098 & n1181;
  assign n1183 = n1101 & n1125;
  assign n1184 = n1132 & n1183;
  assign n1185 = n1114 & ~n1169;
  assign n1186 = n1126 & n1185;
  assign n1187 = n1101 & n1122;
  assign n1188 = n1135 & n1187;
  assign n1189 = n1136 & ~n1169;
  assign n1190 = n1135 & n1189;
  assign n1191 = ~n1098 & n1133;
  assign n1192 = n1131 & n1191;
  assign n1193 = n1127 & n1183;
  assign n1194 = ~n1125 & n1169;
  assign n1195 = n1112 & n1194;
  assign n1196 = ~n1101 & n1128;
  assign n1197 = ~n1104 & n1170;
  assign n1198 = ~n1107 & n1172;
  assign n1199 = ~n1107 & n1173;
  assign n1200 = n1104 & n1137;
  assign n1201 = n1177 & ~n1179;
  assign n1202 = ~n1200 & n1201;
  assign n1203 = ~n1199 & n1202;
  assign n1204 = ~n1198 & n1203;
  assign n1205 = ~n1197 & n1204;
  assign n1206 = ~n1196 & n1205;
  assign n1207 = ~n1195 & n1206;
  assign n1208 = ~n1193 & n1207;
  assign n1209 = ~n1192 & n1208;
  assign n1210 = ~n1190 & n1209;
  assign n1211 = ~n1188 & n1210;
  assign n1212 = ~n1186 & n1211;
  assign n1213 = ~n1184 & n1212;
  assign n1214 = ~n1182 & n1213;
  assign n1215 = ~\data<21>  & ~n1214;
  assign n1216 = \data<21>  & n1214;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = n504 & ~n1217;
  assign n1219 = \outreg<29>  & n508;
  assign n1220 = \outreg<21>  & ~\count<0> ;
  assign n1221 = ~n1219 & ~n1220;
  assign \outreg_new<21>  = n1218 | ~n1221;
  assign n1223 = \outreg<30>  & n508;
  assign n1224 = \outreg<22>  & ~\count<0> ;
  assign n1225 = \data<61>  & n504;
  assign n1226 = ~n1224 & ~n1225;
  assign \outreg_new<22>  = n1223 | ~n1226;
  assign n1228 = ~\data<29>  & ~n1042;
  assign n1229 = \data<29>  & n1042;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = n504 & ~n1230;
  assign n1232 = \outreg<31>  & n508;
  assign n1233 = \outreg<23>  & ~\count<0> ;
  assign n1234 = ~n1232 & ~n1233;
  assign \outreg_new<23>  = n1231 | ~n1234;
  assign n1236 = \outreg<32>  & n508;
  assign n1237 = \outreg<24>  & ~\count<0> ;
  assign n1238 = \data<36>  & n504;
  assign n1239 = ~n1237 & ~n1238;
  assign \outreg_new<24>  = n1236 | ~n1239;
  assign n1241 = \outreg<28>  & n508;
  assign n1242 = \outreg<20>  & ~\count<0> ;
  assign n1243 = \data<53>  & n504;
  assign n1244 = ~n1242 & ~n1243;
  assign \outreg_new<20>  = n1241 | ~n1244;
  assign n1246 = n547 & n560;
  assign n1247 = n564 & ~n601;
  assign n1248 = ~n562 & n1247;
  assign n1249 = ~n549 & n1248;
  assign n1250 = ~n538 & n601;
  assign n1251 = n555 & n1250;
  assign n1252 = n549 & n1251;
  assign n1253 = ~n555 & ~n601;
  assign n1254 = n535 & n1253;
  assign n1255 = n565 & n1254;
  assign n1256 = n538 & n601;
  assign n1257 = ~n555 & n1256;
  assign n1258 = n565 & n1257;
  assign n1259 = n538 & n555;
  assign n1260 = ~n552 & n1259;
  assign n1261 = ~n565 & n1260;
  assign n1262 = n538 & ~n601;
  assign n1263 = n555 & n1262;
  assign n1264 = n542 & n1263;
  assign n1265 = n542 & n555;
  assign n1266 = n604 & n1265;
  assign n1267 = n567 & n616;
  assign n1268 = ~n538 & ~n546;
  assign n1269 = n567 & n1268;
  assign n1270 = ~n538 & ~n555;
  assign n1271 = n562 & n1270;
  assign n1272 = n535 & n601;
  assign n1273 = n556 & n1272;
  assign n1274 = ~n535 & n557;
  assign n1275 = ~n535 & n1246;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = ~n1273 & n1276;
  assign n1278 = ~n1271 & n1277;
  assign n1279 = ~n1269 & n1278;
  assign n1280 = ~n1267 & n1279;
  assign n1281 = ~n1266 & n1280;
  assign n1282 = ~n1264 & n1281;
  assign n1283 = ~n1261 & n1282;
  assign n1284 = ~n1258 & n1283;
  assign n1285 = ~n1255 & n1284;
  assign n1286 = ~n1252 & n1285;
  assign n1287 = ~n1249 & n1286;
  assign n1288 = ~\data<20>  & ~n1287;
  assign n1289 = \data<20>  & n1287;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = n504 & ~n1290;
  assign n1292 = \outreg<37>  & n508;
  assign n1293 = \outreg<29>  & ~\count<0> ;
  assign n1294 = ~n1292 & ~n1293;
  assign \outreg_new<29>  = n1291 | ~n1294;
  assign n1296 = n557 & n559;
  assign n1297 = n546 & ~n560;
  assign n1298 = n559 & n1297;
  assign n1299 = ~n558 & n1298;
  assign n1300 = ~n557 & n1299;
  assign n1301 = n535 & ~n546;
  assign n1302 = ~n547 & n1301;
  assign n1303 = ~n558 & n1302;
  assign n1304 = ~n603 & n1303;
  assign n1305 = ~n564 & n585;
  assign n1306 = n560 & n1305;
  assign n1307 = ~n559 & n1306;
  assign n1308 = ~n538 & ~n560;
  assign n1309 = n549 & n1308;
  assign n1310 = ~n558 & n1309;
  assign n1311 = n535 & n546;
  assign n1312 = ~n549 & n1311;
  assign n1313 = n558 & n1312;
  assign n1314 = n538 & ~n1296;
  assign n1315 = n552 & n1314;
  assign n1316 = n549 & n1315;
  assign n1317 = ~n538 & ~n552;
  assign n1318 = n547 & n1317;
  assign n1319 = ~n561 & n1318;
  assign n1320 = ~n538 & n542;
  assign n1321 = ~n565 & n1320;
  assign n1322 = n561 & n1321;
  assign n1323 = n555 & n604;
  assign n1324 = n603 & n1323;
  assign n1325 = ~n538 & n547;
  assign n1326 = n558 & n1325;
  assign n1327 = ~n546 & n560;
  assign n1328 = n559 & n1327;
  assign n1329 = n547 & n552;
  assign n1330 = n559 & n1329;
  assign n1331 = n547 & n556;
  assign n1332 = n543 & n1331;
  assign n1333 = ~n1330 & ~n1332;
  assign n1334 = ~n1328 & n1333;
  assign n1335 = ~n1326 & n1334;
  assign n1336 = ~n1324 & n1335;
  assign n1337 = ~n1322 & n1336;
  assign n1338 = ~n1319 & n1337;
  assign n1339 = ~n1316 & n1338;
  assign n1340 = ~n1313 & n1339;
  assign n1341 = ~n1310 & n1340;
  assign n1342 = ~n1307 & n1341;
  assign n1343 = ~n1304 & n1342;
  assign n1344 = ~n1300 & n1343;
  assign n1345 = ~\data<4>  & ~n1344;
  assign n1346 = \data<4>  & n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = n504 & ~n1347;
  assign n1349 = \outreg<33>  & n508;
  assign n1350 = \outreg<25>  & ~\count<0> ;
  assign n1351 = ~n1349 & ~n1350;
  assign \outreg_new<25>  = n1348 | ~n1351;
  assign n1353 = \outreg<34>  & n508;
  assign n1354 = \outreg<26>  & ~\count<0> ;
  assign n1355 = \data<44>  & n504;
  assign n1356 = ~n1354 & ~n1355;
  assign \outreg_new<26>  = n1353 | ~n1356;
  assign n1358 = \data<40>  & ~\C<9> ;
  assign n1359 = ~\data<40>  & \C<9> ;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~\C<20>  & \data<39> ;
  assign n1362 = \C<20>  & ~\data<39> ;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1360 & ~n1363;
  assign n1365 = ~\C<14>  & \data<37> ;
  assign n1366 = \C<14>  & ~\data<37> ;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n1364 & ~n1367;
  assign n1369 = \data<35>  & ~\C<2> ;
  assign n1370 = ~\data<35>  & \C<2> ;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1363 & n1371;
  assign n1373 = n1363 & n1371;
  assign n1374 = ~n1367 & n1373;
  assign n1375 = n1367 & ~n1371;
  assign n1376 = n1363 & n1375;
  assign n1377 = \data<38>  & ~\C<5> ;
  assign n1378 = ~\data<38>  & \C<5> ;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = ~\C<27>  & \data<36> ;
  assign n1381 = \C<27>  & ~\data<36> ;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = ~n1379 & ~n1382;
  assign n1384 = ~n1363 & ~n1371;
  assign n1385 = ~n1379 & n1382;
  assign n1386 = n1360 & n1385;
  assign n1387 = n1376 & n1386;
  assign n1388 = ~n1360 & n1379;
  assign n1389 = ~n1382 & n1388;
  assign n1390 = n1363 & ~n1371;
  assign n1391 = ~n1360 & ~n1367;
  assign n1392 = n1383 & n1391;
  assign n1393 = n1379 & n1382;
  assign n1394 = n1371 & n1393;
  assign n1395 = n1368 & n1394;
  assign n1396 = n1360 & ~n1383;
  assign n1397 = ~n1376 & n1396;
  assign n1398 = ~n1374 & n1397;
  assign n1399 = ~n1372 & n1398;
  assign n1400 = ~n1368 & n1399;
  assign n1401 = n1360 & ~n1387;
  assign n1402 = n1367 & n1401;
  assign n1403 = ~n1379 & n1402;
  assign n1404 = ~n1373 & n1403;
  assign n1405 = ~n1384 & n1404;
  assign n1406 = ~n1385 & n1391;
  assign n1407 = ~n1390 & n1406;
  assign n1408 = ~n1372 & n1407;
  assign n1409 = ~n1389 & n1408;
  assign n1410 = ~n1360 & ~n1363;
  assign n1411 = n1367 & n1410;
  assign n1412 = ~n1385 & n1411;
  assign n1413 = ~n1389 & n1412;
  assign n1414 = n1360 & ~n1382;
  assign n1415 = ~n1383 & n1414;
  assign n1416 = n1374 & n1415;
  assign n1417 = n1372 & n1391;
  assign n1418 = n1389 & n1417;
  assign n1419 = n1363 & n1367;
  assign n1420 = n1389 & n1419;
  assign n1421 = n1371 & n1385;
  assign n1422 = n1391 & n1421;
  assign n1423 = ~n1360 & n1382;
  assign n1424 = n1376 & n1423;
  assign n1425 = n1368 & n1383;
  assign n1426 = n1390 & n1392;
  assign n1427 = ~n1395 & ~n1426;
  assign n1428 = ~n1425 & n1427;
  assign n1429 = ~n1424 & n1428;
  assign n1430 = ~n1422 & n1429;
  assign n1431 = ~n1420 & n1430;
  assign n1432 = ~n1418 & n1431;
  assign n1433 = ~n1416 & n1432;
  assign n1434 = ~n1413 & n1433;
  assign n1435 = ~n1409 & n1434;
  assign n1436 = ~n1405 & n1435;
  assign n1437 = ~n1400 & n1436;
  assign n1438 = ~\data<12>  & ~n1437;
  assign n1439 = \data<12>  & n1437;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = n504 & ~n1440;
  assign n1442 = \outreg<35>  & n508;
  assign n1443 = \outreg<27>  & ~\count<0> ;
  assign n1444 = ~n1442 & ~n1443;
  assign \outreg_new<27>  = n1441 | ~n1444;
  assign n1446 = \outreg<36>  & n508;
  assign n1447 = \outreg<28>  & ~\count<0> ;
  assign n1448 = \data<52>  & n504;
  assign n1449 = ~n1447 & ~n1448;
  assign \outreg_new<28>  = n1446 | ~n1449;
  assign n1451 = ~\D<22>  & \data<53> ;
  assign n1452 = \D<22>  & ~\data<53> ;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~\D<1>  & \data<51> ;
  assign n1455 = \D<1>  & ~\data<51> ;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1453 & n1456;
  assign n1458 = ~\D<11>  & \data<52> ;
  assign n1459 = \D<11>  & ~\data<52> ;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = n1457 & ~n1460;
  assign n1462 = ~n1453 & ~n1456;
  assign n1463 = ~\D<4>  & \data<55> ;
  assign n1464 = \D<4>  & ~\data<55> ;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~\D<16>  & \data<54> ;
  assign n1467 = \D<16>  & ~\data<54> ;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = n1465 & ~n1468;
  assign n1470 = ~n1465 & n1468;
  assign n1471 = n1453 & n1456;
  assign n1472 = ~n1456 & ~n1460;
  assign n1473 = ~\D<19>  & \data<56> ;
  assign n1474 = \D<19>  & ~\data<56> ;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n1472 & ~n1475;
  assign n1477 = n1453 & n1476;
  assign n1478 = ~n1465 & ~n1468;
  assign n1479 = n1470 & n1475;
  assign n1480 = n1460 & ~n1475;
  assign n1481 = n1475 & n1478;
  assign n1482 = ~n1460 & ~n1475;
  assign n1483 = n1465 & n1475;
  assign n1484 = ~n1453 & n1480;
  assign n1485 = n1460 & n1481;
  assign n1486 = n1468 & n1483;
  assign n1487 = n1453 & ~n1456;
  assign n1488 = n1460 & n1487;
  assign n1489 = n1479 & n1488;
  assign n1490 = ~n1456 & ~n1475;
  assign n1491 = n1478 & n1490;
  assign n1492 = ~n1477 & n1491;
  assign n1493 = ~n1460 & n1471;
  assign n1494 = n1479 & n1493;
  assign n1495 = n1465 & n1480;
  assign n1496 = n1462 & n1495;
  assign n1497 = n1453 & n1472;
  assign n1498 = n1481 & n1497;
  assign n1499 = ~n1468 & n1471;
  assign n1500 = n1482 & n1499;
  assign n1501 = n1453 & n1460;
  assign n1502 = n1483 & n1501;
  assign n1503 = n1468 & n1471;
  assign n1504 = n1480 & n1503;
  assign n1505 = n1457 & ~n1475;
  assign n1506 = n1470 & n1505;
  assign n1507 = n1469 & n1484;
  assign n1508 = n1456 & n1485;
  assign n1509 = n1461 & n1478;
  assign n1510 = n1462 & n1479;
  assign n1511 = n1457 & n1486;
  assign n1512 = n1462 & n1469;
  assign n1513 = n1468 & n1477;
  assign n1514 = ~n1489 & ~n1513;
  assign n1515 = ~n1512 & n1514;
  assign n1516 = ~n1511 & n1515;
  assign n1517 = ~n1510 & n1516;
  assign n1518 = ~n1509 & n1517;
  assign n1519 = ~n1508 & n1518;
  assign n1520 = ~n1507 & n1519;
  assign n1521 = ~n1506 & n1520;
  assign n1522 = ~n1504 & n1521;
  assign n1523 = ~n1502 & n1522;
  assign n1524 = ~n1500 & n1523;
  assign n1525 = ~n1498 & n1524;
  assign n1526 = ~n1496 & n1525;
  assign n1527 = ~n1494 & n1526;
  assign n1528 = ~n1492 & n1527;
  assign n1529 = ~n1468 & n1483;
  assign n1530 = n1465 & n1468;
  assign n1531 = ~n1453 & n1472;
  assign n1532 = n1470 & n1480;
  assign n1533 = ~n1471 & n1528;
  assign n1534 = ~n1470 & n1533;
  assign n1535 = ~n1469 & n1534;
  assign n1536 = ~n1462 & n1535;
  assign n1537 = ~n1461 & n1536;
  assign n1538 = n1453 & ~n1528;
  assign n1539 = ~n1481 & n1538;
  assign n1540 = ~n1530 & n1539;
  assign n1541 = ~n1529 & n1540;
  assign n1542 = ~n1470 & n1476;
  assign n1543 = ~n1469 & n1542;
  assign n1544 = n1531 & n1543;
  assign n1545 = n1475 & ~n1528;
  assign n1546 = n1471 & n1545;
  assign n1547 = n1530 & n1546;
  assign n1548 = n1465 & n1528;
  assign n1549 = ~n1475 & n1548;
  assign n1550 = n1471 & n1549;
  assign n1551 = n1484 & n1512;
  assign n1552 = n1475 & ~n1481;
  assign n1553 = n1461 & n1552;
  assign n1554 = ~n1471 & n1529;
  assign n1555 = ~n1531 & n1554;
  assign n1556 = ~n1465 & ~n1476;
  assign n1557 = n1531 & n1556;
  assign n1558 = n1484 & n1532;
  assign n1559 = n1471 & n1481;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1557 & n1560;
  assign n1562 = ~n1555 & n1561;
  assign n1563 = ~n1553 & n1562;
  assign n1564 = ~n1551 & n1563;
  assign n1565 = ~n1550 & n1564;
  assign n1566 = ~n1547 & n1565;
  assign n1567 = ~n1544 & n1566;
  assign n1568 = ~n1541 & n1567;
  assign n1569 = ~n1537 & n1568;
  assign n1570 = ~\data<28>  & ~n1569;
  assign n1571 = \data<28>  & n1569;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = n504 & ~n1572;
  assign n1574 = \outreg<39>  & n508;
  assign n1575 = \outreg<31>  & ~\count<0> ;
  assign n1576 = ~n1574 & ~n1575;
  assign \outreg_new<31>  = n1573 | ~n1576;
  assign n1578 = \outreg<40>  & n508;
  assign n1579 = \outreg<32>  & ~\count<0> ;
  assign n1580 = \data<35>  & n504;
  assign n1581 = ~n1579 & ~n1580;
  assign \outreg_new<32>  = n1578 | ~n1581;
  assign n1583 = ~\data<3>  & ~n1528;
  assign n1584 = \data<3>  & n1528;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = n504 & ~n1585;
  assign n1587 = \outreg<41>  & n508;
  assign n1588 = \outreg<33>  & ~\count<0> ;
  assign n1589 = ~n1587 & ~n1588;
  assign \outreg_new<33>  = n1586 | ~n1589;
  assign n1591 = \outreg<42>  & n508;
  assign n1592 = \outreg<34>  & ~\count<0> ;
  assign n1593 = \data<43>  & n504;
  assign n1594 = ~n1592 & ~n1593;
  assign \outreg_new<34>  = n1591 | ~n1594;
  assign n1596 = \outreg<38>  & n508;
  assign n1597 = \outreg<30>  & ~\count<0> ;
  assign n1598 = \data<60>  & n504;
  assign n1599 = ~n1597 & ~n1598;
  assign \outreg_new<30>  = n1596 | ~n1599;
  assign n1601 = ~n1360 & n1383;
  assign n1602 = n1382 & n1388;
  assign n1603 = n1367 & n1371;
  assign n1604 = ~n1367 & ~n1385;
  assign n1605 = ~n1364 & n1604;
  assign n1606 = ~n1390 & n1605;
  assign n1607 = ~n1601 & n1606;
  assign n1608 = ~n1372 & n1607;
  assign n1609 = n1360 & n1367;
  assign n1610 = ~n1373 & n1609;
  assign n1611 = ~n1393 & n1610;
  assign n1612 = ~n1384 & n1611;
  assign n1613 = ~n1360 & n1373;
  assign n1614 = n1603 & n1613;
  assign n1615 = ~n1602 & n1614;
  assign n1616 = ~n1601 & n1615;
  assign n1617 = ~n1374 & ~n1603;
  assign n1618 = n1601 & n1617;
  assign n1619 = ~n1384 & n1618;
  assign n1620 = n1367 & ~n1373;
  assign n1621 = n1602 & n1620;
  assign n1622 = ~n1384 & n1621;
  assign n1623 = ~n1373 & n1385;
  assign n1624 = ~n1376 & n1623;
  assign n1625 = ~n1384 & n1624;
  assign n1626 = ~n1360 & ~n1382;
  assign n1627 = n1375 & n1626;
  assign n1628 = n1384 & n1627;
  assign n1629 = n1360 & n1393;
  assign n1630 = ~n1390 & n1629;
  assign n1631 = ~n1372 & n1630;
  assign n1632 = n1364 & n1383;
  assign n1633 = n1384 & n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign n1635 = ~n1628 & n1634;
  assign n1636 = ~n1625 & n1635;
  assign n1637 = ~n1622 & n1636;
  assign n1638 = ~n1619 & n1637;
  assign n1639 = ~n1616 & n1638;
  assign n1640 = ~n1612 & n1639;
  assign n1641 = ~n1608 & n1640;
  assign n1642 = ~\data<27>  & ~n1641;
  assign n1643 = \data<27>  & n1641;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = n504 & ~n1644;
  assign n1646 = \outreg<47>  & n508;
  assign n1647 = \outreg<39>  & ~\count<0> ;
  assign n1648 = ~n1646 & ~n1647;
  assign \outreg_new<39>  = n1645 | ~n1648;
  assign n1650 = ~\data<11>  & ~n1169;
  assign n1651 = \data<11>  & n1169;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n504 & ~n1652;
  assign n1654 = \outreg<43>  & n508;
  assign n1655 = \outreg<35>  & ~\count<0> ;
  assign n1656 = ~n1654 & ~n1655;
  assign \outreg_new<35>  = n1653 | ~n1656;
  assign n1658 = \outreg<44>  & n508;
  assign n1659 = \outreg<36>  & ~\count<0> ;
  assign n1660 = \data<51>  & n504;
  assign n1661 = ~n1659 & ~n1660;
  assign \outreg_new<36>  = n1658 | ~n1661;
  assign n1663 = \data<48>  & ~\C<1> ;
  assign n1664 = ~\data<48>  & \C<1> ;
  assign n1665 = ~n1663 & ~n1664;
  assign n1666 = ~\C<12>  & \data<47> ;
  assign n1667 = \C<12>  & ~\data<47> ;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~n1665 & ~n1668;
  assign n1670 = \data<44>  & ~\C<6> ;
  assign n1671 = ~\data<44>  & \C<6> ;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~\C<15>  & \data<43> ;
  assign n1674 = \C<15>  & ~\data<43> ;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~n1672 & ~n1675;
  assign n1677 = ~\C<19>  & \data<46> ;
  assign n1678 = \C<19>  & ~\data<46> ;
  assign n1679 = ~n1677 & ~n1678;
  assign n1680 = ~\C<26>  & \data<45> ;
  assign n1681 = \C<26>  & ~\data<45> ;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = ~n1672 & n1675;
  assign n1684 = ~n1682 & n1683;
  assign n1685 = n1668 & n1679;
  assign n1686 = n1665 & n1685;
  assign n1687 = n1684 & n1686;
  assign n1688 = n1675 & n1682;
  assign n1689 = n1679 & n1688;
  assign n1690 = n1665 & ~n1668;
  assign n1691 = n1665 & n1672;
  assign n1692 = ~n1668 & n1691;
  assign n1693 = ~n1675 & ~n1682;
  assign n1694 = n1679 & n1693;
  assign n1695 = n1692 & n1694;
  assign n1696 = ~n1665 & n1672;
  assign n1697 = n1685 & n1696;
  assign n1698 = n1676 & n1682;
  assign n1699 = ~n1679 & n1698;
  assign n1700 = ~n1665 & n1668;
  assign n1701 = n1668 & n1691;
  assign n1702 = ~n1675 & n1682;
  assign n1703 = n1669 & n1679;
  assign n1704 = ~n1679 & ~n1682;
  assign n1705 = n1669 & n1676;
  assign n1706 = n1704 & n1705;
  assign n1707 = ~n1675 & n1704;
  assign n1708 = n1672 & n1700;
  assign n1709 = n1707 & n1708;
  assign n1710 = n1683 & n1704;
  assign n1711 = n1700 & n1710;
  assign n1712 = n1672 & n1675;
  assign n1713 = ~n1682 & n1703;
  assign n1714 = n1712 & n1713;
  assign n1715 = ~n1679 & n1682;
  assign n1716 = ~n1676 & n1715;
  assign n1717 = n1669 & n1716;
  assign n1718 = n1679 & ~n1682;
  assign n1719 = ~n1665 & n1718;
  assign n1720 = n1676 & n1719;
  assign n1721 = n1665 & ~n1687;
  assign n1722 = n1684 & n1721;
  assign n1723 = ~n1665 & ~n1672;
  assign n1724 = n1689 & n1723;
  assign n1725 = ~n1672 & ~n1679;
  assign n1726 = n1690 & n1725;
  assign n1727 = n1679 & ~n1695;
  assign n1728 = n1692 & n1727;
  assign n1729 = n1691 & ~n1695;
  assign n1730 = n1693 & n1729;
  assign n1731 = n1675 & n1697;
  assign n1732 = n1699 & n1700;
  assign n1733 = n1676 & n1686;
  assign n1734 = n1688 & n1701;
  assign n1735 = n1702 & n1703;
  assign n1736 = ~n1711 & ~n1714;
  assign n1737 = ~n1709 & n1736;
  assign n1738 = ~n1706 & n1737;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = ~n1734 & n1739;
  assign n1741 = ~n1733 & n1740;
  assign n1742 = ~n1732 & n1741;
  assign n1743 = ~n1731 & n1742;
  assign n1744 = ~n1730 & n1743;
  assign n1745 = ~n1728 & n1744;
  assign n1746 = ~n1726 & n1745;
  assign n1747 = ~n1724 & n1746;
  assign n1748 = ~n1722 & n1747;
  assign n1749 = ~n1720 & n1748;
  assign n1750 = ~n1717 & n1749;
  assign n1751 = ~\data<19>  & ~n1750;
  assign n1752 = \data<19>  & n1750;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = n504 & ~n1753;
  assign n1755 = \outreg<45>  & n508;
  assign n1756 = \outreg<37>  & ~\count<0> ;
  assign n1757 = ~n1755 & ~n1756;
  assign \outreg_new<37>  = n1754 | ~n1757;
  assign n1759 = \outreg<46>  & n508;
  assign n1760 = \outreg<38>  & ~\count<0> ;
  assign n1761 = \data<59>  & n504;
  assign n1762 = ~n1760 & ~n1761;
  assign \outreg_new<38>  = n1759 | ~n1762;
  assign n1764 = n811 & n814;
  assign n1765 = n810 & n811;
  assign n1766 = ~n788 & n808;
  assign n1767 = n797 & ~n800;
  assign n1768 = n788 & ~n812;
  assign n1769 = ~n797 & n1768;
  assign n1770 = ~n796 & n1769;
  assign n1771 = ~n1764 & n1770;
  assign n1772 = ~n797 & ~n800;
  assign n1773 = n807 & n1772;
  assign n1774 = ~n1765 & n1773;
  assign n1775 = ~n797 & n811;
  assign n1776 = ~n796 & n1775;
  assign n1777 = n806 & n1776;
  assign n1778 = n797 & ~n803;
  assign n1779 = n806 & n1778;
  assign n1780 = ~n800 & n814;
  assign n1781 = n789 & n1780;
  assign n1782 = n807 & n825;
  assign n1783 = ~n785 & n812;
  assign n1784 = n796 & n1783;
  assign n1785 = ~n795 & n813;
  assign n1786 = n808 & n1785;
  assign n1787 = n810 & n1766;
  assign n1788 = n804 & n1767;
  assign n1789 = n805 & n1767;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1787 & n1790;
  assign n1792 = ~n1786 & n1791;
  assign n1793 = ~n1784 & n1792;
  assign n1794 = ~n1782 & n1793;
  assign n1795 = ~n1781 & n1794;
  assign n1796 = ~n1779 & n1795;
  assign n1797 = ~n1777 & n1796;
  assign n1798 = ~n1774 & n1797;
  assign n1799 = ~n1771 & n1798;
  assign n1800 = ~\data<2>  & ~n1799;
  assign n1801 = \data<2>  & n1799;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n504 & ~n1802;
  assign n1804 = \outreg<49>  & n508;
  assign n1805 = \outreg<41>  & ~\count<0> ;
  assign n1806 = ~n1804 & ~n1805;
  assign \outreg_new<41>  = n1803 | ~n1806;
  assign n1808 = \outreg<50>  & n508;
  assign n1809 = \outreg<42>  & ~\count<0> ;
  assign n1810 = \data<42>  & n504;
  assign n1811 = ~n1809 & ~n1810;
  assign \outreg_new<42>  = n1808 | ~n1811;
  assign n1813 = n1529 & n1531;
  assign n1814 = n1457 & n1470;
  assign n1815 = n1482 & n1814;
  assign n1816 = n1486 & n1497;
  assign n1817 = n1488 & n1529;
  assign n1818 = n1471 & n1485;
  assign n1819 = n1456 & n1460;
  assign n1820 = n1529 & n1819;
  assign n1821 = ~n1457 & n1482;
  assign n1822 = n1530 & n1821;
  assign n1823 = n1456 & n1480;
  assign n1824 = n1530 & n1823;
  assign n1825 = n1460 & n1462;
  assign n1826 = n1486 & n1825;
  assign n1827 = n1460 & n1478;
  assign n1828 = n1462 & n1827;
  assign n1829 = ~n1460 & ~n1471;
  assign n1830 = n1481 & n1829;
  assign n1831 = n1457 & n1469;
  assign n1832 = n1482 & n1831;
  assign n1833 = ~n1456 & n1480;
  assign n1834 = n1469 & n1833;
  assign n1835 = n1471 & ~n1475;
  assign n1836 = n1478 & n1835;
  assign n1837 = n1453 & n1532;
  assign n1838 = n1461 & n1486;
  assign n1839 = n1471 & n1529;
  assign n1840 = n1457 & n1479;
  assign n1841 = ~n1465 & n1477;
  assign n1842 = ~n1489 & ~n1818;
  assign n1843 = ~n1817 & n1842;
  assign n1844 = ~n1816 & n1843;
  assign n1845 = ~n1815 & n1844;
  assign n1846 = ~n1813 & n1845;
  assign n1847 = ~n1841 & n1846;
  assign n1848 = ~n1840 & n1847;
  assign n1849 = ~n1839 & n1848;
  assign n1850 = ~n1838 & n1849;
  assign n1851 = ~n1837 & n1850;
  assign n1852 = ~n1836 & n1851;
  assign n1853 = ~n1834 & n1852;
  assign n1854 = ~n1832 & n1853;
  assign n1855 = ~n1830 & n1854;
  assign n1856 = ~n1828 & n1855;
  assign n1857 = ~n1826 & n1856;
  assign n1858 = ~n1824 & n1857;
  assign n1859 = ~n1822 & n1858;
  assign n1860 = ~n1820 & n1859;
  assign n1861 = ~\data<10>  & ~n1860;
  assign n1862 = \data<10>  & n1860;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = n504 & ~n1863;
  assign n1865 = \outreg<51>  & n508;
  assign n1866 = \outreg<43>  & ~\count<0> ;
  assign n1867 = ~n1865 & ~n1866;
  assign \outreg_new<43>  = n1864 | ~n1867;
  assign n1869 = \outreg<52>  & n508;
  assign n1870 = \outreg<44>  & ~\count<0> ;
  assign n1871 = \data<50>  & n504;
  assign n1872 = ~n1870 & ~n1871;
  assign \outreg_new<44>  = n1869 | ~n1872;
  assign n1874 = \outreg<48>  & n508;
  assign n1875 = \outreg<40>  & ~\count<0> ;
  assign n1876 = \data<34>  & n504;
  assign n1877 = ~n1875 & ~n1876;
  assign \outreg_new<40>  = n1874 | ~n1877;
  assign n1879 = ~n1363 & n1603;
  assign n1880 = n1364 & n1603;
  assign n1881 = n1383 & n1880;
  assign n1882 = n1360 & n1383;
  assign n1883 = ~n1375 & n1882;
  assign n1884 = ~n1374 & n1883;
  assign n1885 = ~n1879 & n1884;
  assign n1886 = ~n1393 & ~n1881;
  assign n1887 = ~n1389 & n1886;
  assign n1888 = n1879 & n1887;
  assign n1889 = ~n1371 & ~n1382;
  assign n1890 = n1368 & n1889;
  assign n1891 = ~n1382 & n1391;
  assign n1892 = n1374 & n1891;
  assign n1893 = n1374 & n1386;
  assign n1894 = n1364 & n1375;
  assign n1895 = n1393 & n1894;
  assign n1896 = n1363 & ~n1375;
  assign n1897 = n1393 & n1896;
  assign n1898 = ~n1363 & n1382;
  assign n1899 = n1391 & n1898;
  assign n1900 = n1375 & ~n1379;
  assign n1901 = n1364 & n1900;
  assign n1902 = n1375 & n1389;
  assign n1903 = n1376 & n1385;
  assign n1904 = ~n1395 & ~n1903;
  assign n1905 = n1390 & n1601;
  assign n1906 = n1904 & ~n1905;
  assign n1907 = ~n1902 & n1906;
  assign n1908 = ~n1901 & n1907;
  assign n1909 = ~n1899 & n1908;
  assign n1910 = ~n1897 & n1909;
  assign n1911 = ~n1895 & n1910;
  assign n1912 = ~n1893 & n1911;
  assign n1913 = ~n1892 & n1912;
  assign n1914 = ~n1890 & n1913;
  assign n1915 = ~n1888 & n1914;
  assign n1916 = ~n1885 & n1915;
  assign n1917 = ~\data<1>  & ~n1916;
  assign n1918 = \data<1>  & n1916;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = n504 & ~n1919;
  assign n1921 = \outreg<57>  & n508;
  assign n1922 = \outreg<49>  & ~\count<0> ;
  assign n1923 = ~n1921 & ~n1922;
  assign \outreg_new<49>  = n1920 | ~n1923;
  assign n1925 = n1457 & n1460;
  assign n1926 = ~n1470 & n1925;
  assign n1927 = ~n1469 & n1926;
  assign n1928 = ~n1485 & n1927;
  assign n1929 = ~n1460 & ~n1478;
  assign n1930 = ~n1476 & n1929;
  assign n1931 = ~n1530 & n1930;
  assign n1932 = ~n1487 & n1931;
  assign n1933 = n1461 & n1481;
  assign n1934 = n1465 & n1484;
  assign n1935 = ~n1457 & n1485;
  assign n1936 = ~n1456 & n1532;
  assign n1937 = n1486 & n1487;
  assign n1938 = n1486 & n1531;
  assign n1939 = ~n1470 & n1477;
  assign n1940 = n1476 & n1478;
  assign n1941 = n1470 & n1471;
  assign n1942 = ~n1817 & ~n1941;
  assign n1943 = ~n1940 & n1942;
  assign n1944 = ~n1939 & n1943;
  assign n1945 = ~n1938 & n1944;
  assign n1946 = ~n1937 & n1945;
  assign n1947 = ~n1936 & n1946;
  assign n1948 = ~n1935 & n1947;
  assign n1949 = ~n1934 & n1948;
  assign n1950 = ~n1933 & n1949;
  assign n1951 = ~n1932 & n1950;
  assign n1952 = ~n1928 & n1951;
  assign n1953 = ~\data<18>  & ~n1952;
  assign n1954 = \data<18>  & n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = n504 & ~n1955;
  assign n1957 = \outreg<53>  & n508;
  assign n1958 = \outreg<45>  & ~\count<0> ;
  assign n1959 = ~n1957 & ~n1958;
  assign \outreg_new<45>  = n1956 | ~n1959;
  assign n1961 = \outreg<54>  & n508;
  assign n1962 = \outreg<46>  & ~\count<0> ;
  assign n1963 = \data<58>  & n504;
  assign n1964 = ~n1962 & ~n1963;
  assign \outreg_new<46>  = n1961 | ~n1964;
  assign n1966 = ~\data<26>  & ~n601;
  assign n1967 = \data<26>  & n601;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = n504 & ~n1968;
  assign n1970 = \outreg<55>  & n508;
  assign n1971 = \outreg<47>  & ~\count<0> ;
  assign n1972 = ~n1970 & ~n1971;
  assign \outreg_new<47>  = n1969 | ~n1972;
  assign n1974 = \outreg<56>  & n508;
  assign n1975 = \outreg<48>  & ~\count<0> ;
  assign n1976 = \data<33>  & n504;
  assign n1977 = ~n1975 & ~n1976;
  assign \outreg_new<48>  = n1974 | ~n1977;
  assign n1979 = \encrypt_mode<0>  & ~\encrypt<0> ;
  assign n1980 = n504 & n1979;
  assign n1981 = ~\encrypt_mode<0>  & \encrypt<0> ;
  assign n1982 = n504 & n1981;
  assign n1983 = ~n1980 & ~n1982;
  assign n1984 = n645 & n1983;
  assign n1985 = ~\encrypt_mode<0>  & n1984;
  assign n1986 = ~n745 & n1985;
  assign n1987 = \encrypt_mode<0>  & n1984;
  assign n1988 = ~n745 & n1987;
  assign n1989 = n745 & n1987;
  assign n1990 = n745 & n1985;
  assign n1991 = n645 & ~n1983;
  assign n1992 = ~\reset<0>  & n644;
  assign n1993 = \encrypt<0>  & n1992;
  assign n1994 = ~\encrypt<0>  & n1992;
  assign n1995 = \C<22>  & n1986;
  assign n1996 = \C<24>  & n1988;
  assign n1997 = \C<25>  & n1989;
  assign n1998 = \C<21>  & n1990;
  assign n1999 = \C<23>  & n1991;
  assign n2000 = \inreg<51>  & n1993;
  assign n2001 = \data_in<2>  & n1994;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1999 & n2002;
  assign n2004 = ~n1998 & n2003;
  assign n2005 = ~n1997 & n2004;
  assign n2006 = ~n1996 & n2005;
  assign \C_new<23>  = n1995 | ~n2006;
  assign n2008 = \C<23>  & n1986;
  assign n2009 = \C<25>  & n1988;
  assign n2010 = \C<26>  & n1989;
  assign n2011 = \C<22>  & n1990;
  assign n2012 = \C<24>  & n1991;
  assign n2013 = \inreg<43>  & n1993;
  assign n2014 = \inreg<51>  & n1994;
  assign n2015 = ~n2013 & ~n2014;
  assign n2016 = ~n2012 & n2015;
  assign n2017 = ~n2011 & n2016;
  assign n2018 = ~n2010 & n2017;
  assign n2019 = ~n2009 & n2018;
  assign \C_new<24>  = n2008 | ~n2019;
  assign n2021 = \C<20>  & n1986;
  assign n2022 = \C<22>  & n1988;
  assign n2023 = \C<23>  & n1989;
  assign n2024 = \C<19>  & n1990;
  assign n2025 = \C<21>  & n1991;
  assign n2026 = \inreg<2>  & n1993;
  assign n2027 = \inreg<10>  & n1994;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = ~n2025 & n2028;
  assign n2030 = ~n2024 & n2029;
  assign n2031 = ~n2023 & n2030;
  assign n2032 = ~n2022 & n2031;
  assign \C_new<21>  = n2021 | ~n2032;
  assign n2034 = \C<21>  & n1986;
  assign n2035 = \C<23>  & n1988;
  assign n2036 = \C<24>  & n1989;
  assign n2037 = \C<20>  & n1990;
  assign n2038 = \C<22>  & n1991;
  assign n2039 = \data_in<2>  & n1993;
  assign n2040 = \inreg<2>  & n1994;
  assign n2041 = ~n2039 & ~n2040;
  assign n2042 = ~n2038 & n2041;
  assign n2043 = ~n2037 & n2042;
  assign n2044 = ~n2036 & n2043;
  assign n2045 = ~n2035 & n2044;
  assign \C_new<22>  = n2034 | ~n2045;
  assign n2047 = \C<19>  & n1986;
  assign n2048 = \C<21>  & n1988;
  assign n2049 = \C<22>  & n1989;
  assign n2050 = \C<18>  & n1990;
  assign n2051 = \C<20>  & n1991;
  assign n2052 = \inreg<10>  & n1993;
  assign n2053 = \inreg<18>  & n1994;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = ~n2051 & n2054;
  assign n2056 = ~n2050 & n2055;
  assign n2057 = ~n2049 & n2056;
  assign n2058 = ~n2048 & n2057;
  assign \C_new<20>  = n2047 | ~n2058;
  assign n2060 = \inreg<17>  & n504;
  assign n2061 = \data<36>  & ~n504;
  assign \data_new<4>  = n2060 | n2061;
  assign n2063 = \inreg<25>  & n504;
  assign n2064 = \data<35>  & ~n504;
  assign \data_new<3>  = n2063 | n2064;
  assign n2066 = \C<26>  & n1986;
  assign n2067 = \C<0>  & n1988;
  assign n2068 = \C<1>  & n1989;
  assign n2069 = \C<25>  & n1990;
  assign n2070 = \C<27>  & n1991;
  assign n2071 = \inreg<48>  & n1993;
  assign n2072 = \inreg<27>  & n1994;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2070 & n2073;
  assign n2075 = ~n2069 & n2074;
  assign n2076 = ~n2068 & n2075;
  assign n2077 = ~n2067 & n2076;
  assign \C_new<27>  = n2066 | ~n2077;
  assign n2079 = \inreg<33>  & n504;
  assign n2080 = \data<34>  & ~n504;
  assign \data_new<2>  = n2079 | n2080;
  assign n2082 = \inreg<41>  & n504;
  assign n2083 = \data<33>  & ~n504;
  assign \data_new<1>  = n2082 | n2083;
  assign n2085 = \C<24>  & n1986;
  assign n2086 = \C<26>  & n1988;
  assign n2087 = \C<27>  & n1989;
  assign n2088 = \C<23>  & n1990;
  assign n2089 = \C<25>  & n1991;
  assign n2090 = \inreg<35>  & n1993;
  assign n2091 = \inreg<43>  & n1994;
  assign n2092 = ~n2090 & ~n2091;
  assign n2093 = ~n2089 & n2092;
  assign n2094 = ~n2088 & n2093;
  assign n2095 = ~n2087 & n2094;
  assign n2096 = ~n2086 & n2095;
  assign \C_new<25>  = n2085 | ~n2096;
  assign n2098 = \inreg<49>  & n504;
  assign n2099 = \data<32>  & ~n504;
  assign \data_new<0>  = n2098 | n2099;
  assign n2101 = \C<25>  & n1986;
  assign n2102 = \C<27>  & n1988;
  assign n2103 = \C<0>  & n1989;
  assign n2104 = \C<24>  & n1990;
  assign n2105 = \C<26>  & n1991;
  assign n2106 = \inreg<27>  & n1993;
  assign n2107 = \inreg<35>  & n1994;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = ~n2105 & n2108;
  assign n2110 = ~n2104 & n2109;
  assign n2111 = ~n2103 & n2110;
  assign n2112 = ~n2102 & n2111;
  assign \C_new<26>  = n2101 | ~n2112;
  assign n2114 = \C<12>  & n1986;
  assign n2115 = \C<14>  & n1988;
  assign n2116 = \C<15>  & n1989;
  assign n2117 = \C<11>  & n1990;
  assign n2118 = \C<13>  & n1991;
  assign n2119 = \inreg<1>  & n1993;
  assign n2120 = \inreg<9>  & n1994;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~n2118 & n2121;
  assign n2123 = ~n2117 & n2122;
  assign n2124 = ~n2116 & n2123;
  assign n2125 = ~n2115 & n2124;
  assign \C_new<13>  = n2114 | ~n2125;
  assign n2127 = \C<13>  & n1986;
  assign n2128 = \C<15>  & n1988;
  assign n2129 = \C<16>  & n1989;
  assign n2130 = \C<12>  & n1990;
  assign n2131 = \C<14>  & n1991;
  assign n2132 = \data_in<1>  & n1993;
  assign n2133 = \inreg<1>  & n1994;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~n2131 & n2134;
  assign n2136 = ~n2130 & n2135;
  assign n2137 = ~n2129 & n2136;
  assign n2138 = ~n2128 & n2137;
  assign \C_new<14>  = n2127 | ~n2138;
  assign n2140 = \C<10>  & n1986;
  assign n2141 = \C<12>  & n1988;
  assign n2142 = \C<13>  & n1989;
  assign n2143 = \C<9>  & n1990;
  assign n2144 = \C<11>  & n1991;
  assign n2145 = \inreg<17>  & n1993;
  assign n2146 = \inreg<25>  & n1994;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2144 & n2147;
  assign n2149 = ~n2143 & n2148;
  assign n2150 = ~n2142 & n2149;
  assign n2151 = ~n2141 & n2150;
  assign \C_new<11>  = n2140 | ~n2151;
  assign n2153 = \C<11>  & n1986;
  assign n2154 = \C<13>  & n1988;
  assign n2155 = \C<14>  & n1989;
  assign n2156 = \C<10>  & n1990;
  assign n2157 = \C<12>  & n1991;
  assign n2158 = \inreg<9>  & n1993;
  assign n2159 = \inreg<17>  & n1994;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = ~n2157 & n2160;
  assign n2162 = ~n2156 & n2161;
  assign n2163 = ~n2155 & n2162;
  assign n2164 = ~n2154 & n2163;
  assign \C_new<12>  = n2153 | ~n2164;
  assign n2166 = \C<9>  & n1986;
  assign n2167 = \C<11>  & n1988;
  assign n2168 = \C<12>  & n1989;
  assign n2169 = \C<8>  & n1990;
  assign n2170 = \C<10>  & n1991;
  assign n2171 = \inreg<25>  & n1993;
  assign n2172 = \inreg<33>  & n1994;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = ~n2170 & n2173;
  assign n2175 = ~n2169 & n2174;
  assign n2176 = ~n2168 & n2175;
  assign n2177 = ~n2167 & n2176;
  assign \C_new<10>  = n2166 | ~n2177;
  assign n2179 = \inreg<43>  & n504;
  assign n2180 = \data<41>  & ~n504;
  assign \data_new<9>  = n2179 | n2180;
  assign n2182 = \inreg<51>  & n504;
  assign n2183 = \data<40>  & ~n504;
  assign \data_new<8>  = n2182 | n2183;
  assign n2185 = \data_in<1>  & n504;
  assign n2186 = \data<39>  & ~n504;
  assign \data_new<7>  = n2185 | n2186;
  assign n2188 = \inreg<1>  & n504;
  assign n2189 = \data<38>  & ~n504;
  assign \data_new<6>  = n2188 | n2189;
  assign n2191 = \inreg<9>  & n504;
  assign n2192 = \data<37>  & ~n504;
  assign \data_new<5>  = n2191 | n2192;
  assign n2194 = \C<18>  & n1986;
  assign n2195 = \C<20>  & n1988;
  assign n2196 = \C<21>  & n1989;
  assign n2197 = \C<17>  & n1990;
  assign n2198 = \C<19>  & n1991;
  assign n2199 = \inreg<18>  & n1993;
  assign n2200 = \inreg<26>  & n1994;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~n2198 & n2201;
  assign n2203 = ~n2197 & n2202;
  assign n2204 = ~n2196 & n2203;
  assign n2205 = ~n2195 & n2204;
  assign \C_new<19>  = n2194 | ~n2205;
  assign n2207 = \C<16>  & n1986;
  assign n2208 = \C<18>  & n1988;
  assign n2209 = \C<19>  & n1989;
  assign n2210 = \C<15>  & n1990;
  assign n2211 = \C<17>  & n1991;
  assign n2212 = \inreg<34>  & n1993;
  assign n2213 = \inreg<42>  & n1994;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n2211 & n2214;
  assign n2216 = ~n2210 & n2215;
  assign n2217 = ~n2209 & n2216;
  assign n2218 = ~n2208 & n2217;
  assign \C_new<17>  = n2207 | ~n2218;
  assign n2220 = \C<17>  & n1986;
  assign n2221 = \C<19>  & n1988;
  assign n2222 = \C<20>  & n1989;
  assign n2223 = \C<16>  & n1990;
  assign n2224 = \C<18>  & n1991;
  assign n2225 = \inreg<26>  & n1993;
  assign n2226 = \inreg<34>  & n1994;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = ~n2224 & n2227;
  assign n2229 = ~n2223 & n2228;
  assign n2230 = ~n2222 & n2229;
  assign n2231 = ~n2221 & n2230;
  assign \C_new<18>  = n2220 | ~n2231;
  assign n2233 = \C<14>  & n1986;
  assign n2234 = \C<16>  & n1988;
  assign n2235 = \C<17>  & n1989;
  assign n2236 = \C<13>  & n1990;
  assign n2237 = \C<15>  & n1991;
  assign n2238 = \inreg<50>  & n1993;
  assign n2239 = \data_in<1>  & n1994;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n2237 & n2240;
  assign n2242 = ~n2236 & n2241;
  assign n2243 = ~n2235 & n2242;
  assign n2244 = ~n2234 & n2243;
  assign \C_new<15>  = n2233 | ~n2244;
  assign n2246 = \C<15>  & n1986;
  assign n2247 = \C<17>  & n1988;
  assign n2248 = \C<18>  & n1989;
  assign n2249 = \C<14>  & n1990;
  assign n2250 = \C<16>  & n1991;
  assign n2251 = \inreg<42>  & n1993;
  assign n2252 = \inreg<50>  & n1994;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = ~n2250 & n2253;
  assign n2255 = ~n2249 & n2254;
  assign n2256 = ~n2248 & n2255;
  assign n2257 = ~n2247 & n2256;
  assign \C_new<16>  = n2246 | ~n2257;
  assign n2259 = \D<12>  & n1986;
  assign n2260 = \D<14>  & n1988;
  assign n2261 = \D<15>  & n1989;
  assign n2262 = \D<11>  & n1990;
  assign n2263 = \D<13>  & n1991;
  assign n2264 = \inreg<5>  & n1993;
  assign n2265 = \inreg<13>  & n1994;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n2263 & n2266;
  assign n2268 = ~n2262 & n2267;
  assign n2269 = ~n2261 & n2268;
  assign n2270 = ~n2260 & n2269;
  assign \D_new<13>  = n2259 | ~n2270;
  assign n2272 = \D<13>  & n1986;
  assign n2273 = \D<15>  & n1988;
  assign n2274 = \D<16>  & n1989;
  assign n2275 = \D<12>  & n1990;
  assign n2276 = \D<14>  & n1991;
  assign n2277 = \data_in<5>  & n1993;
  assign n2278 = \inreg<5>  & n1994;
  assign n2279 = ~n2277 & ~n2278;
  assign n2280 = ~n2276 & n2279;
  assign n2281 = ~n2275 & n2280;
  assign n2282 = ~n2274 & n2281;
  assign n2283 = ~n2273 & n2282;
  assign \D_new<14>  = n2272 | ~n2283;
  assign n2285 = \D<10>  & n1986;
  assign n2286 = \D<12>  & n1988;
  assign n2287 = \D<13>  & n1989;
  assign n2288 = \D<9>  & n1990;
  assign n2289 = \D<11>  & n1991;
  assign n2290 = \inreg<21>  & n1993;
  assign n2291 = \inreg<29>  & n1994;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = ~n2289 & n2292;
  assign n2294 = ~n2288 & n2293;
  assign n2295 = ~n2287 & n2294;
  assign n2296 = ~n2286 & n2295;
  assign \D_new<11>  = n2285 | ~n2296;
  assign n2298 = \D<11>  & n1986;
  assign n2299 = \D<13>  & n1988;
  assign n2300 = \D<14>  & n1989;
  assign n2301 = \D<10>  & n1990;
  assign n2302 = \D<12>  & n1991;
  assign n2303 = \inreg<13>  & n1993;
  assign n2304 = \inreg<21>  & n1994;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n2302 & n2305;
  assign n2307 = ~n2301 & n2306;
  assign n2308 = ~n2300 & n2307;
  assign n2309 = ~n2299 & n2308;
  assign \D_new<12>  = n2298 | ~n2309;
  assign n2311 = \D<9>  & n1986;
  assign n2312 = \D<11>  & n1988;
  assign n2313 = \D<12>  & n1989;
  assign n2314 = \D<8>  & n1990;
  assign n2315 = \D<10>  & n1991;
  assign n2316 = \inreg<29>  & n1993;
  assign n2317 = \inreg<37>  & n1994;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = ~n2315 & n2318;
  assign n2320 = ~n2314 & n2319;
  assign n2321 = ~n2313 & n2320;
  assign n2322 = ~n2312 & n2321;
  assign \D_new<10>  = n2311 | ~n2322;
  assign n2324 = n1101 & n1130;
  assign n2325 = n1129 & n2324;
  assign n2326 = ~n1104 & n1169;
  assign n2327 = ~n1101 & n2326;
  assign n2328 = n1129 & n2327;
  assign n2329 = ~n1107 & ~n1169;
  assign n2330 = n1101 & n2329;
  assign n2331 = n1127 & n2330;
  assign n2332 = n1107 & n1194;
  assign n2333 = ~n1111 & n2332;
  assign n2334 = n1111 & n1135;
  assign n2335 = n1126 & n2334;
  assign n2336 = n1132 & ~n1137;
  assign n2337 = ~n1108 & n1132;
  assign n2338 = n1104 & n1173;
  assign n2339 = n1137 & n1169;
  assign n2340 = ~n1121 & n1125;
  assign n2341 = n1127 & n1171;
  assign n2342 = n1130 & n1133;
  assign n2343 = n1177 & ~n2325;
  assign n2344 = ~n2342 & n2343;
  assign n2345 = ~n2341 & n2344;
  assign n2346 = ~n2340 & n2345;
  assign n2347 = ~n2339 & n2346;
  assign n2348 = ~n2338 & n2347;
  assign n2349 = ~n1157 & n2348;
  assign n2350 = ~n2337 & n2349;
  assign n2351 = ~n2336 & n2350;
  assign n2352 = ~n2335 & n2351;
  assign n2353 = ~n2333 & n2352;
  assign n2354 = ~n2331 & n2353;
  assign n2355 = ~n2328 & n2354;
  assign n2356 = ~\data<31>  & ~n2355;
  assign n2357 = \data<31>  & n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n504 & ~n2358;
  assign n2360 = \data_in<6>  & n504;
  assign \data_new<63>  = n2359 | n2360;
  assign n2362 = ~n504 & ~n1230;
  assign n2363 = \inreg<14>  & n504;
  assign \data_new<61>  = n2362 | n2363;
  assign n2365 = ~n504 & ~n957;
  assign n2366 = \inreg<6>  & n504;
  assign \data_new<62>  = n2365 | n2366;
  assign n2368 = \D<18>  & n1986;
  assign n2369 = \D<20>  & n1988;
  assign n2370 = \D<21>  & n1989;
  assign n2371 = \D<17>  & n1990;
  assign n2372 = \D<19>  & n1991;
  assign n2373 = \inreg<20>  & n1993;
  assign n2374 = \inreg<28>  & n1994;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n2372 & n2375;
  assign n2377 = ~n2371 & n2376;
  assign n2378 = ~n2370 & n2377;
  assign n2379 = ~n2369 & n2378;
  assign \D_new<19>  = n2368 | ~n2379;
  assign n2381 = ~n504 & ~n1572;
  assign n2382 = \inreg<22>  & n504;
  assign \data_new<60>  = n2381 | n2382;
  assign n2384 = \D<16>  & n1986;
  assign n2385 = \D<18>  & n1988;
  assign n2386 = \D<19>  & n1989;
  assign n2387 = \D<15>  & n1990;
  assign n2388 = \D<17>  & n1991;
  assign n2389 = \inreg<36>  & n1993;
  assign n2390 = \inreg<44>  & n1994;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = ~n2388 & n2391;
  assign n2393 = ~n2387 & n2392;
  assign n2394 = ~n2386 & n2393;
  assign n2395 = ~n2385 & n2394;
  assign \D_new<17>  = n2384 | ~n2395;
  assign n2397 = \D<17>  & n1986;
  assign n2398 = \D<19>  & n1988;
  assign n2399 = \D<20>  & n1989;
  assign n2400 = \D<16>  & n1990;
  assign n2401 = \D<18>  & n1991;
  assign n2402 = \inreg<28>  & n1993;
  assign n2403 = \inreg<36>  & n1994;
  assign n2404 = ~n2402 & ~n2403;
  assign n2405 = ~n2401 & n2404;
  assign n2406 = ~n2400 & n2405;
  assign n2407 = ~n2399 & n2406;
  assign n2408 = ~n2398 & n2407;
  assign \D_new<18>  = n2397 | ~n2408;
  assign n2410 = \D<14>  & n1986;
  assign n2411 = \D<16>  & n1988;
  assign n2412 = \D<17>  & n1989;
  assign n2413 = \D<13>  & n1990;
  assign n2414 = \D<15>  & n1991;
  assign n2415 = \inreg<52>  & n1993;
  assign n2416 = \data_in<5>  & n1994;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = ~n2414 & n2417;
  assign n2419 = ~n2413 & n2418;
  assign n2420 = ~n2412 & n2419;
  assign n2421 = ~n2411 & n2420;
  assign \D_new<15>  = n2410 | ~n2421;
  assign n2423 = \D<15>  & n1986;
  assign n2424 = \D<17>  & n1988;
  assign n2425 = \D<18>  & n1989;
  assign n2426 = \D<14>  & n1990;
  assign n2427 = \D<16>  & n1991;
  assign n2428 = \inreg<44>  & n1993;
  assign n2429 = \inreg<52>  & n1994;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = ~n2427 & n2430;
  assign n2432 = ~n2426 & n2431;
  assign n2433 = ~n2425 & n2432;
  assign n2434 = ~n2424 & n2433;
  assign \D_new<16>  = n2423 | ~n2434;
  assign n2436 = \D<22>  & n1986;
  assign n2437 = \D<24>  & n1988;
  assign n2438 = \D<25>  & n1989;
  assign n2439 = \D<21>  & n1990;
  assign n2440 = \D<23>  & n1991;
  assign n2441 = \inreg<19>  & n1993;
  assign n2442 = \data_in<4>  & n1994;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2440 & n2443;
  assign n2445 = ~n2439 & n2444;
  assign n2446 = ~n2438 & n2445;
  assign n2447 = ~n2437 & n2446;
  assign \D_new<23>  = n2436 | ~n2447;
  assign n2449 = \D<23>  & n1986;
  assign n2450 = \D<25>  & n1988;
  assign n2451 = \D<26>  & n1989;
  assign n2452 = \D<22>  & n1990;
  assign n2453 = \D<24>  & n1991;
  assign n2454 = \inreg<11>  & n1993;
  assign n2455 = \inreg<19>  & n1994;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = ~n2453 & n2456;
  assign n2458 = ~n2452 & n2457;
  assign n2459 = ~n2451 & n2458;
  assign n2460 = ~n2450 & n2459;
  assign \D_new<24>  = n2449 | ~n2460;
  assign n2462 = \D<20>  & n1986;
  assign n2463 = \D<22>  & n1988;
  assign n2464 = \D<23>  & n1989;
  assign n2465 = \D<19>  & n1990;
  assign n2466 = \D<21>  & n1991;
  assign n2467 = \inreg<4>  & n1993;
  assign n2468 = \inreg<12>  & n1994;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = ~n2466 & n2469;
  assign n2471 = ~n2465 & n2470;
  assign n2472 = ~n2464 & n2471;
  assign n2473 = ~n2463 & n2472;
  assign \D_new<21>  = n2462 | ~n2473;
  assign n2475 = \D<21>  & n1986;
  assign n2476 = \D<23>  & n1988;
  assign n2477 = \D<24>  & n1989;
  assign n2478 = \D<20>  & n1990;
  assign n2479 = \D<22>  & n1991;
  assign n2480 = \data_in<4>  & n1993;
  assign n2481 = \inreg<4>  & n1994;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = ~n2479 & n2482;
  assign n2484 = ~n2478 & n2483;
  assign n2485 = ~n2477 & n2484;
  assign n2486 = ~n2476 & n2485;
  assign \D_new<22>  = n2475 | ~n2486;
  assign n2488 = \D<19>  & n1986;
  assign n2489 = \D<21>  & n1988;
  assign n2490 = \D<22>  & n1989;
  assign n2491 = \D<18>  & n1990;
  assign n2492 = \D<20>  & n1991;
  assign n2493 = \inreg<12>  & n1993;
  assign n2494 = \inreg<20>  & n1994;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2492 & n2495;
  assign n2497 = ~n2491 & n2496;
  assign n2498 = ~n2490 & n2497;
  assign n2499 = ~n2489 & n2498;
  assign \D_new<20>  = n2488 | ~n2499;
  assign n2501 = ~n504 & ~n1217;
  assign n2502 = \inreg<12>  & n504;
  assign \data_new<53>  = n2501 | n2502;
  assign n2504 = ~n504 & ~n726;
  assign n2505 = \inreg<4>  & n504;
  assign \data_new<54>  = n2504 | n2505;
  assign n2507 = ~n504 & ~n1753;
  assign n2508 = \inreg<28>  & n504;
  assign \data_new<51>  = n2507 | n2508;
  assign n2510 = ~n504 & ~n1290;
  assign n2511 = \inreg<20>  & n504;
  assign \data_new<52>  = n2510 | n2511;
  assign n2513 = ~n504 & ~n1955;
  assign n2514 = \inreg<36>  & n504;
  assign \data_new<50>  = n2513 | n2514;
  assign n2516 = \D<26>  & n1986;
  assign n2517 = \D<0>  & n1988;
  assign n2518 = \D<1>  & n1989;
  assign n2519 = \D<25>  & n1990;
  assign n2520 = \D<27>  & n1991;
  assign n2521 = \inreg<54>  & n1993;
  assign n2522 = \data_in<3>  & n1994;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = ~n2520 & n2523;
  assign n2525 = ~n2519 & n2524;
  assign n2526 = ~n2518 & n2525;
  assign n2527 = ~n2517 & n2526;
  assign \D_new<27>  = n2516 | ~n2527;
  assign n2529 = \D<24>  & n1986;
  assign n2530 = \D<26>  & n1988;
  assign n2531 = \D<27>  & n1989;
  assign n2532 = \D<23>  & n1990;
  assign n2533 = \D<25>  & n1991;
  assign n2534 = \inreg<3>  & n1993;
  assign n2535 = \inreg<11>  & n1994;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = ~n2533 & n2536;
  assign n2538 = ~n2532 & n2537;
  assign n2539 = ~n2531 & n2538;
  assign n2540 = ~n2530 & n2539;
  assign \D_new<25>  = n2529 | ~n2540;
  assign n2542 = \D<25>  & n1986;
  assign n2543 = \D<27>  & n1988;
  assign n2544 = \D<0>  & n1989;
  assign n2545 = \D<24>  & n1990;
  assign n2546 = \D<26>  & n1991;
  assign n2547 = \data_in<3>  & n1993;
  assign n2548 = \inreg<3>  & n1994;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = ~n2546 & n2549;
  assign n2551 = ~n2545 & n2550;
  assign n2552 = ~n2544 & n2551;
  assign n2553 = ~n2543 & n2552;
  assign \D_new<26>  = n2542 | ~n2553;
  assign n2555 = ~n504 & ~n1644;
  assign n2556 = \inreg<30>  & n504;
  assign \data_new<59>  = n2555 | n2556;
  assign n2558 = n1665 & n1668;
  assign n2559 = n1701 & n1707;
  assign n2560 = n1690 & n1699;
  assign n2561 = n1689 & n1692;
  assign n2562 = ~n1679 & ~n2559;
  assign n2563 = ~n1702 & n2562;
  assign n2564 = n2558 & n2563;
  assign n2565 = ~n1684 & n2564;
  assign n2566 = ~n1672 & ~n1688;
  assign n2567 = ~n1693 & n2566;
  assign n2568 = n1686 & n2567;
  assign n2569 = n1672 & ~n2559;
  assign n2570 = ~n1703 & n2569;
  assign n2571 = n1693 & n2570;
  assign n2572 = n1688 & n1700;
  assign n2573 = n1712 & n2572;
  assign n2574 = n1691 & n1704;
  assign n2575 = n1712 & n2574;
  assign n2576 = ~n1685 & ~n2558;
  assign n2577 = n1684 & n2576;
  assign n2578 = n1672 & n1703;
  assign n2579 = ~n1693 & n2578;
  assign n2580 = n1676 & n1685;
  assign n2581 = n1700 & n2580;
  assign n2582 = n1669 & n1725;
  assign n2583 = n1701 & n1702;
  assign n2584 = ~n2560 & ~n2561;
  assign n2585 = ~n2583 & n2584;
  assign n2586 = ~n2582 & n2585;
  assign n2587 = ~n2581 & n2586;
  assign n2588 = ~n2579 & n2587;
  assign n2589 = ~n2577 & n2588;
  assign n2590 = ~n2575 & n2589;
  assign n2591 = ~n2573 & n2590;
  assign n2592 = ~n2571 & n2591;
  assign n2593 = ~n2568 & n2592;
  assign n2594 = ~n2565 & n2593;
  assign n2595 = ~\data<25>  & ~n2594;
  assign n2596 = \data<25>  & n2594;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~n504 & ~n2597;
  assign n2599 = \inreg<46>  & n504;
  assign \data_new<57>  = n2598 | n2599;
  assign n2601 = ~n504 & ~n1968;
  assign n2602 = \inreg<38>  & n504;
  assign \data_new<58>  = n2601 | n2602;
  assign n2604 = n973 & n994;
  assign n2605 = ~n974 & n991;
  assign n2606 = n998 & n2605;
  assign n2607 = ~n2604 & n2606;
  assign n2608 = ~n1000 & n2607;
  assign n2609 = ~n970 & n1042;
  assign n2610 = ~n1003 & n2609;
  assign n2611 = ~n1002 & n2610;
  assign n2612 = ~n2604 & n2611;
  assign n2613 = n994 & n1003;
  assign n2614 = ~n1000 & n2613;
  assign n2615 = n970 & n990;
  assign n2616 = n986 & n2615;
  assign n2617 = n980 & n2616;
  assign n2618 = n1003 & ~n1042;
  assign n2619 = n1000 & n2618;
  assign n2620 = ~n980 & n990;
  assign n2621 = n993 & n2620;
  assign n2622 = n999 & ~n1042;
  assign n2623 = n1043 & n2622;
  assign n2624 = ~n980 & n1002;
  assign n2625 = n1004 & n2624;
  assign n2626 = n1001 & n1002;
  assign n2627 = n1005 & n2626;
  assign n2628 = ~n990 & ~n1042;
  assign n2629 = n974 & n2628;
  assign n2630 = ~n998 & n1002;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = ~n2627 & n2631;
  assign n2633 = ~n2625 & n2632;
  assign n2634 = ~n2623 & n2633;
  assign n2635 = ~n2621 & n2634;
  assign n2636 = ~n2619 & n2635;
  assign n2637 = ~n2617 & n2636;
  assign n2638 = ~n2614 & n2637;
  assign n2639 = ~n2612 & n2638;
  assign n2640 = ~n2608 & n2639;
  assign n2641 = ~\data<23>  & ~n2640;
  assign n2642 = \data<23>  & n2640;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = ~n504 & ~n2643;
  assign n2645 = \data_in<4>  & n504;
  assign \data_new<55>  = n2644 | n2645;
  assign n2647 = ~n810 & ~n814;
  assign n2648 = ~n811 & n2647;
  assign n2649 = ~n809 & n2648;
  assign n2650 = n789 & n2649;
  assign n2651 = ~n795 & n803;
  assign n2652 = n807 & n2651;
  assign n2653 = n797 & n805;
  assign n2654 = n809 & n2653;
  assign n2655 = ~n788 & n795;
  assign n2656 = n809 & n2655;
  assign n2657 = n804 & n813;
  assign n2658 = n810 & n2657;
  assign n2659 = n800 & ~n813;
  assign n2660 = n810 & n2659;
  assign n2661 = n792 & ~n813;
  assign n2662 = n804 & n2661;
  assign n2663 = n792 & n805;
  assign n2664 = ~n804 & n2663;
  assign n2665 = n814 & n1766;
  assign n2666 = n788 & n1765;
  assign n2667 = n806 & n1767;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n2665 & n2668;
  assign n2670 = ~n2664 & n2669;
  assign n2671 = ~n2662 & n2670;
  assign n2672 = ~n2660 & n2671;
  assign n2673 = ~n2658 & n2672;
  assign n2674 = ~n2656 & n2673;
  assign n2675 = ~n2654 & n2674;
  assign n2676 = ~n2652 & n2675;
  assign n2677 = ~n2650 & n2676;
  assign n2678 = ~\data<24>  & ~n2677;
  assign n2679 = \data<24>  & n2677;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = ~n504 & ~n2680;
  assign n2682 = \inreg<54>  & n504;
  assign \data_new<56>  = n2681 | n2682;
  assign n2684 = \D<6>  & n1986;
  assign n2685 = \D<8>  & n1988;
  assign n2686 = \D<9>  & n1989;
  assign n2687 = \D<5>  & n1990;
  assign n2688 = \D<7>  & n1991;
  assign n2689 = \inreg<53>  & n1993;
  assign n2690 = \data_in<6>  & n1994;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = ~n2688 & n2691;
  assign n2693 = ~n2687 & n2692;
  assign n2694 = ~n2686 & n2693;
  assign n2695 = ~n2685 & n2694;
  assign \D_new<7>  = n2684 | ~n2695;
  assign n2697 = \C<5>  & n1986;
  assign n2698 = \C<7>  & n1988;
  assign n2699 = \C<8>  & n1989;
  assign n2700 = \C<4>  & n1990;
  assign n2701 = \C<6>  & n1991;
  assign n2702 = \data_in<0>  & n1993;
  assign n2703 = \inreg<0>  & n1994;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~n2701 & n2704;
  assign n2706 = ~n2700 & n2705;
  assign n2707 = ~n2699 & n2706;
  assign n2708 = ~n2698 & n2707;
  assign \C_new<6>  = n2697 | ~n2708;
  assign n2710 = \D<7>  & n1986;
  assign n2711 = \D<9>  & n1988;
  assign n2712 = \D<10>  & n1989;
  assign n2713 = \D<6>  & n1990;
  assign n2714 = \D<8>  & n1991;
  assign n2715 = \inreg<45>  & n1993;
  assign n2716 = \inreg<53>  & n1994;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = ~n2714 & n2717;
  assign n2719 = ~n2713 & n2718;
  assign n2720 = ~n2712 & n2719;
  assign n2721 = ~n2711 & n2720;
  assign \D_new<8>  = n2710 | ~n2721;
  assign n2723 = \C<4>  & n1986;
  assign n2724 = \C<6>  & n1988;
  assign n2725 = \C<7>  & n1989;
  assign n2726 = \C<3>  & n1990;
  assign n2727 = \C<5>  & n1991;
  assign n2728 = \inreg<0>  & n1993;
  assign n2729 = \inreg<8>  & n1994;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2727 & n2730;
  assign n2732 = ~n2726 & n2731;
  assign n2733 = ~n2725 & n2732;
  assign n2734 = ~n2724 & n2733;
  assign \C_new<5>  = n2723 | ~n2734;
  assign n2736 = \D<4>  & n1986;
  assign n2737 = \D<6>  & n1988;
  assign n2738 = \D<7>  & n1989;
  assign n2739 = \D<3>  & n1990;
  assign n2740 = \D<5>  & n1991;
  assign n2741 = \inreg<6>  & n1993;
  assign n2742 = \inreg<14>  & n1994;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~n2740 & n2743;
  assign n2745 = ~n2739 & n2744;
  assign n2746 = ~n2738 & n2745;
  assign n2747 = ~n2737 & n2746;
  assign \D_new<5>  = n2736 | ~n2747;
  assign n2749 = \C<7>  & n1986;
  assign n2750 = \C<9>  & n1988;
  assign n2751 = \C<10>  & n1989;
  assign n2752 = \C<6>  & n1990;
  assign n2753 = \C<8>  & n1991;
  assign n2754 = \inreg<41>  & n1993;
  assign n2755 = \inreg<49>  & n1994;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = ~n2753 & n2756;
  assign n2758 = ~n2752 & n2757;
  assign n2759 = ~n2751 & n2758;
  assign n2760 = ~n2750 & n2759;
  assign \C_new<8>  = n2749 | ~n2760;
  assign n2762 = \D<5>  & n1986;
  assign n2763 = \D<7>  & n1988;
  assign n2764 = \D<8>  & n1989;
  assign n2765 = \D<4>  & n1990;
  assign n2766 = \D<6>  & n1991;
  assign n2767 = \data_in<6>  & n1993;
  assign n2768 = \inreg<6>  & n1994;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2766 & n2769;
  assign n2771 = ~n2765 & n2770;
  assign n2772 = ~n2764 & n2771;
  assign n2773 = ~n2763 & n2772;
  assign \D_new<6>  = n2762 | ~n2773;
  assign n2775 = \C<6>  & n1986;
  assign n2776 = \C<8>  & n1988;
  assign n2777 = \C<9>  & n1989;
  assign n2778 = \C<5>  & n1990;
  assign n2779 = \C<7>  & n1991;
  assign n2780 = \inreg<49>  & n1993;
  assign n2781 = \data_in<0>  & n1994;
  assign n2782 = ~n2780 & ~n2781;
  assign n2783 = ~n2779 & n2782;
  assign n2784 = ~n2778 & n2783;
  assign n2785 = ~n2777 & n2784;
  assign n2786 = ~n2776 & n2785;
  assign \C_new<7>  = n2775 | ~n2786;
  assign n2788 = \C<8>  & n1986;
  assign n2789 = \C<10>  & n1988;
  assign n2790 = \C<11>  & n1989;
  assign n2791 = \C<7>  & n1990;
  assign n2792 = \C<9>  & n1991;
  assign n2793 = \inreg<33>  & n1993;
  assign n2794 = \inreg<41>  & n1994;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2792 & n2795;
  assign n2797 = ~n2791 & n2796;
  assign n2798 = ~n2790 & n2797;
  assign n2799 = ~n2789 & n2798;
  assign \C_new<9>  = n2788 | ~n2799;
  assign n2801 = \D<8>  & n1986;
  assign n2802 = \D<10>  & n1988;
  assign n2803 = \D<11>  & n1989;
  assign n2804 = \D<7>  & n1990;
  assign n2805 = \D<9>  & n1991;
  assign n2806 = \inreg<37>  & n1993;
  assign n2807 = \inreg<45>  & n1994;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = ~n2805 & n2808;
  assign n2810 = ~n2804 & n2809;
  assign n2811 = ~n2803 & n2810;
  assign n2812 = ~n2802 & n2811;
  assign \D_new<9>  = n2801 | ~n2812;
  assign n2814 = \D<27>  & n1986;
  assign n2815 = \D<1>  & n1988;
  assign n2816 = \D<2>  & n1989;
  assign n2817 = \D<26>  & n1990;
  assign n2818 = \D<0>  & n1991;
  assign n2819 = \inreg<46>  & n1993;
  assign n2820 = \inreg<54>  & n1994;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2818 & n2821;
  assign n2823 = ~n2817 & n2822;
  assign n2824 = ~n2816 & n2823;
  assign n2825 = ~n2815 & n2824;
  assign \D_new<0>  = n2814 | ~n2825;
  assign n2827 = \C<27>  & n1986;
  assign n2828 = \C<1>  & n1988;
  assign n2829 = \C<2>  & n1989;
  assign n2830 = \C<26>  & n1990;
  assign n2831 = \C<0>  & n1991;
  assign n2832 = \inreg<40>  & n1993;
  assign n2833 = \inreg<48>  & n1994;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = ~n2831 & n2834;
  assign n2836 = ~n2830 & n2835;
  assign n2837 = ~n2829 & n2836;
  assign n2838 = ~n2828 & n2837;
  assign \C_new<0>  = n2827 | ~n2838;
  assign n2840 = \D<2>  & n1986;
  assign n2841 = \D<4>  & n1988;
  assign n2842 = \D<5>  & n1989;
  assign n2843 = \D<1>  & n1990;
  assign n2844 = \D<3>  & n1991;
  assign n2845 = \inreg<22>  & n1993;
  assign n2846 = \inreg<30>  & n1994;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = ~n2844 & n2847;
  assign n2849 = ~n2843 & n2848;
  assign n2850 = ~n2842 & n2849;
  assign n2851 = ~n2841 & n2850;
  assign \D_new<3>  = n2840 | ~n2851;
  assign n2853 = \C<1>  & n1986;
  assign n2854 = \C<3>  & n1988;
  assign n2855 = \C<4>  & n1989;
  assign n2856 = \C<0>  & n1990;
  assign n2857 = \C<2>  & n1991;
  assign n2858 = \inreg<24>  & n1993;
  assign n2859 = \inreg<32>  & n1994;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = ~n2857 & n2860;
  assign n2862 = ~n2856 & n2861;
  assign n2863 = ~n2855 & n2862;
  assign n2864 = ~n2854 & n2863;
  assign \C_new<2>  = n2853 | ~n2864;
  assign n2866 = \D<3>  & n1986;
  assign n2867 = \D<5>  & n1988;
  assign n2868 = \D<6>  & n1989;
  assign n2869 = \D<2>  & n1990;
  assign n2870 = \D<4>  & n1991;
  assign n2871 = \inreg<14>  & n1993;
  assign n2872 = \inreg<22>  & n1994;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = ~n2870 & n2873;
  assign n2875 = ~n2869 & n2874;
  assign n2876 = ~n2868 & n2875;
  assign n2877 = ~n2867 & n2876;
  assign \D_new<4>  = n2866 | ~n2877;
  assign n2879 = \C<0>  & n1986;
  assign n2880 = \C<2>  & n1988;
  assign n2881 = \C<3>  & n1989;
  assign n2882 = \C<27>  & n1990;
  assign n2883 = \C<1>  & n1991;
  assign n2884 = \inreg<32>  & n1993;
  assign n2885 = \inreg<40>  & n1994;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = ~n2883 & n2886;
  assign n2888 = ~n2882 & n2887;
  assign n2889 = ~n2881 & n2888;
  assign n2890 = ~n2880 & n2889;
  assign \C_new<1>  = n2879 | ~n2890;
  assign n2892 = \D<0>  & n1986;
  assign n2893 = \D<2>  & n1988;
  assign n2894 = \D<3>  & n1989;
  assign n2895 = \D<27>  & n1990;
  assign n2896 = \D<1>  & n1991;
  assign n2897 = \inreg<38>  & n1993;
  assign n2898 = \inreg<46>  & n1994;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & n2899;
  assign n2901 = ~n2895 & n2900;
  assign n2902 = ~n2894 & n2901;
  assign n2903 = ~n2893 & n2902;
  assign \D_new<1>  = n2892 | ~n2903;
  assign n2905 = \C<3>  & n1986;
  assign n2906 = \C<5>  & n1988;
  assign n2907 = \C<6>  & n1989;
  assign n2908 = \C<2>  & n1990;
  assign n2909 = \C<4>  & n1991;
  assign n2910 = \inreg<8>  & n1993;
  assign n2911 = \inreg<16>  & n1994;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = ~n2909 & n2912;
  assign n2914 = ~n2908 & n2913;
  assign n2915 = ~n2907 & n2914;
  assign n2916 = ~n2906 & n2915;
  assign \C_new<4>  = n2905 | ~n2916;
  assign n2918 = \D<1>  & n1986;
  assign n2919 = \D<3>  & n1988;
  assign n2920 = \D<4>  & n1989;
  assign n2921 = \D<0>  & n1990;
  assign n2922 = \D<2>  & n1991;
  assign n2923 = \inreg<30>  & n1993;
  assign n2924 = \inreg<38>  & n1994;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = ~n2922 & n2925;
  assign n2927 = ~n2921 & n2926;
  assign n2928 = ~n2920 & n2927;
  assign n2929 = ~n2919 & n2928;
  assign \D_new<2>  = n2918 | ~n2929;
  assign n2931 = \C<2>  & n1986;
  assign n2932 = \C<4>  & n1988;
  assign n2933 = \C<5>  & n1989;
  assign n2934 = \C<1>  & n1990;
  assign n2935 = \C<3>  & n1991;
  assign n2936 = \inreg<16>  & n1993;
  assign n2937 = \inreg<24>  & n1994;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = ~n2935 & n2938;
  assign n2940 = ~n2934 & n2939;
  assign n2941 = ~n2933 & n2940;
  assign n2942 = ~n2932 & n2941;
  assign \C_new<3>  = n2931 | ~n2942;
  assign n2944 = \inreg<42>  & n508;
  assign n2945 = ~\count<0>  & \inreg<50> ;
  assign \inreg_new<50>  = n2944 | n2945;
  assign n2947 = \inreg<1>  & n508;
  assign n2948 = \inreg<9>  & ~\count<0> ;
  assign \inreg_new<9>  = n2947 | n2948;
  assign n2950 = \inreg<46>  & n508;
  assign n2951 = ~\count<0>  & \inreg<54> ;
  assign \inreg_new<54>  = n2950 | n2951;
  assign n2953 = \inreg<45>  & n508;
  assign n2954 = ~\count<0>  & \inreg<53> ;
  assign \inreg_new<53>  = n2953 | n2954;
  assign n2956 = \inreg<44>  & n508;
  assign n2957 = ~\count<0>  & \inreg<52> ;
  assign \inreg_new<52>  = n2956 | n2957;
  assign n2959 = \data_in<6>  & n508;
  assign n2960 = \inreg<6>  & ~\count<0> ;
  assign \inreg_new<6>  = n2959 | n2960;
  assign n2962 = \inreg<43>  & n508;
  assign n2963 = ~\count<0>  & \inreg<51> ;
  assign \inreg_new<51>  = n2962 | n2963;
  assign n2965 = \data_in<5>  & n508;
  assign n2966 = \inreg<5>  & ~\count<0> ;
  assign \inreg_new<5>  = n2965 | n2966;
  assign n2968 = \inreg<0>  & n508;
  assign n2969 = \inreg<8>  & ~\count<0> ;
  assign \inreg_new<8>  = n2968 | n2969;
  assign n2971 = \data_in<7>  & n508;
  assign n2972 = \inreg<7>  & ~\count<0> ;
  assign \inreg_new<7>  = n2971 | n2972;
  assign n2974 = \data_in<2>  & n508;
  assign n2975 = \inreg<2>  & ~\count<0> ;
  assign \inreg_new<2>  = n2974 | n2975;
  assign n2977 = \inreg<47>  & n508;
  assign n2978 = ~\count<0>  & \inreg<55> ;
  assign \inreg_new<55>  = n2977 | n2978;
  assign n2980 = \data_in<1>  & n508;
  assign n2981 = \inreg<1>  & ~\count<0> ;
  assign \inreg_new<1>  = n2980 | n2981;
  assign n2983 = \data_in<4>  & n508;
  assign n2984 = \inreg<4>  & ~\count<0> ;
  assign \inreg_new<4>  = n2983 | n2984;
  assign n2986 = \data_in<3>  & n508;
  assign n2987 = \inreg<3>  & ~\count<0> ;
  assign \inreg_new<3>  = n2986 | n2987;
  assign n2989 = \data_in<0>  & n508;
  assign n2990 = \inreg<0>  & ~\count<0> ;
  assign \inreg_new<0>  = n2989 | n2990;
  assign n2992 = \encrypt_mode<0>  & n1983;
  assign n2993 = \encrypt<0>  & ~n1983;
  assign \encrypt_mode_new<0>  = n2992 | n2993;
  assign n2995 = ~n1098 & ~n1125;
  assign n2996 = ~n1112 & n2995;
  assign n2997 = n1108 & n2996;
  assign n2998 = ~n1173 & n2997;
  assign n2999 = ~n1098 & n1112;
  assign n3000 = n1115 & n2999;
  assign n3001 = n1126 & n3000;
  assign n3002 = ~n1101 & n1108;
  assign n3003 = n1114 & n3002;
  assign n3004 = n1129 & n3003;
  assign n3005 = n1111 & n1136;
  assign n3006 = ~n1108 & n3005;
  assign n3007 = ~n1135 & n3006;
  assign n3008 = n1101 & ~n1114;
  assign n3009 = n1131 & n3008;
  assign n3010 = ~n1113 & n3009;
  assign n3011 = n1098 & ~n1125;
  assign n3012 = n1115 & n3011;
  assign n3013 = ~n1113 & n3012;
  assign n3014 = ~n1098 & ~n1112;
  assign n3015 = n1128 & n3014;
  assign n3016 = ~n1115 & n1125;
  assign n3017 = n1134 & n3016;
  assign n3018 = ~n1107 & n1113;
  assign n3019 = n1126 & n3018;
  assign n3020 = ~n1129 & n2324;
  assign n3021 = n1135 & ~n2325;
  assign n3022 = n1129 & n3021;
  assign n3023 = n1108 & n1137;
  assign n3024 = n1130 & n1171;
  assign n3025 = n1177 & ~n3024;
  assign n3026 = ~n3023 & n3025;
  assign n3027 = ~n3022 & n3026;
  assign n3028 = ~n3020 & n3027;
  assign n3029 = ~n3019 & n3028;
  assign n3030 = ~n3017 & n3029;
  assign n3031 = ~n3015 & n3030;
  assign n3032 = ~n3013 & n3031;
  assign n3033 = ~n3010 & n3032;
  assign n3034 = ~n3007 & n3033;
  assign n3035 = ~n3004 & n3034;
  assign n3036 = ~n3001 & n3035;
  assign n3037 = ~n2998 & n3036;
  assign n3038 = ~\data<6>  & ~n3037;
  assign n3039 = \data<6>  & n3037;
  assign n3040 = ~n3038 & ~n3039;
  assign n3041 = n504 & ~n3040;
  assign n3042 = \outreg<17>  & n508;
  assign n3043 = ~\count<0>  & \outreg<9> ;
  assign n3044 = ~n3042 & ~n3043;
  assign \outreg_new<9>  = n3041 | ~n3044;
  assign n3046 = ~n1679 & n1688;
  assign n3047 = n1669 & n1699;
  assign n3048 = n1690 & n1710;
  assign n3049 = ~n1668 & ~n1682;
  assign n3050 = n1712 & n3049;
  assign n3051 = ~n1668 & ~n1672;
  assign n3052 = n1689 & n3051;
  assign n3053 = n1690 & n1694;
  assign n3054 = ~n1672 & n1704;
  assign n3055 = n1700 & n3054;
  assign n3056 = n1669 & n1672;
  assign n3057 = n1702 & n3056;
  assign n3058 = n1672 & n1679;
  assign n3059 = n1702 & n3058;
  assign n3060 = n1691 & ~n2561;
  assign n3061 = n1688 & n3060;
  assign n3062 = ~n1682 & n1697;
  assign n3063 = ~n1672 & n1713;
  assign n3064 = n1698 & n2558;
  assign n3065 = ~n2559 & ~n3048;
  assign n3066 = ~n2560 & n3065;
  assign n3067 = ~n1706 & n3066;
  assign n3068 = ~n1687 & n3067;
  assign n3069 = ~n3047 & n3068;
  assign n3070 = ~n3064 & n3069;
  assign n3071 = n1700 & n3046;
  assign n3072 = n3070 & ~n3071;
  assign n3073 = ~n3063 & n3072;
  assign n3074 = ~n3062 & n3073;
  assign n3075 = ~n3061 & n3074;
  assign n3076 = ~n3059 & n3075;
  assign n3077 = ~n3057 & n3076;
  assign n3078 = ~n3055 & n3077;
  assign n3079 = ~n3053 & n3078;
  assign n3080 = ~n3052 & n3079;
  assign n3081 = ~n3050 & n3080;
  assign n3082 = ~\data<9>  & ~n3081;
  assign n3083 = \data<9>  & n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n504 & ~n3084;
  assign n3086 = \outreg<59>  & n508;
  assign n3087 = \outreg<51>  & ~\count<0> ;
  assign n3088 = ~n3086 & ~n3087;
  assign \outreg_new<51>  = n3085 | ~n3088;
  assign n3090 = \outreg<60>  & n508;
  assign n3091 = \outreg<52>  & ~\count<0> ;
  assign n3092 = \data<49>  & n504;
  assign n3093 = ~n3091 & ~n3092;
  assign \outreg_new<52>  = n3090 | ~n3093;
  assign n3095 = ~n1363 & n1367;
  assign n3096 = n1385 & n3095;
  assign n3097 = ~n1880 & n3096;
  assign n3098 = n1379 & n1414;
  assign n3099 = n1390 & n3098;
  assign n3100 = ~n1367 & ~n1382;
  assign n3101 = n1384 & n3100;
  assign n3102 = n1363 & ~n1367;
  assign n3103 = n1386 & n3102;
  assign n3104 = n1371 & ~n1437;
  assign n3105 = n1393 & n3104;
  assign n3106 = n1360 & n1379;
  assign n3107 = n1603 & n3106;
  assign n3108 = ~n1367 & ~n1437;
  assign n3109 = n1388 & n3108;
  assign n3110 = ~n1371 & n1386;
  assign n3111 = n1437 & n1601;
  assign n3112 = n1363 & n1602;
  assign n3113 = n1374 & n1383;
  assign n3114 = n1376 & n1388;
  assign n3115 = ~n1881 & ~n3114;
  assign n3116 = ~n3113 & n3115;
  assign n3117 = ~n3112 & n3116;
  assign n3118 = ~n3111 & n3117;
  assign n3119 = ~n3110 & n3118;
  assign n3120 = ~n3109 & n3119;
  assign n3121 = ~n3107 & n3120;
  assign n3122 = ~n3105 & n3121;
  assign n3123 = ~n3103 & n3122;
  assign n3124 = ~n3101 & n3123;
  assign n3125 = ~n3099 & n3124;
  assign n3126 = ~n3097 & n3125;
  assign n3127 = ~\data<17>  & ~n3126;
  assign n3128 = \data<17>  & n3126;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n504 & ~n3129;
  assign n3131 = \outreg<61>  & n508;
  assign n3132 = \outreg<53>  & ~\count<0> ;
  assign n3133 = ~n3131 & ~n3132;
  assign \outreg_new<53>  = n3130 | ~n3133;
  assign n3135 = n504 & ~n2643;
  assign n3136 = \outreg<13>  & n508;
  assign n3137 = ~\count<0>  & \outreg<5> ;
  assign n3138 = ~n3136 & ~n3137;
  assign \outreg_new<5>  = n3135 | ~n3138;
  assign n3140 = \outreg<62>  & n508;
  assign n3141 = \outreg<54>  & ~\count<0> ;
  assign n3142 = \data<57>  & n504;
  assign n3143 = ~n3141 & ~n3142;
  assign \outreg_new<54>  = n3140 | ~n3143;
  assign n3145 = \outreg<14>  & n508;
  assign n3146 = ~\count<0>  & \outreg<6> ;
  assign n3147 = \data<63>  & n504;
  assign n3148 = ~n3146 & ~n3147;
  assign \outreg_new<6>  = n3145 | ~n3148;
  assign n3150 = n504 & ~n2358;
  assign n3151 = \outreg<15>  & n508;
  assign n3152 = ~\count<0>  & \outreg<7> ;
  assign n3153 = ~n3151 & ~n3152;
  assign \outreg_new<7>  = n3150 | ~n3153;
  assign n3155 = \outreg<16>  & n508;
  assign n3156 = ~\count<0>  & \outreg<8> ;
  assign n3157 = \data<38>  & n504;
  assign n3158 = ~n3156 & ~n3157;
  assign \outreg_new<8>  = n3155 | ~n3158;
  assign n3160 = n789 & n804;
  assign n3161 = n804 & n805;
  assign n3162 = ~n804 & ~n805;
  assign n3163 = n810 & n3162;
  assign n3164 = ~n807 & n3163;
  assign n3165 = ~n1766 & n3164;
  assign n3166 = n792 & n1799;
  assign n3167 = ~n789 & n3166;
  assign n3168 = ~n806 & n3167;
  assign n3169 = ~n1764 & n3168;
  assign n3170 = ~n792 & ~n803;
  assign n3171 = n789 & n3170;
  assign n3172 = ~n1767 & n3171;
  assign n3173 = ~n803 & ~n1799;
  assign n3174 = n795 & n3173;
  assign n3175 = n807 & n3174;
  assign n3176 = n1766 & n2647;
  assign n3177 = n785 & ~n3160;
  assign n3178 = n1767 & n3177;
  assign n3179 = n796 & n811;
  assign n3180 = n789 & n3179;
  assign n3181 = n804 & n814;
  assign n3182 = ~n807 & n3181;
  assign n3183 = ~n785 & ~n795;
  assign n3184 = n808 & n3183;
  assign n3185 = ~n788 & n1764;
  assign n3186 = ~n3161 & ~n3185;
  assign n3187 = ~n3184 & n3186;
  assign n3188 = ~n3182 & n3187;
  assign n3189 = ~n3180 & n3188;
  assign n3190 = ~n3178 & n3189;
  assign n3191 = ~n3176 & n3190;
  assign n3192 = ~n3175 & n3191;
  assign n3193 = ~n3172 & n3192;
  assign n3194 = ~n3169 & n3193;
  assign n3195 = ~n3165 & n3194;
  assign n3196 = ~\data<7>  & ~n3195;
  assign n3197 = \data<7>  & n3195;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = n504 & ~n3198;
  assign n3200 = \outreg<9>  & n508;
  assign n3201 = ~\count<0>  & \outreg<1> ;
  assign n3202 = ~n3200 & ~n3201;
  assign \outreg_new<1>  = n3199 | ~n3202;
  assign n3204 = \outreg<58>  & n508;
  assign n3205 = \outreg<50>  & ~\count<0> ;
  assign n3206 = \data<41>  & n504;
  assign n3207 = ~n3205 & ~n3206;
  assign \outreg_new<50>  = n3204 | ~n3207;
  assign n3209 = \outreg<10>  & n508;
  assign n3210 = ~\count<0>  & \outreg<2> ;
  assign n3211 = \data<47>  & n504;
  assign n3212 = ~n3210 & ~n3211;
  assign \outreg_new<2>  = n3209 | ~n3212;
  assign n3214 = ~\data<8>  & ~n918;
  assign n3215 = \data<8>  & n918;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = n504 & ~n3216;
  assign n3218 = \outreg<59>  & ~\count<0> ;
  assign \outreg_new<59>  = n3217 | n3218;
  assign n3220 = n1020 & ~n2604;
  assign n3221 = ~n993 & n3220;
  assign n3222 = n991 & ~n1001;
  assign n3223 = n998 & n3222;
  assign n3224 = ~n1004 & n3223;
  assign n3225 = n973 & n999;
  assign n3226 = ~n987 & n3225;
  assign n3227 = ~n1004 & n3226;
  assign n3228 = n990 & n1005;
  assign n3229 = n978 & n3228;
  assign n3230 = n1001 & n1003;
  assign n3231 = n998 & n3230;
  assign n3232 = n991 & n1001;
  assign n3233 = ~n998 & n3232;
  assign n3234 = n995 & n1003;
  assign n3235 = ~n1001 & n3234;
  assign n3236 = n980 & n986;
  assign n3237 = n1002 & n3236;
  assign n3238 = n993 & n999;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3235 & n3239;
  assign n3241 = ~n3233 & n3240;
  assign n3242 = ~n3231 & n3241;
  assign n3243 = ~n3229 & n3242;
  assign n3244 = ~n3227 & n3243;
  assign n3245 = ~n3224 & n3244;
  assign n3246 = ~n3221 & n3245;
  assign n3247 = ~\data<15>  & ~n3246;
  assign n3248 = \data<15>  & n3246;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = n504 & ~n3249;
  assign n3251 = \outreg<11>  & n508;
  assign n3252 = ~\count<0>  & \outreg<3> ;
  assign n3253 = ~n3251 & ~n3252;
  assign \outreg_new<3>  = n3250 | ~n3253;
  assign n3255 = \outreg<12>  & n508;
  assign n3256 = ~\count<0>  & \outreg<4> ;
  assign n3257 = \data<55>  & n504;
  assign n3258 = ~n3256 & ~n3257;
  assign \outreg_new<4>  = n3255 | ~n3258;
  assign n3260 = n504 & ~n2597;
  assign n3261 = \outreg<63>  & n508;
  assign n3262 = \outreg<55>  & ~\count<0> ;
  assign n3263 = ~n3261 & ~n3262;
  assign \outreg_new<55>  = n3260 | ~n3263;
  assign n3265 = ~n504 & ~n1652;
  assign n3266 = \inreg<26>  & n504;
  assign \data_new<43>  = n3265 | n3266;
  assign n3268 = \outreg<56>  & ~\count<0> ;
  assign n3269 = \data<32>  & n504;
  assign \outreg_new<56>  = n3268 | n3269;
  assign n3271 = ~n504 & ~n1440;
  assign n3272 = \inreg<18>  & n504;
  assign \data_new<44>  = n3271 | n3272;
  assign n3274 = \outreg<8>  & n508;
  assign n3275 = ~\count<0>  & \outreg<0> ;
  assign n3276 = \data<39>  & n504;
  assign n3277 = ~n3275 & ~n3276;
  assign \outreg_new<0>  = n3274 | ~n3277;
  assign n3279 = n1702 & n2578;
  assign n3280 = ~n1679 & n1702;
  assign n3281 = n2558 & n3280;
  assign n3282 = n1665 & n1679;
  assign n3283 = n1698 & n3282;
  assign n3284 = ~n1672 & n1688;
  assign n3285 = n1703 & n3284;
  assign n3286 = n1669 & n1675;
  assign n3287 = n1704 & n3286;
  assign n3288 = n1682 & n1697;
  assign n3289 = ~n1672 & n1686;
  assign n3290 = n1696 & n3046;
  assign n3291 = n1684 & n1685;
  assign n3292 = n1690 & n3046;
  assign n3293 = n1689 & n1691;
  assign n3294 = n1701 & n1704;
  assign n3295 = n1692 & n1693;
  assign n3296 = n1693 & n1703;
  assign n3297 = n1668 & n1698;
  assign n3298 = ~n1714 & ~n3048;
  assign n3299 = ~n3279 & n3298;
  assign n3300 = ~n1709 & n3299;
  assign n3301 = ~n3047 & n3300;
  assign n3302 = ~n3297 & n3301;
  assign n3303 = ~n3296 & n3302;
  assign n3304 = ~n3295 & n3303;
  assign n3305 = ~n3294 & n3304;
  assign n3306 = ~n3293 & n3305;
  assign n3307 = ~n3292 & n3306;
  assign n3308 = ~n3291 & n3307;
  assign n3309 = ~n3290 & n3308;
  assign n3310 = ~n3289 & n3309;
  assign n3311 = ~n3288 & n3310;
  assign n3312 = ~n3287 & n3311;
  assign n3313 = ~n3285 & n3312;
  assign n3314 = ~n3283 & n3313;
  assign n3315 = ~n3281 & n3314;
  assign n3316 = ~\data<0>  & ~n3315;
  assign n3317 = \data<0>  & n3315;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = n504 & ~n3318;
  assign n3320 = \outreg<57>  & ~\count<0> ;
  assign \outreg_new<57>  = n3319 | n3320;
  assign n3322 = ~n504 & ~n3084;
  assign n3323 = \inreg<42>  & n504;
  assign \data_new<41>  = n3322 | n3323;
  assign n3325 = \outreg<58>  & ~\count<0> ;
  assign n3326 = \data<40>  & n504;
  assign \outreg_new<58>  = n3325 | n3326;
  assign n3328 = ~n504 & ~n1863;
  assign n3329 = \inreg<34>  & n504;
  assign \data_new<42>  = n3328 | n3329;
  assign n3331 = \inreg<12>  & n508;
  assign n3332 = ~\count<0>  & \inreg<20> ;
  assign \inreg_new<20>  = n3331 | n3332;
  assign n3334 = n677 & n682;
  assign n3335 = n687 & n3334;
  assign n3336 = n660 & ~n673;
  assign n3337 = n668 & n3336;
  assign n3338 = ~n685 & n3337;
  assign n3339 = n676 & n680;
  assign n3340 = n678 & n3339;
  assign n3341 = n667 & n684;
  assign n3342 = n661 & n3341;
  assign n3343 = n669 & n681;
  assign n3344 = ~n668 & n3343;
  assign n3345 = n657 & n723;
  assign n3346 = n687 & n3345;
  assign n3347 = n670 & ~n673;
  assign n3348 = n669 & n3347;
  assign n3349 = ~n660 & n677;
  assign n3350 = n670 & n3349;
  assign n3351 = n657 & n667;
  assign n3352 = n677 & n3351;
  assign n3353 = ~n657 & n667;
  assign n3354 = n681 & n3353;
  assign n3355 = n680 & n685;
  assign n3356 = n676 & n683;
  assign n3357 = n688 & n723;
  assign n3358 = ~n676 & n883;
  assign n3359 = ~n3335 & ~n3358;
  assign n3360 = ~n3357 & n3359;
  assign n3361 = ~n3356 & n3360;
  assign n3362 = ~n3355 & n3361;
  assign n3363 = ~n3354 & n3362;
  assign n3364 = ~n3352 & n3363;
  assign n3365 = ~n3350 & n3364;
  assign n3366 = ~n3348 & n3365;
  assign n3367 = ~n3346 & n3366;
  assign n3368 = ~n3344 & n3367;
  assign n3369 = ~n3342 & n3368;
  assign n3370 = ~n3340 & n3369;
  assign n3371 = ~n3338 & n3370;
  assign n3372 = ~\data<16>  & ~n3371;
  assign n3373 = \data<16>  & n3371;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = n504 & ~n3374;
  assign n3376 = \outreg<61>  & ~\count<0> ;
  assign \outreg_new<61>  = n3375 | n3376;
  assign n3378 = \outreg<62>  & ~\count<0> ;
  assign n3379 = \data<56>  & n504;
  assign \outreg_new<62>  = n3378 | n3379;
  assign n3381 = ~n504 & ~n3216;
  assign n3382 = \inreg<50>  & n504;
  assign \data_new<40>  = n3381 | n3382;
  assign n3384 = n504 & ~n2680;
  assign n3385 = \outreg<63>  & ~\count<0> ;
  assign \outreg_new<63>  = n3384 | n3385;
  assign n3387 = \inreg<16>  & n508;
  assign n3388 = ~\count<0>  & \inreg<24> ;
  assign \inreg_new<24>  = n3387 | n3388;
  assign n3390 = \inreg<15>  & n508;
  assign n3391 = ~\count<0>  & \inreg<23> ;
  assign \inreg_new<23>  = n3390 | n3391;
  assign n3393 = \inreg<14>  & n508;
  assign n3394 = ~\count<0>  & \inreg<22> ;
  assign \inreg_new<22>  = n3393 | n3394;
  assign n3396 = ~n504 & ~n3129;
  assign n3397 = \inreg<44>  & n504;
  assign \data_new<49>  = n3396 | n3397;
  assign n3399 = \inreg<13>  & n508;
  assign n3400 = ~\count<0>  & \inreg<21> ;
  assign \inreg_new<21>  = n3399 | n3400;
  assign n3402 = \outreg<60>  & ~\count<0> ;
  assign n3403 = \data<48>  & n504;
  assign \outreg_new<60>  = n3402 | n3403;
  assign n3405 = \inreg<20>  & n508;
  assign n3406 = ~\count<0>  & \inreg<28> ;
  assign \inreg_new<28>  = n3405 | n3406;
  assign n3408 = ~n504 & ~n3249;
  assign n3409 = \data_in<2>  & n504;
  assign \data_new<47>  = n3408 | n3409;
  assign n3411 = \inreg<19>  & n508;
  assign n3412 = ~\count<0>  & \inreg<27> ;
  assign \inreg_new<27>  = n3411 | n3412;
  assign n3414 = ~n504 & ~n3374;
  assign n3415 = \inreg<52>  & n504;
  assign \data_new<48>  = n3414 | n3415;
  assign n3417 = \inreg<18>  & n508;
  assign n3418 = ~\count<0>  & \inreg<26> ;
  assign \inreg_new<26>  = n3417 | n3418;
  assign n3420 = ~n504 & ~n856;
  assign n3421 = \inreg<10>  & n504;
  assign \data_new<45>  = n3420 | n3421;
  assign n3423 = \inreg<17>  & n508;
  assign n3424 = ~\count<0>  & \inreg<25> ;
  assign \inreg_new<25>  = n3423 | n3424;
  assign n3426 = ~n504 & ~n638;
  assign n3427 = \inreg<2>  & n504;
  assign \data_new<46>  = n3426 | n3427;
  assign n3429 = ~n504 & ~n1919;
  assign n3430 = \inreg<40>  & n504;
  assign \data_new<33>  = n3429 | n3430;
  assign n3432 = ~n504 & ~n1802;
  assign n3433 = \inreg<32>  & n504;
  assign \data_new<34>  = n3432 | n3433;
  assign n3435 = \data_in<7>  & n504;
  assign n3436 = \data<63>  & ~n504;
  assign \data_new<31>  = n3435 | n3436;
  assign n3438 = \inreg<21>  & n508;
  assign n3439 = ~\count<0>  & \inreg<29> ;
  assign \inreg_new<29>  = n3438 | n3439;
  assign n3441 = ~n504 & ~n3318;
  assign n3442 = \inreg<48>  & n504;
  assign \data_new<32>  = n3441 | n3442;
  assign n3444 = \inreg<2>  & n508;
  assign n3445 = ~\count<0>  & \inreg<10> ;
  assign \inreg_new<10>  = n3444 | n3445;
  assign n3447 = \inreg<7>  & n504;
  assign n3448 = \data<62>  & ~n504;
  assign \data_new<30>  = n3447 | n3448;
  assign n3450 = \inreg<6>  & n508;
  assign n3451 = ~\count<0>  & \inreg<14> ;
  assign \inreg_new<14>  = n3450 | n3451;
  assign n3453 = \inreg<5>  & n508;
  assign n3454 = ~\count<0>  & \inreg<13> ;
  assign \inreg_new<13>  = n3453 | n3454;
  assign n3456 = \inreg<4>  & n508;
  assign n3457 = ~\count<0>  & \inreg<12> ;
  assign \inreg_new<12>  = n3456 | n3457;
  assign n3459 = ~n504 & ~n3198;
  assign n3460 = \data_in<0>  & n504;
  assign \data_new<39>  = n3459 | n3460;
  assign n3462 = \inreg<3>  & n508;
  assign n3463 = ~\count<0>  & \inreg<11> ;
  assign \inreg_new<11>  = n3462 | n3463;
  assign n3465 = \inreg<10>  & n508;
  assign n3466 = ~\count<0>  & \inreg<18> ;
  assign \inreg_new<18>  = n3465 | n3466;
  assign n3468 = ~n504 & ~n1082;
  assign n3469 = \inreg<8>  & n504;
  assign \data_new<37>  = n3468 | n3469;
  assign n3471 = \inreg<9>  & n508;
  assign n3472 = ~\count<0>  & \inreg<17> ;
  assign \inreg_new<17>  = n3471 | n3472;
  assign n3474 = ~n504 & ~n3040;
  assign n3475 = \inreg<0>  & n504;
  assign \data_new<38>  = n3474 | n3475;
  assign n3477 = \inreg<8>  & n508;
  assign n3478 = ~\count<0>  & \inreg<16> ;
  assign \inreg_new<16>  = n3477 | n3478;
  assign n3480 = ~n504 & ~n1585;
  assign n3481 = \inreg<24>  & n504;
  assign \data_new<35>  = n3480 | n3481;
  assign n3483 = \inreg<7>  & n508;
  assign n3484 = ~\count<0>  & \inreg<15> ;
  assign \inreg_new<15>  = n3483 | n3484;
  assign n3486 = ~n504 & ~n1347;
  assign n3487 = \inreg<16>  & n504;
  assign \data_new<36>  = n3486 | n3487;
  assign n3489 = \data_in<5>  & n504;
  assign n3490 = \data<55>  & ~n504;
  assign \data_new<23>  = n3489 | n3490;
  assign n3492 = \inreg<55>  & n504;
  assign n3493 = \data<56>  & ~n504;
  assign \data_new<24>  = n3492 | n3493;
  assign n3495 = \inreg<13>  & n504;
  assign n3496 = \data<53>  & ~n504;
  assign \data_new<21>  = n3495 | n3496;
  assign n3498 = \inreg<11>  & n508;
  assign n3499 = ~\count<0>  & \inreg<19> ;
  assign \inreg_new<19>  = n3498 | n3499;
  assign n3501 = \inreg<5>  & n504;
  assign n3502 = \data<54>  & ~n504;
  assign \data_new<22>  = n3501 | n3502;
  assign n3504 = \inreg<32>  & n508;
  assign n3505 = ~\count<0>  & \inreg<40> ;
  assign \inreg_new<40>  = n3504 | n3505;
  assign n3507 = \inreg<21>  & n504;
  assign n3508 = \data<52>  & ~n504;
  assign \data_new<20>  = n3507 | n3508;
  assign n3510 = \inreg<36>  & n508;
  assign n3511 = ~\count<0>  & \inreg<44> ;
  assign \inreg_new<44>  = n3510 | n3511;
  assign n3513 = \inreg<35>  & n508;
  assign n3514 = ~\count<0>  & \inreg<43> ;
  assign \inreg_new<43>  = n3513 | n3514;
  assign n3516 = \inreg<34>  & n508;
  assign n3517 = ~\count<0>  & \inreg<42> ;
  assign \inreg_new<42>  = n3516 | n3517;
  assign n3519 = \inreg<15>  & n504;
  assign n3520 = \data<61>  & ~n504;
  assign \data_new<29>  = n3519 | n3520;
  assign n3522 = \inreg<33>  & n508;
  assign n3523 = ~\count<0>  & \inreg<41> ;
  assign \inreg_new<41>  = n3522 | n3523;
  assign n3525 = \inreg<40>  & n508;
  assign n3526 = ~\count<0>  & \inreg<48> ;
  assign \inreg_new<48>  = n3525 | n3526;
  assign n3528 = \inreg<31>  & n504;
  assign n3529 = \data<59>  & ~n504;
  assign \data_new<27>  = n3528 | n3529;
  assign n3531 = \inreg<39>  & n508;
  assign n3532 = ~\count<0>  & \inreg<47> ;
  assign \inreg_new<47>  = n3531 | n3532;
  assign n3534 = \inreg<23>  & n504;
  assign n3535 = \data<60>  & ~n504;
  assign \data_new<28>  = n3534 | n3535;
  assign n3537 = \inreg<38>  & n508;
  assign n3538 = ~\count<0>  & \inreg<46> ;
  assign \inreg_new<46>  = n3537 | n3538;
endmodule


