// Benchmark "i9" written by ABC on Tue May 16 16:07:51 2017

module i9 ( 
    \V88(11) , \V88(10) , \V88(17) , \V88(16) , \V88(19) , \V88(18) ,
    \V88(23) , \V56(0) , \V88(22) , \V56(13) , \V56(1) , \V88(25) ,
    \V56(12) , \V56(2) , \V88(24) , \V56(15) , \V56(3) , \V56(14) ,
    \V56(4) , \V56(5) , \V88(21) , \V56(6) , \V88(20) , \V56(11) ,
    \V56(7) , \V56(10) , \V56(8) , \V56(9) , \V88(27) , \V88(26) ,
    \V56(17) , \V88(29) , \V56(16) , \V88(28) , \V56(19) , \V56(18) ,
    \V56(23) , \V56(22) , \V24(13) , \V56(25) , \V24(12) , \V56(24) ,
    \V24(14) , \V88(31) , \V88(30) , \V56(21) , \V56(20) , \V24(11) ,
    \V24(10) , \V56(27) , \V56(26) , \V56(29) , \V56(28) , \V56(31) ,
    \V56(30) , \V24(0) , \V24(1) , \V24(2) , \V24(3) , \V24(4) , \V24(5) ,
    \V24(6) , \V24(7) , \V24(8) , \V24(9) , \V88(0) , \V88(1) , \V88(2) ,
    \V88(3) , \V88(4) , \V88(5) , \V88(6) , \V88(7) , \V88(8) , \V9(0) ,
    \V88(9) , \V9(1) , \V9(2) , \V9(3) , \V9(5) , \V9(6) , \V9(7) ,
    \V9(8) , \V9(10) , \V88(13) , \V88(12) , \V88(15) , \V88(14) ,
    \V119(30) , \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) ,
    \V151(0) , \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V119(3) ,
    \V119(2) , \V119(5) , \V119(4) , \V151(27) , \V151(26) , \V151(29) ,
    \V119(1) , \V151(28) , \V119(0) , \V119(7) , \V119(6) , \V151(21) ,
    \V119(9) , \V151(20) , \V119(8) , \V151(23) , \V151(22) , \V151(25) ,
    \V151(24) , \V151(17) , \V151(16) , \V151(19) , \V151(18) , \V151(11) ,
    \V151(10) , \V151(13) , \V151(12) , \V119(27) , \V151(15) , \V119(26) ,
    \V151(14) , \V119(29) , \V119(28) , \V119(21) , \V119(20) , \V119(23) ,
    \V119(22) , \V119(25) , \V119(24) , \V119(17) , \V119(16) , \V119(19) ,
    \V119(18) , \V119(11) , \V119(10) , \V119(13) , \V151(31) , \V119(12) ,
    \V151(30) , \V119(15) , \V119(14)   );
  input  \V88(11) , \V88(10) , \V88(17) , \V88(16) , \V88(19) ,
    \V88(18) , \V88(23) , \V56(0) , \V88(22) , \V56(13) , \V56(1) ,
    \V88(25) , \V56(12) , \V56(2) , \V88(24) , \V56(15) , \V56(3) ,
    \V56(14) , \V56(4) , \V56(5) , \V88(21) , \V56(6) , \V88(20) ,
    \V56(11) , \V56(7) , \V56(10) , \V56(8) , \V56(9) , \V88(27) ,
    \V88(26) , \V56(17) , \V88(29) , \V56(16) , \V88(28) , \V56(19) ,
    \V56(18) , \V56(23) , \V56(22) , \V24(13) , \V56(25) , \V24(12) ,
    \V56(24) , \V24(14) , \V88(31) , \V88(30) , \V56(21) , \V56(20) ,
    \V24(11) , \V24(10) , \V56(27) , \V56(26) , \V56(29) , \V56(28) ,
    \V56(31) , \V56(30) , \V24(0) , \V24(1) , \V24(2) , \V24(3) , \V24(4) ,
    \V24(5) , \V24(6) , \V24(7) , \V24(8) , \V24(9) , \V88(0) , \V88(1) ,
    \V88(2) , \V88(3) , \V88(4) , \V88(5) , \V88(6) , \V88(7) , \V88(8) ,
    \V9(0) , \V88(9) , \V9(1) , \V9(2) , \V9(3) , \V9(5) , \V9(6) ,
    \V9(7) , \V9(8) , \V9(10) , \V88(13) , \V88(12) , \V88(15) , \V88(14) ;
  output \V119(30) , \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) ,
    \V151(0) , \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V119(3) ,
    \V119(2) , \V119(5) , \V119(4) , \V151(27) , \V151(26) , \V151(29) ,
    \V119(1) , \V151(28) , \V119(0) , \V119(7) , \V119(6) , \V151(21) ,
    \V119(9) , \V151(20) , \V119(8) , \V151(23) , \V151(22) , \V151(25) ,
    \V151(24) , \V151(17) , \V151(16) , \V151(19) , \V151(18) , \V151(11) ,
    \V151(10) , \V151(13) , \V151(12) , \V119(27) , \V151(15) , \V119(26) ,
    \V151(14) , \V119(29) , \V119(28) , \V119(21) , \V119(20) , \V119(23) ,
    \V119(22) , \V119(25) , \V119(24) , \V119(17) , \V119(16) , \V119(19) ,
    \V119(18) , \V119(11) , \V119(10) , \V119(13) , \V151(31) , \V119(12) ,
    \V151(30) , \V119(15) , \V119(14) ;
  wire n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n216, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n636, n637,
    n638, n639, n640, n641, n642, n643, n645, n646, n647, n648, n649, n650,
    n651, n652, n654, n655, n656, n657, n658, n659, n660, n661, n662, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n696, n697, n698, n699, n700, n701, n702, n703,
    n705, n706, n707, n708, n709, n710, n711, n712, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n726, n727, n728, n729, n730,
    n731, n732, n733, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n747, n748, n749, n750, n751, n752, n753, n754, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996;
  assign n152 = ~\V9(1)  & \V9(2) ;
  assign n153 = ~\V9(10)  & n152;
  assign n154 = \V9(8)  & n153;
  assign n155 = \V9(0)  & n153;
  assign n156 = ~\V9(5)  & n155;
  assign n157 = ~\V9(6)  & n156;
  assign n158 = \V9(1)  & ~\V9(3) ;
  assign n159 = \V9(2)  & n158;
  assign n160 = ~\V9(10)  & n159;
  assign n161 = \V9(1)  & ~\V9(10) ;
  assign n162 = \V9(8)  & n161;
  assign n163 = \V9(1)  & ~\V9(2) ;
  assign n164 = ~\V9(10)  & n163;
  assign n165 = ~\V9(5)  & n164;
  assign n166 = ~\V9(6)  & n165;
  assign n167 = ~\V9(0)  & ~\V9(10) ;
  assign n168 = ~\V9(5)  & n167;
  assign n169 = \V9(7)  & n167;
  assign n170 = \V9(1)  & \V9(3) ;
  assign n171 = \V9(2)  & n170;
  assign n172 = \V9(1)  & \V9(10) ;
  assign n173 = \V9(2)  & \V9(10) ;
  assign n174 = ~\V9(1)  & ~\V9(2) ;
  assign n175 = ~\V9(5)  & n174;
  assign n176 = ~\V9(6)  & n175;
  assign n177 = \V9(7)  & n174;
  assign n178 = \V9(10)  & n174;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n176 & n179;
  assign n181 = ~n173 & n180;
  assign n182 = ~n172 & n181;
  assign n183 = ~n171 & n182;
  assign n184 = ~n169 & n183;
  assign n185 = ~n168 & n184;
  assign n186 = ~n166 & n185;
  assign n187 = ~n162 & n186;
  assign n188 = ~n160 & n187;
  assign n189 = ~n157 & n188;
  assign n190 = ~n154 & n189;
  assign n191 = ~n154 & ~n157;
  assign n192 = ~n160 & n191;
  assign n193 = ~n177 & n192;
  assign n194 = ~n176 & n193;
  assign n195 = ~n178 & n194;
  assign n196 = ~n162 & ~n169;
  assign n197 = ~n168 & n196;
  assign n198 = ~n166 & n197;
  assign n199 = ~n177 & n198;
  assign n200 = ~n176 & n199;
  assign n201 = ~n178 & n200;
  assign n202 = \V56(16)  & ~n201;
  assign n203 = ~n195 & n202;
  assign n204 = ~n190 & n203;
  assign n205 = \V56(20)  & ~n190;
  assign n206 = ~n195 & n205;
  assign n207 = n201 & n206;
  assign n208 = ~n190 & n195;
  assign n209 = ~n201 & n208;
  assign n210 = \V56(23)  & n209;
  assign n211 = \V56(31)  & ~n190;
  assign n212 = n195 & n211;
  assign n213 = n201 & n212;
  assign n214 = ~n190 & ~n213;
  assign n215 = ~n210 & n214;
  assign n216 = ~n207 & n215;
  assign \V119(30)  = n204 | ~n216;
  assign n218 = \V56(20)  & ~n201;
  assign n219 = ~n195 & n218;
  assign n220 = ~n190 & n219;
  assign n221 = \V56(24)  & ~n190;
  assign n222 = ~n195 & n221;
  assign n223 = n201 & n222;
  assign n224 = \V56(27)  & ~n190;
  assign n225 = n195 & n224;
  assign n226 = ~n201 & n225;
  assign n227 = \V88(3)  & ~n190;
  assign n228 = n195 & n227;
  assign n229 = n201 & n228;
  assign n230 = n190 & ~n195;
  assign n231 = ~n201 & n230;
  assign n232 = n201 & n230;
  assign n233 = n190 & n195;
  assign n234 = ~n201 & n233;
  assign n235 = n201 & n233;
  assign n236 = ~n234 & ~n235;
  assign n237 = ~n232 & n236;
  assign n238 = ~n231 & n237;
  assign n239 = ~n229 & n238;
  assign n240 = ~n226 & n239;
  assign n241 = ~n223 & n240;
  assign \V151(3)  = n220 | ~n241;
  assign n243 = \V56(19)  & ~n201;
  assign n244 = ~n195 & n243;
  assign n245 = ~n190 & n244;
  assign n246 = \V56(23)  & ~n190;
  assign n247 = ~n195 & n246;
  assign n248 = n201 & n247;
  assign n249 = \V56(26)  & ~n190;
  assign n250 = n195 & n249;
  assign n251 = ~n201 & n250;
  assign n252 = \V88(2)  & ~n190;
  assign n253 = n195 & n252;
  assign n254 = n201 & n253;
  assign n255 = n238 & ~n254;
  assign n256 = ~n251 & n255;
  assign n257 = ~n248 & n256;
  assign \V151(2)  = n245 | ~n257;
  assign n259 = \V56(22)  & ~n201;
  assign n260 = ~n195 & n259;
  assign n261 = ~n190 & n260;
  assign n262 = ~n195 & n249;
  assign n263 = n201 & n262;
  assign n264 = \V56(29)  & ~n190;
  assign n265 = n195 & n264;
  assign n266 = ~n201 & n265;
  assign n267 = \V88(5)  & ~n190;
  assign n268 = n195 & n267;
  assign n269 = n201 & n268;
  assign n270 = n238 & ~n269;
  assign n271 = ~n266 & n270;
  assign n272 = ~n263 & n271;
  assign \V151(5)  = n261 | ~n272;
  assign n274 = \V56(21)  & ~n201;
  assign n275 = ~n195 & n274;
  assign n276 = ~n190 & n275;
  assign n277 = \V56(25)  & ~n190;
  assign n278 = ~n195 & n277;
  assign n279 = n201 & n278;
  assign n280 = \V56(28)  & ~n190;
  assign n281 = n195 & n280;
  assign n282 = ~n201 & n281;
  assign n283 = \V88(4)  & ~n190;
  assign n284 = n195 & n283;
  assign n285 = n201 & n284;
  assign n286 = n238 & ~n285;
  assign n287 = ~n282 & n286;
  assign n288 = ~n279 & n287;
  assign \V151(4)  = n276 | ~n288;
  assign n290 = \V56(18)  & ~n201;
  assign n291 = ~n195 & n290;
  assign n292 = ~n190 & n291;
  assign n293 = \V56(22)  & ~n190;
  assign n294 = ~n195 & n293;
  assign n295 = n201 & n294;
  assign n296 = n195 & n277;
  assign n297 = ~n201 & n296;
  assign n298 = \V88(1)  & ~n190;
  assign n299 = n195 & n298;
  assign n300 = n201 & n299;
  assign n301 = n238 & ~n300;
  assign n302 = ~n297 & n301;
  assign n303 = ~n295 & n302;
  assign \V151(1)  = n292 | ~n303;
  assign n305 = \V56(17)  & ~n201;
  assign n306 = ~n195 & n305;
  assign n307 = ~n190 & n306;
  assign n308 = \V56(21)  & ~n190;
  assign n309 = ~n195 & n308;
  assign n310 = n201 & n309;
  assign n311 = n195 & n221;
  assign n312 = ~n201 & n311;
  assign n313 = \V88(0)  & ~n190;
  assign n314 = n195 & n313;
  assign n315 = n201 & n314;
  assign n316 = n238 & ~n315;
  assign n317 = ~n312 & n316;
  assign n318 = ~n310 & n317;
  assign \V151(0)  = n307 | ~n318;
  assign n320 = \V56(24)  & ~n201;
  assign n321 = ~n195 & n320;
  assign n322 = ~n190 & n321;
  assign n323 = ~n195 & n280;
  assign n324 = n201 & n323;
  assign n325 = ~n201 & n212;
  assign n326 = \V88(7)  & ~n190;
  assign n327 = n195 & n326;
  assign n328 = n201 & n327;
  assign n329 = n238 & ~n328;
  assign n330 = ~n325 & n329;
  assign n331 = ~n324 & n330;
  assign \V151(7)  = n322 | ~n331;
  assign n333 = \V56(23)  & ~n201;
  assign n334 = ~n195 & n333;
  assign n335 = ~n190 & n334;
  assign n336 = ~n195 & n224;
  assign n337 = n201 & n336;
  assign n338 = \V56(30)  & ~n190;
  assign n339 = n195 & n338;
  assign n340 = ~n201 & n339;
  assign n341 = \V88(6)  & ~n190;
  assign n342 = n195 & n341;
  assign n343 = n201 & n342;
  assign n344 = n238 & ~n343;
  assign n345 = ~n340 & n344;
  assign n346 = ~n337 & n345;
  assign \V151(6)  = n335 | ~n346;
  assign n348 = \V56(26)  & ~n201;
  assign n349 = ~n195 & n348;
  assign n350 = ~n190 & n349;
  assign n351 = ~n195 & n338;
  assign n352 = n201 & n351;
  assign n353 = ~n201 & n299;
  assign n354 = \V88(9)  & ~n190;
  assign n355 = n195 & n354;
  assign n356 = n201 & n355;
  assign n357 = n238 & ~n356;
  assign n358 = ~n353 & n357;
  assign n359 = ~n352 & n358;
  assign \V151(9)  = n350 | ~n359;
  assign n361 = \V56(25)  & ~n201;
  assign n362 = ~n195 & n361;
  assign n363 = ~n190 & n362;
  assign n364 = ~n195 & n264;
  assign n365 = n201 & n364;
  assign n366 = ~n201 & n314;
  assign n367 = \V88(8)  & ~n190;
  assign n368 = n195 & n367;
  assign n369 = n201 & n368;
  assign n370 = n238 & ~n369;
  assign n371 = ~n366 & n370;
  assign n372 = ~n365 & n371;
  assign \V151(8)  = n363 | ~n372;
  assign n374 = \V24(3)  & ~n201;
  assign n375 = ~n195 & n374;
  assign n376 = ~n190 & n375;
  assign n377 = ~n195 & n283;
  assign n378 = n201 & n377;
  assign n379 = \V56(4)  & ~n190;
  assign n380 = n195 & n379;
  assign n381 = n201 & n380;
  assign n382 = ~n190 & ~n209;
  assign n383 = ~n381 & n382;
  assign n384 = ~n378 & n383;
  assign \V119(3)  = n376 | ~n384;
  assign n386 = \V24(2)  & ~n201;
  assign n387 = ~n195 & n386;
  assign n388 = ~n190 & n387;
  assign n389 = ~n195 & n227;
  assign n390 = n201 & n389;
  assign n391 = \V56(3)  & ~n190;
  assign n392 = n195 & n391;
  assign n393 = n201 & n392;
  assign n394 = n382 & ~n393;
  assign n395 = ~n390 & n394;
  assign \V119(2)  = n388 | ~n395;
  assign n397 = \V24(5)  & ~n201;
  assign n398 = ~n195 & n397;
  assign n399 = ~n190 & n398;
  assign n400 = ~n195 & n341;
  assign n401 = n201 & n400;
  assign n402 = \V56(6)  & ~n190;
  assign n403 = n195 & n402;
  assign n404 = n201 & n403;
  assign n405 = n382 & ~n404;
  assign n406 = ~n401 & n405;
  assign \V119(5)  = n399 | ~n406;
  assign n408 = \V24(4)  & ~n201;
  assign n409 = ~n195 & n408;
  assign n410 = ~n190 & n409;
  assign n411 = ~n195 & n267;
  assign n412 = n201 & n411;
  assign n413 = \V56(5)  & ~n190;
  assign n414 = n195 & n413;
  assign n415 = n201 & n414;
  assign n416 = n382 & ~n415;
  assign n417 = ~n412 & n416;
  assign \V119(4)  = n410 | ~n417;
  assign n419 = \V88(12)  & ~n201;
  assign n420 = ~n195 & n419;
  assign n421 = ~n190 & n420;
  assign n422 = \V88(16)  & ~n190;
  assign n423 = ~n195 & n422;
  assign n424 = n201 & n423;
  assign n425 = \V88(19)  & ~n190;
  assign n426 = n195 & n425;
  assign n427 = ~n201 & n426;
  assign n428 = \V88(27)  & ~n190;
  assign n429 = n195 & n428;
  assign n430 = n201 & n429;
  assign n431 = n238 & ~n430;
  assign n432 = ~n427 & n431;
  assign n433 = ~n424 & n432;
  assign \V151(27)  = n421 | ~n433;
  assign n435 = \V88(11)  & ~n201;
  assign n436 = ~n195 & n435;
  assign n437 = ~n190 & n436;
  assign n438 = \V88(15)  & ~n190;
  assign n439 = ~n195 & n438;
  assign n440 = n201 & n439;
  assign n441 = \V88(18)  & ~n190;
  assign n442 = n195 & n441;
  assign n443 = ~n201 & n442;
  assign n444 = \V88(26)  & ~n190;
  assign n445 = n195 & n444;
  assign n446 = n201 & n445;
  assign n447 = n238 & ~n446;
  assign n448 = ~n443 & n447;
  assign n449 = ~n440 & n448;
  assign \V151(26)  = n437 | ~n449;
  assign n451 = \V88(14)  & ~n201;
  assign n452 = ~n195 & n451;
  assign n453 = ~n190 & n452;
  assign n454 = ~n195 & n441;
  assign n455 = n201 & n454;
  assign n456 = \V88(21)  & ~n190;
  assign n457 = n195 & n456;
  assign n458 = ~n201 & n457;
  assign n459 = \V88(29)  & ~n190;
  assign n460 = n195 & n459;
  assign n461 = n201 & n460;
  assign n462 = n238 & ~n461;
  assign n463 = ~n458 & n462;
  assign n464 = ~n455 & n463;
  assign \V151(29)  = n453 | ~n464;
  assign n466 = \V24(1)  & ~n201;
  assign n467 = ~n195 & n466;
  assign n468 = ~n190 & n467;
  assign n469 = ~n195 & n252;
  assign n470 = n201 & n469;
  assign n471 = \V56(2)  & ~n190;
  assign n472 = n195 & n471;
  assign n473 = n201 & n472;
  assign n474 = n382 & ~n473;
  assign n475 = ~n470 & n474;
  assign \V119(1)  = n468 | ~n475;
  assign n477 = \V88(13)  & ~n201;
  assign n478 = ~n195 & n477;
  assign n479 = ~n190 & n478;
  assign n480 = \V88(17)  & ~n190;
  assign n481 = ~n195 & n480;
  assign n482 = n201 & n481;
  assign n483 = \V88(20)  & ~n190;
  assign n484 = n195 & n483;
  assign n485 = ~n201 & n484;
  assign n486 = \V88(28)  & ~n190;
  assign n487 = n195 & n486;
  assign n488 = n201 & n487;
  assign n489 = n238 & ~n488;
  assign n490 = ~n485 & n489;
  assign n491 = ~n482 & n490;
  assign \V151(28)  = n479 | ~n491;
  assign n493 = \V24(0)  & ~n201;
  assign n494 = ~n195 & n493;
  assign n495 = ~n190 & n494;
  assign n496 = ~n195 & n298;
  assign n497 = n201 & n496;
  assign n498 = \V56(1)  & ~n190;
  assign n499 = n195 & n498;
  assign n500 = n201 & n499;
  assign n501 = n382 & ~n500;
  assign n502 = ~n497 & n501;
  assign \V119(0)  = n495 | ~n502;
  assign n504 = \V24(7)  & ~n201;
  assign n505 = ~n195 & n504;
  assign n506 = ~n190 & n505;
  assign n507 = ~n195 & n367;
  assign n508 = n201 & n507;
  assign n509 = \V56(0)  & n209;
  assign n510 = \V56(8)  & ~n190;
  assign n511 = n195 & n510;
  assign n512 = n201 & n511;
  assign n513 = ~n190 & ~n512;
  assign n514 = ~n509 & n513;
  assign n515 = ~n508 & n514;
  assign \V119(7)  = n506 | ~n515;
  assign n517 = \V24(6)  & ~n201;
  assign n518 = ~n195 & n517;
  assign n519 = ~n190 & n518;
  assign n520 = ~n195 & n326;
  assign n521 = n201 & n520;
  assign n522 = \V56(7)  & ~n190;
  assign n523 = n195 & n522;
  assign n524 = n201 & n523;
  assign n525 = ~n190 & ~n524;
  assign n526 = ~n209 & n525;
  assign n527 = ~n521 & n526;
  assign \V119(6)  = n519 | ~n527;
  assign n529 = \V88(6)  & ~n201;
  assign n530 = ~n195 & n529;
  assign n531 = ~n190 & n530;
  assign n532 = \V88(10)  & ~n190;
  assign n533 = ~n195 & n532;
  assign n534 = n201 & n533;
  assign n535 = \V88(13)  & ~n190;
  assign n536 = n195 & n535;
  assign n537 = ~n201 & n536;
  assign n538 = n201 & n457;
  assign n539 = n238 & ~n538;
  assign n540 = ~n537 & n539;
  assign n541 = ~n534 & n540;
  assign \V151(21)  = n531 | ~n541;
  assign n543 = \V24(9)  & ~n201;
  assign n544 = ~n195 & n543;
  assign n545 = ~n190 & n544;
  assign n546 = \V56(2)  & n209;
  assign n547 = \V56(10)  & ~n190;
  assign n548 = n195 & n547;
  assign n549 = n201 & n548;
  assign n550 = ~n190 & ~n549;
  assign n551 = ~n546 & n550;
  assign n552 = ~n534 & n551;
  assign \V119(9)  = n545 | ~n552;
  assign n554 = \V88(5)  & ~n201;
  assign n555 = ~n195 & n554;
  assign n556 = ~n190 & n555;
  assign n557 = ~n195 & n354;
  assign n558 = n201 & n557;
  assign n559 = \V88(12)  & ~n190;
  assign n560 = n195 & n559;
  assign n561 = ~n201 & n560;
  assign n562 = n201 & n484;
  assign n563 = n238 & ~n562;
  assign n564 = ~n561 & n563;
  assign n565 = ~n558 & n564;
  assign \V151(20)  = n556 | ~n565;
  assign n567 = \V24(8)  & ~n201;
  assign n568 = ~n195 & n567;
  assign n569 = ~n190 & n568;
  assign n570 = \V56(1)  & n209;
  assign n571 = \V56(9)  & ~n190;
  assign n572 = n195 & n571;
  assign n573 = n201 & n572;
  assign n574 = ~n190 & ~n573;
  assign n575 = ~n570 & n574;
  assign n576 = ~n558 & n575;
  assign \V119(8)  = n569 | ~n576;
  assign n578 = \V88(8)  & ~n201;
  assign n579 = ~n195 & n578;
  assign n580 = ~n190 & n579;
  assign n581 = ~n195 & n559;
  assign n582 = n201 & n581;
  assign n583 = n195 & n438;
  assign n584 = ~n201 & n583;
  assign n585 = \V88(23)  & ~n190;
  assign n586 = n195 & n585;
  assign n587 = n201 & n586;
  assign n588 = n238 & ~n587;
  assign n589 = ~n584 & n588;
  assign n590 = ~n582 & n589;
  assign \V151(23)  = n580 | ~n590;
  assign n592 = \V88(7)  & ~n201;
  assign n593 = ~n195 & n592;
  assign n594 = ~n190 & n593;
  assign n595 = \V88(11)  & ~n190;
  assign n596 = ~n195 & n595;
  assign n597 = n201 & n596;
  assign n598 = \V88(14)  & ~n190;
  assign n599 = n195 & n598;
  assign n600 = ~n201 & n599;
  assign n601 = \V88(22)  & ~n190;
  assign n602 = n195 & n601;
  assign n603 = n201 & n602;
  assign n604 = n238 & ~n603;
  assign n605 = ~n600 & n604;
  assign n606 = ~n597 & n605;
  assign \V151(22)  = n594 | ~n606;
  assign n608 = \V88(10)  & ~n201;
  assign n609 = ~n195 & n608;
  assign n610 = ~n190 & n609;
  assign n611 = ~n195 & n598;
  assign n612 = n201 & n611;
  assign n613 = n195 & n480;
  assign n614 = ~n201 & n613;
  assign n615 = \V88(25)  & ~n190;
  assign n616 = n195 & n615;
  assign n617 = n201 & n616;
  assign n618 = n238 & ~n617;
  assign n619 = ~n614 & n618;
  assign n620 = ~n612 & n619;
  assign \V151(25)  = n610 | ~n620;
  assign n622 = \V88(9)  & ~n201;
  assign n623 = ~n195 & n622;
  assign n624 = ~n190 & n623;
  assign n625 = ~n195 & n535;
  assign n626 = n201 & n625;
  assign n627 = n195 & n422;
  assign n628 = ~n201 & n627;
  assign n629 = \V88(24)  & ~n190;
  assign n630 = n195 & n629;
  assign n631 = n201 & n630;
  assign n632 = n238 & ~n631;
  assign n633 = ~n628 & n632;
  assign n634 = ~n626 & n633;
  assign \V151(24)  = n624 | ~n634;
  assign n636 = \V88(2)  & ~n201;
  assign n637 = ~n195 & n636;
  assign n638 = ~n190 & n637;
  assign n639 = ~n201 & n355;
  assign n640 = n201 & n613;
  assign n641 = n238 & ~n640;
  assign n642 = ~n639 & n641;
  assign n643 = ~n401 & n642;
  assign \V151(17)  = n638 | ~n643;
  assign n645 = \V88(1)  & ~n201;
  assign n646 = ~n195 & n645;
  assign n647 = ~n190 & n646;
  assign n648 = ~n201 & n368;
  assign n649 = n201 & n627;
  assign n650 = n238 & ~n649;
  assign n651 = ~n648 & n650;
  assign n652 = ~n412 & n651;
  assign \V151(16)  = n647 | ~n652;
  assign n654 = \V88(4)  & ~n201;
  assign n655 = ~n195 & n654;
  assign n656 = ~n190 & n655;
  assign n657 = n195 & n595;
  assign n658 = ~n201 & n657;
  assign n659 = n201 & n426;
  assign n660 = n238 & ~n659;
  assign n661 = ~n658 & n660;
  assign n662 = ~n508 & n661;
  assign \V151(19)  = n656 | ~n662;
  assign n664 = \V88(3)  & ~n201;
  assign n665 = ~n195 & n664;
  assign n666 = ~n190 & n665;
  assign n667 = n195 & n532;
  assign n668 = ~n201 & n667;
  assign n669 = n201 & n442;
  assign n670 = n238 & ~n669;
  assign n671 = ~n668 & n670;
  assign n672 = ~n521 & n671;
  assign \V151(18)  = n666 | ~n672;
  assign n674 = \V56(28)  & ~n201;
  assign n675 = ~n195 & n674;
  assign n676 = ~n190 & n675;
  assign n677 = ~n195 & n313;
  assign n678 = n201 & n677;
  assign n679 = ~n201 & n228;
  assign n680 = n201 & n657;
  assign n681 = n238 & ~n680;
  assign n682 = ~n679 & n681;
  assign n683 = ~n678 & n682;
  assign \V151(11)  = n676 | ~n683;
  assign n685 = \V56(27)  & ~n201;
  assign n686 = ~n195 & n685;
  assign n687 = ~n190 & n686;
  assign n688 = ~n195 & n211;
  assign n689 = n201 & n688;
  assign n690 = ~n201 & n253;
  assign n691 = n201 & n667;
  assign n692 = n238 & ~n691;
  assign n693 = ~n690 & n692;
  assign n694 = ~n689 & n693;
  assign \V151(10)  = n687 | ~n694;
  assign n696 = \V56(30)  & ~n201;
  assign n697 = ~n195 & n696;
  assign n698 = ~n190 & n697;
  assign n699 = ~n201 & n268;
  assign n700 = n201 & n536;
  assign n701 = n238 & ~n700;
  assign n702 = ~n699 & n701;
  assign n703 = ~n470 & n702;
  assign \V151(13)  = n698 | ~n703;
  assign n705 = \V56(29)  & ~n201;
  assign n706 = ~n195 & n705;
  assign n707 = ~n190 & n706;
  assign n708 = ~n201 & n284;
  assign n709 = n201 & n560;
  assign n710 = n238 & ~n709;
  assign n711 = ~n708 & n710;
  assign n712 = ~n497 & n711;
  assign \V151(12)  = n707 | ~n712;
  assign n714 = \V56(13)  & ~n201;
  assign n715 = ~n195 & n714;
  assign n716 = ~n190 & n715;
  assign n717 = \V56(17)  & ~n190;
  assign n718 = ~n195 & n717;
  assign n719 = n201 & n718;
  assign n720 = \V56(20)  & n209;
  assign n721 = n201 & n281;
  assign n722 = ~n190 & ~n721;
  assign n723 = ~n720 & n722;
  assign n724 = ~n719 & n723;
  assign \V119(27)  = n716 | ~n724;
  assign n726 = \V88(0)  & ~n201;
  assign n727 = ~n195 & n726;
  assign n728 = ~n190 & n727;
  assign n729 = ~n201 & n327;
  assign n730 = n201 & n583;
  assign n731 = n238 & ~n730;
  assign n732 = ~n729 & n731;
  assign n733 = ~n378 & n732;
  assign \V151(15)  = n728 | ~n733;
  assign n735 = \V56(12)  & ~n201;
  assign n736 = ~n195 & n735;
  assign n737 = ~n190 & n736;
  assign n738 = \V56(16)  & ~n190;
  assign n739 = ~n195 & n738;
  assign n740 = n201 & n739;
  assign n741 = \V56(19)  & n209;
  assign n742 = n201 & n225;
  assign n743 = ~n190 & ~n742;
  assign n744 = ~n741 & n743;
  assign n745 = ~n740 & n744;
  assign \V119(26)  = n737 | ~n745;
  assign n747 = \V56(31)  & ~n201;
  assign n748 = ~n195 & n747;
  assign n749 = ~n190 & n748;
  assign n750 = ~n201 & n342;
  assign n751 = n201 & n599;
  assign n752 = n238 & ~n751;
  assign n753 = ~n750 & n752;
  assign n754 = ~n390 & n753;
  assign \V151(14)  = n749 | ~n754;
  assign n756 = \V56(15)  & ~n201;
  assign n757 = ~n195 & n756;
  assign n758 = ~n190 & n757;
  assign n759 = \V56(19)  & ~n190;
  assign n760 = ~n195 & n759;
  assign n761 = n201 & n760;
  assign n762 = \V56(22)  & n209;
  assign n763 = n201 & n339;
  assign n764 = ~n190 & ~n763;
  assign n765 = ~n762 & n764;
  assign n766 = ~n761 & n765;
  assign \V119(29)  = n758 | ~n766;
  assign n768 = \V56(14)  & ~n201;
  assign n769 = ~n195 & n768;
  assign n770 = ~n190 & n769;
  assign n771 = \V56(18)  & ~n190;
  assign n772 = ~n195 & n771;
  assign n773 = n201 & n772;
  assign n774 = \V56(21)  & n209;
  assign n775 = n201 & n265;
  assign n776 = ~n190 & ~n775;
  assign n777 = ~n774 & n776;
  assign n778 = ~n773 & n777;
  assign \V119(28)  = n770 | ~n778;
  assign n780 = \V56(7)  & ~n201;
  assign n781 = ~n195 & n780;
  assign n782 = ~n190 & n781;
  assign n783 = \V56(11)  & ~n190;
  assign n784 = ~n195 & n783;
  assign n785 = n201 & n784;
  assign n786 = \V56(14)  & n209;
  assign n787 = n195 & n293;
  assign n788 = n201 & n787;
  assign n789 = ~n190 & ~n788;
  assign n790 = ~n786 & n789;
  assign n791 = ~n785 & n790;
  assign \V119(21)  = n782 | ~n791;
  assign n793 = \V56(6)  & ~n201;
  assign n794 = ~n195 & n793;
  assign n795 = ~n190 & n794;
  assign n796 = ~n195 & n547;
  assign n797 = n201 & n796;
  assign n798 = \V56(13)  & n209;
  assign n799 = n195 & n308;
  assign n800 = n201 & n799;
  assign n801 = ~n190 & ~n800;
  assign n802 = ~n798 & n801;
  assign n803 = ~n797 & n802;
  assign \V119(20)  = n795 | ~n803;
  assign n805 = \V56(9)  & ~n201;
  assign n806 = ~n195 & n805;
  assign n807 = ~n190 & n806;
  assign n808 = \V56(13)  & ~n190;
  assign n809 = ~n195 & n808;
  assign n810 = n201 & n809;
  assign n811 = \V56(16)  & n209;
  assign n812 = n201 & n311;
  assign n813 = ~n190 & ~n812;
  assign n814 = ~n811 & n813;
  assign n815 = ~n810 & n814;
  assign \V119(23)  = n807 | ~n815;
  assign n817 = \V56(8)  & ~n201;
  assign n818 = ~n195 & n817;
  assign n819 = ~n190 & n818;
  assign n820 = \V56(12)  & ~n190;
  assign n821 = ~n195 & n820;
  assign n822 = n201 & n821;
  assign n823 = \V56(15)  & n209;
  assign n824 = n195 & n246;
  assign n825 = n201 & n824;
  assign n826 = ~n190 & ~n825;
  assign n827 = ~n823 & n826;
  assign n828 = ~n822 & n827;
  assign \V119(22)  = n819 | ~n828;
  assign n830 = \V56(11)  & ~n201;
  assign n831 = ~n195 & n830;
  assign n832 = ~n190 & n831;
  assign n833 = \V56(15)  & ~n190;
  assign n834 = ~n195 & n833;
  assign n835 = n201 & n834;
  assign n836 = \V56(18)  & n209;
  assign n837 = n201 & n250;
  assign n838 = ~n190 & ~n837;
  assign n839 = ~n836 & n838;
  assign n840 = ~n835 & n839;
  assign \V119(25)  = n832 | ~n840;
  assign n842 = \V56(10)  & ~n201;
  assign n843 = ~n195 & n842;
  assign n844 = ~n190 & n843;
  assign n845 = \V56(14)  & ~n190;
  assign n846 = ~n195 & n845;
  assign n847 = n201 & n846;
  assign n848 = \V56(17)  & n209;
  assign n849 = n201 & n296;
  assign n850 = ~n190 & ~n849;
  assign n851 = ~n848 & n850;
  assign n852 = ~n847 & n851;
  assign \V119(24)  = n844 | ~n852;
  assign n854 = \V56(3)  & ~n201;
  assign n855 = ~n195 & n854;
  assign n856 = ~n190 & n855;
  assign n857 = ~n195 & n522;
  assign n858 = n201 & n857;
  assign n859 = \V56(10)  & n209;
  assign n860 = n195 & n771;
  assign n861 = n201 & n860;
  assign n862 = ~n190 & ~n861;
  assign n863 = ~n859 & n862;
  assign n864 = ~n858 & n863;
  assign \V119(17)  = n856 | ~n864;
  assign n866 = \V56(2)  & ~n201;
  assign n867 = ~n195 & n866;
  assign n868 = ~n190 & n867;
  assign n869 = ~n195 & n402;
  assign n870 = n201 & n869;
  assign n871 = \V56(9)  & n209;
  assign n872 = n195 & n717;
  assign n873 = n201 & n872;
  assign n874 = ~n190 & ~n873;
  assign n875 = ~n871 & n874;
  assign n876 = ~n870 & n875;
  assign \V119(16)  = n868 | ~n876;
  assign n878 = \V56(5)  & ~n201;
  assign n879 = ~n195 & n878;
  assign n880 = ~n190 & n879;
  assign n881 = ~n195 & n571;
  assign n882 = n201 & n881;
  assign n883 = \V56(12)  & n209;
  assign n884 = n195 & n205;
  assign n885 = n201 & n884;
  assign n886 = ~n190 & ~n885;
  assign n887 = ~n883 & n886;
  assign n888 = ~n882 & n887;
  assign \V119(19)  = n880 | ~n888;
  assign n890 = \V56(4)  & ~n201;
  assign n891 = ~n195 & n890;
  assign n892 = ~n190 & n891;
  assign n893 = ~n195 & n510;
  assign n894 = n201 & n893;
  assign n895 = \V56(11)  & n209;
  assign n896 = n195 & n759;
  assign n897 = n201 & n896;
  assign n898 = ~n190 & ~n897;
  assign n899 = ~n895 & n898;
  assign n900 = ~n894 & n899;
  assign \V119(18)  = n892 | ~n900;
  assign n902 = \V24(11)  & ~n201;
  assign n903 = ~n195 & n902;
  assign n904 = ~n190 & n903;
  assign n905 = ~n195 & n498;
  assign n906 = n201 & n905;
  assign n907 = \V56(4)  & n209;
  assign n908 = n195 & n820;
  assign n909 = n201 & n908;
  assign n910 = ~n190 & ~n909;
  assign n911 = ~n907 & n910;
  assign n912 = ~n906 & n911;
  assign \V119(11)  = n904 | ~n912;
  assign n914 = \V24(10)  & ~n201;
  assign n915 = ~n195 & n914;
  assign n916 = ~n190 & n915;
  assign n917 = \V56(3)  & n209;
  assign n918 = n195 & n783;
  assign n919 = n201 & n918;
  assign n920 = ~n190 & ~n919;
  assign n921 = ~n917 & n920;
  assign n922 = ~n597 & n921;
  assign \V119(10)  = n916 | ~n922;
  assign n924 = \V24(13)  & ~n201;
  assign n925 = ~n195 & n924;
  assign n926 = ~n190 & n925;
  assign n927 = ~n195 & n391;
  assign n928 = n201 & n927;
  assign n929 = \V56(6)  & n209;
  assign n930 = n195 & n845;
  assign n931 = n201 & n930;
  assign n932 = ~n190 & ~n931;
  assign n933 = ~n929 & n932;
  assign n934 = ~n928 & n933;
  assign \V119(13)  = n926 | ~n934;
  assign n936 = \V88(16)  & ~n201;
  assign n937 = ~n195 & n936;
  assign n938 = ~n190 & n937;
  assign n939 = ~n195 & n483;
  assign n940 = n201 & n939;
  assign n941 = ~n201 & n586;
  assign n942 = \V88(31)  & ~n190;
  assign n943 = n195 & n942;
  assign n944 = n201 & n943;
  assign n945 = n238 & ~n944;
  assign n946 = ~n941 & n945;
  assign n947 = ~n940 & n946;
  assign \V151(31)  = n938 | ~n947;
  assign n949 = \V24(12)  & ~n201;
  assign n950 = ~n195 & n949;
  assign n951 = ~n190 & n950;
  assign n952 = ~n195 & n471;
  assign n953 = n201 & n952;
  assign n954 = \V56(5)  & n209;
  assign n955 = n195 & n808;
  assign n956 = n201 & n955;
  assign n957 = ~n190 & ~n956;
  assign n958 = ~n954 & n957;
  assign n959 = ~n953 & n958;
  assign \V119(12)  = n951 | ~n959;
  assign n961 = \V88(15)  & ~n201;
  assign n962 = ~n195 & n961;
  assign n963 = ~n190 & n962;
  assign n964 = ~n195 & n425;
  assign n965 = n201 & n964;
  assign n966 = ~n201 & n602;
  assign n967 = \V88(30)  & ~n190;
  assign n968 = n195 & n967;
  assign n969 = n201 & n968;
  assign n970 = n238 & ~n969;
  assign n971 = ~n966 & n970;
  assign n972 = ~n965 & n971;
  assign \V151(30)  = n963 | ~n972;
  assign n974 = \V56(1)  & ~n201;
  assign n975 = ~n195 & n974;
  assign n976 = ~n190 & n975;
  assign n977 = ~n195 & n413;
  assign n978 = n201 & n977;
  assign n979 = \V56(8)  & n209;
  assign n980 = n195 & n738;
  assign n981 = n201 & n980;
  assign n982 = ~n190 & ~n981;
  assign n983 = ~n979 & n982;
  assign n984 = ~n978 & n983;
  assign \V119(15)  = n976 | ~n984;
  assign n986 = \V24(14)  & ~n201;
  assign n987 = ~n195 & n986;
  assign n988 = ~n190 & n987;
  assign n989 = ~n195 & n379;
  assign n990 = n201 & n989;
  assign n991 = \V56(7)  & n209;
  assign n992 = n195 & n833;
  assign n993 = n201 & n992;
  assign n994 = ~n190 & ~n993;
  assign n995 = ~n991 & n994;
  assign n996 = ~n990 & n995;
  assign \V119(14)  = n988 | ~n996;
endmodule


