// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:06 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_,
    i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_,
    i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_, i_40_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_,
    i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_,
    i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_,
    i_40_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_;
  wire n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
    n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1053, n1055, n1056, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1083, n1084,
    n1085, n1086, n1087, n1089, n1090, n1091, n1093, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1463, n1464, n1465, n1466,
    n1468, n1470, n1472, n1473, n1475, n1477, n1478, n1479, n1480, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1495, n1496, n1497, n1498, n1499, n1500, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638;
  assign n77 = ~i_32_ & i_33_;
  assign n78 = ~i_34_ & i_35_;
  assign n79 = n77 & n78;
  assign n80 = ~i_7_ & n79;
  assign n81 = i_36_ & n80;
  assign n82 = ~i_25_ & ~i_26_;
  assign n83 = ~i_37_ & ~i_39_;
  assign n84 = ~i_38_ & n83;
  assign n85 = n82 & n84;
  assign n86 = n81 & n85;
  assign n87 = i_12_ & i_15_;
  assign n88 = i_11_ & i_15_;
  assign n89 = ~n87 & ~n88;
  assign n90 = ~i_5_ & ~n89;
  assign n91 = ~i_7_ & n90;
  assign n92 = i_24_ & n77;
  assign n93 = ~i_36_ & n78;
  assign n94 = n92 & n93;
  assign n95 = n91 & n94;
  assign n96 = ~i_38_ & i_40_;
  assign n97 = i_37_ & n96;
  assign n98 = ~i_39_ & n97;
  assign n99 = i_9_ & n98;
  assign n100 = n95 & n99;
  assign n101 = i_24_ & ~i_32_;
  assign n102 = ~i_36_ & n98;
  assign n103 = i_33_ & ~i_34_;
  assign n104 = i_35_ & n103;
  assign n105 = n102 & n104;
  assign n106 = n101 & n105;
  assign n107 = ~i_9_ & n91;
  assign n108 = i_18_ & n107;
  assign n109 = n106 & n108;
  assign n110 = ~n100 & ~n109;
  assign n111 = ~i_21_ & ~i_23_;
  assign n112 = ~i_18_ & ~i_19_;
  assign n113 = i_22_ & ~n112;
  assign n114 = n111 & n113;
  assign n115 = ~n110 & n114;
  assign n116 = i_38_ & i_39_;
  assign n117 = ~i_37_ & n116;
  assign n118 = ~i_36_ & n117;
  assign n119 = n79 & n91;
  assign n120 = i_21_ & n119;
  assign n121 = ~i_5_ & ~i_7_;
  assign n122 = ~i_31_ & n77;
  assign n123 = ~i_34_ & n122;
  assign n124 = n121 & n123;
  assign n125 = ~i_35_ & n124;
  assign n126 = ~i_16_ & ~i_17_;
  assign n127 = ~i_12_ & n88;
  assign n128 = n126 & n127;
  assign n129 = n125 & n128;
  assign n130 = ~n120 & ~n129;
  assign n131 = n118 & ~n130;
  assign n132 = ~i_34_ & ~i_35_;
  assign n133 = ~i_36_ & ~i_37_;
  assign n134 = i_40_ & n116;
  assign n135 = n133 & n134;
  assign n136 = n132 & n135;
  assign n137 = i_12_ & n121;
  assign n138 = i_15_ & n126;
  assign n139 = n122 & n138;
  assign n140 = n137 & n139;
  assign n141 = n136 & n140;
  assign n142 = ~n131 & ~n141;
  assign n143 = ~n115 & n142;
  assign n144 = ~n86 & n143;
  assign n145 = i_36_ & i_40_;
  assign n146 = n117 & n132;
  assign n147 = n145 & n146;
  assign n148 = n77 & n147;
  assign n149 = ~i_35_ & n77;
  assign n150 = i_38_ & ~i_39_;
  assign n151 = i_37_ & n150;
  assign n152 = n145 & n151;
  assign n153 = ~i_34_ & n152;
  assign n154 = n149 & n153;
  assign n155 = ~n148 & ~n154;
  assign n156 = ~i_2_ & ~i_3_;
  assign n157 = ~i_1_ & ~i_4_;
  assign n158 = n156 & n157;
  assign n159 = i_0_ & ~n158;
  assign n160 = ~n155 & n159;
  assign n161 = ~i_7_ & n160;
  assign n162 = ~i_9_ & ~i_18_;
  assign n163 = ~i_9_ & ~i_19_;
  assign n164 = ~n112 & ~n163;
  assign n165 = ~n162 & n164;
  assign n166 = n119 & ~n165;
  assign n167 = n102 & n166;
  assign n168 = i_34_ & n77;
  assign n169 = ~i_35_ & ~i_36_;
  assign n170 = n168 & n169;
  assign n171 = ~i_7_ & n170;
  assign n172 = i_39_ & i_40_;
  assign n173 = ~i_37_ & n172;
  assign n174 = n171 & n173;
  assign n175 = ~i_38_ & n174;
  assign n176 = i_34_ & n169;
  assign n177 = ~i_7_ & n77;
  assign n178 = i_38_ & i_40_;
  assign n179 = ~i_39_ & n178;
  assign n180 = n177 & n179;
  assign n181 = n176 & n180;
  assign n182 = ~n175 & ~n181;
  assign n183 = ~n167 & n182;
  assign n184 = ~n161 & n183;
  assign n185 = i_36_ & ~i_37_;
  assign n186 = ~i_34_ & n185;
  assign n187 = n149 & n186;
  assign n188 = n96 & n187;
  assign n189 = i_39_ & n188;
  assign n190 = i_11_ & n189;
  assign n191 = ~i_7_ & n190;
  assign n192 = ~i_34_ & n77;
  assign n193 = ~i_35_ & i_36_;
  assign n194 = n192 & n193;
  assign n195 = ~i_7_ & n194;
  assign n196 = ~i_40_ & n195;
  assign n197 = ~i_37_ & n150;
  assign n198 = i_10_ & i_27_;
  assign n199 = n197 & n198;
  assign n200 = n196 & n199;
  assign n201 = i_36_ & i_37_;
  assign n202 = i_35_ & n201;
  assign n203 = n192 & n202;
  assign n204 = ~i_3_ & i_4_;
  assign n205 = i_1_ & ~i_2_;
  assign n206 = n204 & n205;
  assign n207 = n203 & ~n206;
  assign n208 = ~i_38_ & ~i_40_;
  assign n209 = i_0_ & ~i_7_;
  assign n210 = n208 & n209;
  assign n211 = n207 & n210;
  assign n212 = i_15_ & ~i_24_;
  assign n213 = n79 & n212;
  assign n214 = i_11_ & n121;
  assign n215 = n213 & n214;
  assign n216 = ~i_38_ & ~i_39_;
  assign n217 = ~i_36_ & n216;
  assign n218 = i_40_ & n217;
  assign n219 = ~n116 & ~n216;
  assign n220 = n133 & ~n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = n215 & ~n221;
  assign n223 = ~n211 & ~n222;
  assign n224 = ~n200 & n223;
  assign n225 = ~n191 & n224;
  assign n226 = n184 & n225;
  assign n227 = n144 & n226;
  assign n228 = n122 & n132;
  assign n229 = ~i_9_ & ~i_16_;
  assign n230 = n91 & n229;
  assign n231 = n228 & n230;
  assign n232 = i_37_ & n217;
  assign n233 = n231 & n232;
  assign n234 = ~i_36_ & i_39_;
  assign n235 = ~i_37_ & n234;
  assign n236 = ~i_36_ & n96;
  assign n237 = ~n235 & ~n236;
  assign n238 = n229 & ~n237;
  assign n239 = n125 & n238;
  assign n240 = n77 & n169;
  assign n241 = ~i_31_ & n240;
  assign n242 = ~i_34_ & n241;
  assign n243 = ~i_5_ & ~i_9_;
  assign n244 = ~i_7_ & n243;
  assign n245 = n116 & n244;
  assign n246 = n242 & n245;
  assign n247 = ~i_17_ & n246;
  assign n248 = ~n239 & ~n247;
  assign n249 = n88 & ~n248;
  assign n250 = ~i_34_ & n169;
  assign n251 = i_37_ & n216;
  assign n252 = n250 & n251;
  assign n253 = ~i_17_ & n252;
  assign n254 = n122 & n253;
  assign n255 = n107 & n254;
  assign n256 = ~n249 & ~n255;
  assign n257 = ~n233 & n256;
  assign n258 = n87 & n239;
  assign n259 = ~i_37_ & i_40_;
  assign n260 = ~i_17_ & n87;
  assign n261 = n259 & ~n260;
  assign n262 = n246 & ~n261;
  assign n263 = n137 & n213;
  assign n264 = n118 & n263;
  assign n265 = ~n262 & ~n264;
  assign n266 = ~n258 & n265;
  assign n267 = ~n118 & ~n232;
  assign n268 = i_34_ & n149;
  assign n269 = ~i_7_ & n268;
  assign n270 = ~n158 & n269;
  assign n271 = ~n267 & n270;
  assign n272 = i_11_ & i_12_;
  assign n273 = i_15_ & n272;
  assign n274 = i_38_ & ~i_40_;
  assign n275 = n133 & n274;
  assign n276 = i_39_ & n275;
  assign n277 = ~n273 & n276;
  assign n278 = n125 & n277;
  assign n279 = n77 & n93;
  assign n280 = n117 & n279;
  assign n281 = ~i_22_ & n280;
  assign n282 = n91 & n281;
  assign n283 = i_13_ & n121;
  assign n284 = n89 & n283;
  assign n285 = n228 & n284;
  assign n286 = ~n232 & n237;
  assign n287 = n285 & ~n286;
  assign n288 = ~n137 & ~n214;
  assign n289 = n139 & ~n288;
  assign n290 = n252 & n289;
  assign n291 = ~n287 & ~n290;
  assign n292 = ~n282 & n291;
  assign n293 = ~n278 & n292;
  assign n294 = ~n271 & n293;
  assign n295 = n266 & n294;
  assign n296 = n257 & n295;
  assign n297 = i_37_ & ~i_40_;
  assign n298 = n217 & n263;
  assign n299 = ~n297 & n298;
  assign n300 = ~i_37_ & ~i_38_;
  assign n301 = i_0_ & ~i_1_;
  assign n302 = ~i_4_ & n301;
  assign n303 = n171 & n302;
  assign n304 = n300 & n303;
  assign n305 = ~i_11_ & ~i_12_;
  assign n306 = ~i_7_ & n305;
  assign n307 = ~i_5_ & n306;
  assign n308 = n79 & n307;
  assign n309 = i_13_ & n218;
  assign n310 = n308 & n309;
  assign n311 = ~n304 & ~n310;
  assign n312 = ~n299 & n311;
  assign n313 = ~i_15_ & n283;
  assign n314 = n79 & n313;
  assign n315 = i_21_ & i_22_;
  assign n316 = n91 & n315;
  assign n317 = n92 & n316;
  assign n318 = i_37_ & n78;
  assign n319 = n317 & n318;
  assign n320 = ~n314 & ~n319;
  assign n321 = n218 & ~n320;
  assign n322 = n231 & n275;
  assign n323 = ~i_18_ & n118;
  assign n324 = n79 & n323;
  assign n325 = n107 & n324;
  assign n326 = ~n322 & ~n325;
  assign n327 = ~n321 & n326;
  assign n328 = n312 & n327;
  assign n329 = n91 & n101;
  assign n330 = ~i_22_ & n329;
  assign n331 = n105 & n330;
  assign n332 = i_38_ & n78;
  assign n333 = n201 & n332;
  assign n334 = i_33_ & n333;
  assign n335 = i_33_ & n169;
  assign n336 = i_34_ & n335;
  assign n337 = n300 & n336;
  assign n338 = ~n334 & ~n337;
  assign n339 = ~i_7_ & ~i_32_;
  assign n340 = i_2_ & n301;
  assign n341 = ~i_3_ & n340;
  assign n342 = n339 & n341;
  assign n343 = ~n338 & n342;
  assign n344 = ~n331 & ~n343;
  assign n345 = i_39_ & n297;
  assign n346 = ~i_7_ & n279;
  assign n347 = i_0_ & n346;
  assign n348 = n345 & n347;
  assign n349 = i_38_ & n348;
  assign n350 = i_37_ & i_38_;
  assign n351 = n81 & n302;
  assign n352 = n350 & n351;
  assign n353 = ~n349 & ~n352;
  assign n354 = n275 & n285;
  assign n355 = i_37_ & i_39_;
  assign n356 = n208 & n355;
  assign n357 = n81 & n356;
  assign n358 = ~n354 & ~n357;
  assign n359 = i_39_ & n236;
  assign n360 = n268 & n359;
  assign n361 = n283 & n360;
  assign n362 = n358 & ~n361;
  assign n363 = n353 & n362;
  assign n364 = i_13_ & n308;
  assign n365 = ~n314 & ~n364;
  assign n366 = n220 & ~n365;
  assign n367 = ~i_7_ & i_38_;
  assign n368 = n194 & n367;
  assign n369 = n345 & n368;
  assign n370 = ~n366 & ~n369;
  assign n371 = n77 & n91;
  assign n372 = ~i_38_ & n169;
  assign n373 = n172 & n372;
  assign n374 = i_34_ & n373;
  assign n375 = n78 & n220;
  assign n376 = ~i_40_ & n375;
  assign n377 = ~n374 & ~n376;
  assign n378 = n371 & ~n377;
  assign n379 = n370 & ~n378;
  assign n380 = n363 & n379;
  assign n381 = n344 & n380;
  assign n382 = i_29_ & i_30_;
  assign n383 = ~i_28_ & ~n382;
  assign n384 = ~i_28_ & n382;
  assign n385 = ~i_29_ & ~i_30_;
  assign n386 = ~n384 & ~n385;
  assign n387 = n121 & ~n386;
  assign n388 = n242 & n356;
  assign n389 = ~i_39_ & i_40_;
  assign n390 = i_38_ & n169;
  assign n391 = n122 & n390;
  assign n392 = n389 & n391;
  assign n393 = ~n388 & ~n392;
  assign n394 = n387 & ~n393;
  assign n395 = ~n383 & n394;
  assign n396 = n381 & ~n395;
  assign n397 = n328 & n396;
  assign n398 = n296 & n397;
  assign o_0_ = ~n227 | ~n398;
  assign n400 = i_16_ & i_17_;
  assign n401 = i_9_ & ~n126;
  assign n402 = ~n400 & ~n401;
  assign n403 = n169 & n192;
  assign n404 = i_31_ & n403;
  assign n405 = n402 & n404;
  assign n406 = ~i_5_ & n405;
  assign n407 = ~i_5_ & n305;
  assign n408 = n77 & n407;
  assign n409 = ~i_13_ & n408;
  assign n410 = n236 & n318;
  assign n411 = ~i_37_ & n169;
  assign n412 = ~i_40_ & n150;
  assign n413 = n411 & n412;
  assign n414 = n96 & n355;
  assign n415 = n169 & n414;
  assign n416 = ~n413 & ~n415;
  assign n417 = ~n410 & n416;
  assign n418 = ~n83 & ~n355;
  assign n419 = ~i_38_ & n418;
  assign n420 = ~n259 & ~n419;
  assign n421 = ~n150 & n250;
  assign n422 = ~n420 & n421;
  assign n423 = n417 & ~n422;
  assign n424 = ~n375 & n423;
  assign n425 = n409 & ~n424;
  assign n426 = i_24_ & n90;
  assign n427 = ~i_37_ & n389;
  assign n428 = n426 & n427;
  assign n429 = n279 & n428;
  assign n430 = ~i_37_ & ~i_40_;
  assign n431 = n150 & n430;
  assign n432 = n170 & n431;
  assign n433 = ~n429 & ~n432;
  assign n434 = n116 & n259;
  assign n435 = n158 & n170;
  assign n436 = n434 & n435;
  assign n437 = i_36_ & n79;
  assign n438 = n300 & n437;
  assign n439 = ~n82 & n438;
  assign n440 = ~n436 & ~n439;
  assign n441 = n433 & n440;
  assign n442 = ~n425 & n441;
  assign n443 = ~n406 & n442;
  assign n444 = ~i_5_ & ~i_15_;
  assign n445 = ~i_13_ & n444;
  assign n446 = ~n173 & ~n251;
  assign n447 = n169 & ~n446;
  assign n448 = ~i_38_ & i_39_;
  assign n449 = ~n96 & ~n448;
  assign n450 = n411 & ~n449;
  assign n451 = ~n447 & ~n450;
  assign n452 = n192 & ~n451;
  assign n453 = n77 & ~n417;
  assign n454 = n79 & n133;
  assign n455 = n216 & n454;
  assign n456 = ~n280 & ~n455;
  assign n457 = ~n453 & n456;
  assign n458 = ~n452 & n457;
  assign n459 = n445 & ~n458;
  assign n460 = i_40_ & n448;
  assign n461 = i_12_ & n460;
  assign n462 = ~i_11_ & n461;
  assign n463 = i_36_ & n462;
  assign n464 = ~i_37_ & n463;
  assign n465 = ~i_36_ & i_37_;
  assign n466 = i_35_ & n465;
  assign n467 = ~n172 & ~n412;
  assign n468 = n466 & ~n467;
  assign n469 = i_37_ & n193;
  assign n470 = n134 & n469;
  assign n471 = ~n468 & ~n470;
  assign n472 = ~i_5_ & i_31_;
  assign n473 = n169 & n472;
  assign n474 = ~n87 & n473;
  assign n475 = i_37_ & ~i_38_;
  assign n476 = n234 & n475;
  assign n477 = i_35_ & n476;
  assign n478 = ~n474 & ~n477;
  assign n479 = i_35_ & ~i_37_;
  assign n480 = n179 & n479;
  assign n481 = i_35_ & n185;
  assign n482 = i_39_ & ~i_40_;
  assign n483 = ~n448 & ~n482;
  assign n484 = n481 & ~n483;
  assign n485 = ~n480 & ~n484;
  assign n486 = n478 & n485;
  assign n487 = n471 & n486;
  assign n488 = n90 & ~n272;
  assign n489 = ~i_14_ & n87;
  assign n490 = ~i_5_ & n489;
  assign n491 = ~n488 & ~n490;
  assign n492 = n169 & n251;
  assign n493 = ~n402 & n492;
  assign n494 = ~n491 & n493;
  assign n495 = n487 & ~n494;
  assign n496 = ~n464 & n495;
  assign n497 = n192 & ~n496;
  assign o_15_ = i_7_ & i_33_;
  assign n499 = n77 & ~n402;
  assign n500 = n90 & n499;
  assign n501 = n136 & n500;
  assign n502 = i_36_ & n300;
  assign n503 = ~i_39_ & ~i_40_;
  assign n504 = n502 & n503;
  assign n505 = n268 & n504;
  assign n506 = ~n501 & ~n505;
  assign n507 = ~i_32_ & n472;
  assign n508 = ~n251 & n507;
  assign n509 = ~i_36_ & n103;
  assign n510 = ~i_35_ & n509;
  assign n511 = n508 & n510;
  assign n512 = ~i_34_ & n149;
  assign n513 = i_14_ & n272;
  assign n514 = i_15_ & n513;
  assign n515 = ~n402 & n514;
  assign n516 = n135 & n515;
  assign n517 = n512 & n516;
  assign n518 = ~n511 & ~n517;
  assign n519 = n506 & n518;
  assign n520 = ~o_15_ & n519;
  assign n521 = ~n497 & n520;
  assign n522 = ~n459 & n521;
  assign o_1_ = ~n443 | ~n522;
  assign n524 = ~i_21_ & n232;
  assign n525 = i_23_ & i_24_;
  assign n526 = n165 & n525;
  assign n527 = i_22_ & n526;
  assign n528 = n90 & n527;
  assign n529 = n524 & n528;
  assign n530 = n79 & n529;
  assign n531 = n84 & n437;
  assign n532 = ~n82 & n531;
  assign n533 = n241 & n356;
  assign n534 = ~i_36_ & n179;
  assign n535 = n228 & n534;
  assign n536 = ~n533 & ~n535;
  assign n537 = ~n383 & ~n386;
  assign n538 = ~i_5_ & ~n537;
  assign n539 = ~n536 & n538;
  assign n540 = ~n532 & ~n539;
  assign n541 = ~n530 & n540;
  assign n542 = i_35_ & n133;
  assign n543 = n445 & n542;
  assign n544 = n389 & n543;
  assign n545 = ~n449 & n469;
  assign n546 = ~n480 & ~n545;
  assign n547 = ~i_40_ & n116;
  assign n548 = n481 & n547;
  assign n549 = ~i_40_ & n216;
  assign n550 = ~n134 & ~n549;
  assign n551 = n466 & ~n550;
  assign n552 = ~n548 & ~n551;
  assign n553 = n546 & n552;
  assign n554 = ~n544 & n553;
  assign n555 = n192 & ~n554;
  assign n556 = i_22_ & ~n162;
  assign n557 = n426 & n556;
  assign n558 = n134 & n557;
  assign n559 = ~i_21_ & n558;
  assign n560 = n279 & n559;
  assign n561 = ~n555 & ~n560;
  assign n562 = n541 & n561;
  assign n563 = ~n136 & ~n252;
  assign n564 = n122 & ~n563;
  assign n565 = n488 & n564;
  assign n566 = ~n402 & n565;
  assign n567 = ~o_15_ & ~n566;
  assign n568 = n179 & n186;
  assign n569 = n77 & n568;
  assign n570 = n150 & n187;
  assign n571 = ~n198 & n570;
  assign n572 = ~n569 & ~n571;
  assign n573 = n93 & n409;
  assign n574 = n427 & n573;
  assign n575 = ~n98 & ~n117;
  assign n576 = n435 & ~n575;
  assign n577 = n268 & n465;
  assign n578 = ~i_38_ & n482;
  assign n579 = n577 & n578;
  assign n580 = ~n576 & ~n579;
  assign n581 = ~n574 & n580;
  assign n582 = n433 & n581;
  assign n583 = n572 & n582;
  assign n584 = n567 & n583;
  assign o_2_ = ~n562 | ~n584;
  assign n586 = ~i_5_ & n126;
  assign n587 = n169 & n434;
  assign n588 = ~n252 & ~n587;
  assign n589 = n586 & ~n588;
  assign n590 = n87 & n589;
  assign n591 = ~i_28_ & n385;
  assign n592 = ~i_5_ & ~n591;
  assign n593 = n534 & n592;
  assign n594 = n243 & n355;
  assign n595 = n243 & n260;
  assign n596 = n234 & n595;
  assign n597 = ~n594 & ~n596;
  assign n598 = i_38_ & ~n597;
  assign n599 = ~n463 & ~n598;
  assign n600 = ~n593 & n599;
  assign n601 = n132 & ~n600;
  assign n602 = n252 & n488;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n590 & n603;
  assign n605 = n77 & ~n604;
  assign n606 = ~n102 & ~n276;
  assign n607 = n445 & ~n606;
  assign n608 = ~i_13_ & n102;
  assign n609 = i_15_ & n276;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~i_5_ & ~i_12_;
  assign n612 = ~n610 & n611;
  assign n613 = ~n607 & ~n612;
  assign n614 = ~n516 & n613;
  assign n615 = n149 & ~n614;
  assign n616 = ~n605 & ~n615;
  assign n617 = n97 & n170;
  assign n618 = ~n315 & n617;
  assign n619 = n192 & n547;
  assign n620 = i_21_ & i_23_;
  assign n621 = n479 & ~n620;
  assign n622 = n619 & n621;
  assign n623 = n117 & n240;
  assign n624 = ~n272 & n623;
  assign n625 = ~n281 & ~n624;
  assign n626 = ~n622 & n625;
  assign n627 = ~n618 & n626;
  assign n628 = n90 & ~n627;
  assign n629 = n90 & n279;
  assign n630 = ~i_24_ & n629;
  assign n631 = n117 & n630;
  assign n632 = ~i_32_ & n204;
  assign n633 = n340 & n632;
  assign n634 = n216 & n336;
  assign n635 = ~n334 & ~n634;
  assign n636 = n633 & ~n635;
  assign n637 = ~n631 & ~n636;
  assign n638 = ~n158 & n170;
  assign n639 = n251 & n638;
  assign n640 = n198 & n412;
  assign n641 = n187 & n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = ~o_15_ & n642;
  assign n644 = n637 & n643;
  assign n645 = ~i_35_ & n103;
  assign n646 = ~i_37_ & ~n116;
  assign n647 = ~i_32_ & n145;
  assign n648 = ~n646 & n647;
  assign n649 = n159 & n648;
  assign n650 = i_15_ & ~i_32_;
  assign n651 = ~i_5_ & n229;
  assign n652 = n650 & n651;
  assign n653 = ~i_36_ & n475;
  assign n654 = i_12_ & n653;
  assign n655 = ~i_12_ & i_38_;
  assign n656 = n234 & ~n655;
  assign n657 = ~n236 & ~n656;
  assign n658 = ~n654 & n657;
  assign n659 = n652 & ~n658;
  assign n660 = ~n305 & n659;
  assign n661 = ~n649 & ~n660;
  assign n662 = n645 & ~n661;
  assign n663 = n644 & ~n662;
  assign n664 = ~n628 & n663;
  assign n665 = n243 & ~n305;
  assign n666 = n240 & n431;
  assign n667 = i_15_ & ~i_16_;
  assign n668 = n666 & n667;
  assign n669 = ~i_21_ & n104;
  assign n670 = n650 & n669;
  assign n671 = n323 & n670;
  assign n672 = ~n668 & ~n671;
  assign n673 = n665 & ~n672;
  assign n674 = i_0_ & n79;
  assign n675 = ~i_38_ & n297;
  assign n676 = n674 & n675;
  assign n677 = ~n206 & n676;
  assign n678 = ~i_25_ & n531;
  assign n679 = ~n677 & ~n678;
  assign n680 = n430 & n633;
  assign n681 = n336 & n680;
  assign n682 = ~i_38_ & ~n302;
  assign n683 = n168 & n411;
  assign n684 = ~n116 & ~n503;
  assign n685 = n683 & ~n684;
  assign n686 = ~n682 & n685;
  assign n687 = ~n681 & ~n686;
  assign n688 = n679 & n687;
  assign n689 = ~n673 & n688;
  assign n690 = n216 & n630;
  assign n691 = n465 & n674;
  assign n692 = n192 & n475;
  assign n693 = ~i_5_ & n692;
  assign n694 = ~n691 & ~n693;
  assign n695 = n482 & ~n694;
  assign n696 = ~n690 & ~n695;
  assign n697 = ~n475 & ~n549;
  assign n698 = ~n315 & n629;
  assign n699 = ~n697 & n698;
  assign n700 = ~i_38_ & n389;
  assign n701 = n577 & n700;
  assign n702 = ~n699 & ~n701;
  assign n703 = n696 & n702;
  assign n704 = n689 & n703;
  assign n705 = i_35_ & n208;
  assign n706 = ~n355 & ~n465;
  assign n707 = n705 & ~n706;
  assign n708 = i_35_ & n503;
  assign n709 = ~n134 & ~n708;
  assign n710 = n201 & n302;
  assign n711 = ~n709 & n710;
  assign n712 = ~n707 & ~n711;
  assign n713 = n492 & n595;
  assign n714 = n243 & n547;
  assign n715 = n169 & n714;
  assign n716 = ~n713 & ~n715;
  assign n717 = ~n179 & ~n547;
  assign n718 = n481 & ~n717;
  assign n719 = ~i_14_ & n473;
  assign n720 = ~i_39_ & ~n96;
  assign n721 = n469 & ~n720;
  assign n722 = ~n719 & ~n721;
  assign n723 = ~n718 & n722;
  assign n724 = n716 & n723;
  assign n725 = n478 & n724;
  assign n726 = n712 & n725;
  assign n727 = n192 & ~n726;
  assign n728 = n704 & ~n727;
  assign n729 = n664 & n728;
  assign n730 = ~n511 & n729;
  assign o_3_ = ~n616 | ~n730;
  assign n732 = ~i_34_ & ~n538;
  assign n733 = n169 & n356;
  assign n734 = ~n732 & n733;
  assign n735 = ~i_34_ & n481;
  assign n736 = n302 & n318;
  assign n737 = ~n735 & ~n736;
  assign n738 = n547 & ~n737;
  assign n739 = ~n460 & ~n503;
  assign n740 = ~i_36_ & n318;
  assign n741 = ~n739 & n740;
  assign n742 = ~n738 & ~n741;
  assign n743 = ~n734 & n742;
  assign n744 = ~n568 & n743;
  assign n745 = n177 & ~n744;
  assign n746 = n303 & n578;
  assign n747 = ~n745 & ~n746;
  assign n748 = n133 & n460;
  assign n749 = ~i_13_ & n512;
  assign n750 = n748 & n749;
  assign n751 = n217 & n259;
  assign n752 = n79 & n751;
  assign n753 = n268 & n476;
  assign n754 = i_13_ & n753;
  assign n755 = ~n752 & ~n754;
  assign n756 = ~n750 & n755;
  assign n757 = n305 & ~n756;
  assign n758 = n534 & n591;
  assign n759 = n512 & n758;
  assign n760 = ~n87 & n404;
  assign n761 = ~n212 & n700;
  assign n762 = n454 & n761;
  assign n763 = ~n760 & ~n762;
  assign n764 = ~n759 & n763;
  assign n765 = ~n757 & n764;
  assign n766 = n121 & ~n765;
  assign n767 = n747 & ~n766;
  assign n768 = n269 & n504;
  assign n769 = ~n414 & ~n462;
  assign n770 = n195 & ~n769;
  assign n771 = ~n768 & ~n770;
  assign n772 = ~i_25_ & i_26_;
  assign n773 = n502 & ~n772;
  assign n774 = n80 & n773;
  assign n775 = ~n198 & n367;
  assign n776 = n187 & n775;
  assign n777 = ~n774 & ~n776;
  assign n778 = ~i_39_ & ~n777;
  assign n779 = n370 & ~n778;
  assign n780 = n499 & ~n563;
  assign n781 = ~n513 & n780;
  assign n782 = n91 & n781;
  assign n783 = n779 & ~n782;
  assign n784 = n347 & n350;
  assign n785 = n171 & n197;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~i_40_ & ~n786;
  assign n788 = ~i_7_ & n510;
  assign n789 = n508 & n788;
  assign n790 = ~n434 & n789;
  assign n791 = ~i_15_ & n77;
  assign n792 = n448 & n791;
  assign n793 = i_37_ & n176;
  assign n794 = n283 & n793;
  assign n795 = n792 & n794;
  assign n796 = n244 & ~n400;
  assign n797 = n404 & n796;
  assign n798 = ~n795 & ~n797;
  assign n799 = ~n790 & n798;
  assign n800 = ~n787 & n799;
  assign n801 = n364 & n653;
  assign n802 = n177 & n445;
  assign n803 = i_39_ & n300;
  assign n804 = n802 & n803;
  assign n805 = n250 & n804;
  assign n806 = ~n801 & ~n805;
  assign n807 = i_40_ & ~n806;
  assign n808 = n179 & n351;
  assign n809 = i_31_ & n339;
  assign n810 = n510 & n809;
  assign n811 = n586 & n810;
  assign n812 = ~n808 & ~n811;
  assign n813 = ~n807 & n812;
  assign n814 = n800 & n813;
  assign n815 = n783 & n814;
  assign n816 = n771 & n815;
  assign n817 = n80 & n133;
  assign n818 = n559 & n817;
  assign n819 = n304 & n389;
  assign n820 = i_22_ & n91;
  assign n821 = ~i_21_ & n820;
  assign n822 = n526 & n821;
  assign n823 = ~n313 & ~n822;
  assign n824 = n97 & n279;
  assign n825 = ~n823 & n824;
  assign n826 = ~n819 & ~n825;
  assign n827 = ~n818 & n826;
  assign n828 = n816 & n827;
  assign o_4_ = ~n767 | ~n828;
  assign n830 = n166 & n524;
  assign n831 = n482 & n736;
  assign n832 = n93 & n675;
  assign n833 = n448 & n735;
  assign n834 = n201 & n578;
  assign n835 = ~i_34_ & n834;
  assign n836 = ~n833 & ~n835;
  assign n837 = ~n832 & n836;
  assign n838 = ~n831 & n837;
  assign n839 = n177 & ~n838;
  assign n840 = ~n830 & ~n839;
  assign n841 = i_40_ & ~n215;
  assign n842 = n217 & ~n841;
  assign n843 = ~n118 & ~n842;
  assign n844 = ~i_21_ & n119;
  assign n845 = ~n215 & ~n844;
  assign n846 = ~n843 & ~n845;
  assign n847 = n185 & n482;
  assign n848 = n80 & n847;
  assign n849 = ~n174 & ~n848;
  assign n850 = n124 & ~n591;
  assign n851 = n356 & n850;
  assign n852 = n122 & n489;
  assign n853 = ~n588 & n852;
  assign n854 = n214 & n853;
  assign n855 = ~n851 & ~n854;
  assign n856 = n849 & n855;
  assign n857 = ~n846 & n856;
  assign n858 = n304 & ~n503;
  assign n859 = n122 & n413;
  assign n860 = n230 & n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = n387 & n535;
  assign n863 = ~i_37_ & n547;
  assign n864 = ~n524 & ~n863;
  assign n865 = ~i_23_ & n79;
  assign n866 = n91 & n865;
  assign n867 = ~n864 & n866;
  assign n868 = ~n862 & ~n867;
  assign n869 = n861 & n868;
  assign n870 = n857 & n869;
  assign n871 = n840 & n870;
  assign n872 = n296 & n871;
  assign n873 = n151 & n351;
  assign n874 = ~i_13_ & n308;
  assign n875 = n80 & n445;
  assign n876 = ~n874 & ~n875;
  assign n877 = n133 & n216;
  assign n878 = ~n876 & n877;
  assign n879 = ~n159 & n418;
  assign n880 = n368 & ~n879;
  assign n881 = n241 & n307;
  assign n882 = i_36_ & n103;
  assign n883 = n339 & n882;
  assign n884 = ~n305 & n883;
  assign n885 = ~n881 & ~n884;
  assign n886 = n803 & ~n885;
  assign n887 = ~n880 & ~n886;
  assign n888 = ~n878 & n887;
  assign n889 = ~n873 & n888;
  assign n890 = i_40_ & ~n889;
  assign n891 = ~i_7_ & n677;
  assign n892 = n289 & n587;
  assign n893 = ~n298 & ~n892;
  assign n894 = ~n98 & ~n199;
  assign n895 = n195 & ~n894;
  assign n896 = n893 & ~n895;
  assign n897 = ~n891 & n896;
  assign n898 = n241 & n313;
  assign n899 = ~n171 & ~n898;
  assign n900 = n431 & ~n899;
  assign n901 = ~i_7_ & n204;
  assign n902 = n340 & n901;
  assign n903 = n170 & n902;
  assign n904 = ~i_38_ & n903;
  assign n905 = ~i_31_ & n444;
  assign n906 = n177 & n905;
  assign n907 = n373 & n906;
  assign n908 = ~n904 & ~n907;
  assign n909 = ~i_37_ & ~n908;
  assign n910 = n268 & ~n315;
  assign n911 = n91 & n910;
  assign n912 = n359 & n911;
  assign n913 = ~n909 & ~n912;
  assign n914 = ~n900 & n913;
  assign n915 = n897 & n914;
  assign n916 = n350 & n437;
  assign n917 = n902 & n916;
  assign n918 = ~i_31_ & n305;
  assign n919 = n283 & n918;
  assign n920 = n666 & n919;
  assign n921 = ~n917 & ~n920;
  assign n922 = ~n348 & ~n774;
  assign n923 = n921 & n922;
  assign n924 = ~i_22_ & ~i_36_;
  assign n925 = n119 & n924;
  assign n926 = n216 & n925;
  assign n927 = ~n259 & n926;
  assign n928 = n923 & ~n927;
  assign n929 = n915 & n928;
  assign n930 = ~n890 & n929;
  assign o_5_ = ~n872 | ~n930;
  assign n932 = n216 & n317;
  assign n933 = ~n180 & ~n932;
  assign n934 = ~i_34_ & n479;
  assign n935 = ~n933 & n934;
  assign n936 = ~n428 & ~n502;
  assign n937 = ~n476 & n936;
  assign n938 = n80 & ~n937;
  assign n939 = n280 & n525;
  assign n940 = n316 & n939;
  assign n941 = ~n848 & ~n940;
  assign n942 = ~n938 & n941;
  assign n943 = ~n935 & n942;
  assign n944 = ~n102 & ~n748;
  assign n945 = n307 & ~n944;
  assign n946 = n133 & n412;
  assign n947 = ~n96 & ~n173;
  assign n948 = ~n419 & n947;
  assign n949 = ~i_36_ & ~n948;
  assign n950 = ~n946 & ~n949;
  assign n951 = n313 & ~n950;
  assign n952 = ~n945 & ~n951;
  assign n953 = n228 & ~n952;
  assign n954 = ~i_40_ & n352;
  assign n955 = n300 & n503;
  assign n956 = ~n118 & ~n955;
  assign n957 = ~n876 & ~n956;
  assign n958 = n460 & n793;
  assign n959 = ~i_7_ & n409;
  assign n960 = n958 & n959;
  assign n961 = ~n410 & ~n958;
  assign n962 = n802 & ~n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~n957 & n963;
  assign n965 = ~n954 & n964;
  assign n966 = ~n953 & n965;
  assign n967 = n943 & n966;
  assign n968 = n351 & ~n717;
  assign n969 = ~i_35_ & n192;
  assign n970 = n919 & n969;
  assign n971 = ~n950 & n970;
  assign n972 = n170 & n460;
  assign n973 = i_37_ & n972;
  assign n974 = n316 & n973;
  assign n975 = ~n971 & ~n974;
  assign n976 = ~n968 & n975;
  assign n977 = n653 & n874;
  assign n978 = n151 & n171;
  assign n979 = ~n977 & ~n978;
  assign n980 = i_40_ & ~n979;
  assign n981 = ~n365 & n427;
  assign n982 = n250 & n906;
  assign n983 = i_11_ & n883;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~i_37_ & n460;
  assign n986 = ~n984 & n985;
  assign n987 = n195 & n356;
  assign n988 = n503 & n776;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~n986 & n989;
  assign n991 = ~n981 & n990;
  assign n992 = ~n980 & n991;
  assign n993 = n976 & n992;
  assign n994 = n158 & n269;
  assign n995 = ~i_36_ & n994;
  assign n996 = n434 & n995;
  assign n997 = n98 & n982;
  assign n998 = i_9_ & n278;
  assign n999 = ~n356 & ~n534;
  assign n1000 = n125 & ~n537;
  assign n1001 = ~n999 & n1000;
  assign n1002 = ~n998 & ~n1001;
  assign n1003 = ~n997 & n1002;
  assign n1004 = ~n996 & n1003;
  assign n1005 = n993 & n1004;
  assign n1006 = n410 & n526;
  assign n1007 = n371 & n1006;
  assign n1008 = n97 & n316;
  assign n1009 = ~i_37_ & n178;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = ~i_21_ & n162;
  assign n1012 = n95 & ~n1011;
  assign n1013 = ~n1010 & n1012;
  assign n1014 = ~n1007 & ~n1013;
  assign n1015 = i_22_ & ~n1014;
  assign n1016 = n1005 & ~n1015;
  assign o_6_ = ~n967 | ~n1016;
  assign n1018 = n464 & n969;
  assign n1019 = ~o_15_ & ~n1018;
  assign n1020 = n90 & n315;
  assign n1021 = n101 & n103;
  assign n1022 = n1020 & n1021;
  assign n1023 = n542 & n1022;
  assign n1024 = ~n550 & n1023;
  assign n1025 = n1019 & ~n1024;
  assign n1026 = ~n566 & n1025;
  assign n1027 = n172 & n542;
  assign n1028 = n557 & n1027;
  assign n1029 = i_38_ & n1028;
  assign n1030 = ~n718 & ~n1029;
  assign n1031 = n192 & ~n1030;
  assign n1032 = n104 & n118;
  assign n1033 = i_23_ & n101;
  assign n1034 = n1032 & n1033;
  assign n1035 = ~n106 & ~n360;
  assign n1036 = ~n1034 & n1035;
  assign n1037 = n1020 & ~n1036;
  assign n1038 = ~n150 & ~n460;
  assign n1039 = n683 & ~n1038;
  assign n1040 = n79 & n102;
  assign n1041 = n528 & n1040;
  assign n1042 = ~n1039 & ~n1041;
  assign n1043 = ~i_5_ & n591;
  assign n1044 = n241 & n1043;
  assign n1045 = ~n170 & ~n1044;
  assign n1046 = n179 & ~n1045;
  assign n1047 = n388 & n1043;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n1042 & n1048;
  assign n1050 = ~n1037 & n1049;
  assign n1051 = ~n1031 & n1050;
  assign o_7_ = ~n1026 | ~n1051;
  assign n1053 = n179 & n577;
  assign o_8_ = ~n1019 | n1053;
  assign n1055 = ~i_21_ & n1041;
  assign n1056 = n567 & ~n1047;
  assign o_9_ = n1055 | ~n1056;
  assign n1058 = ~i_20_ & ~i_25_;
  assign n1059 = ~i_40_ & n877;
  assign n1060 = ~n135 & ~n1059;
  assign n1061 = ~n102 & n1060;
  assign n1062 = n1021 & ~n1061;
  assign n1063 = i_35_ & n1062;
  assign n1064 = ~n939 & ~n972;
  assign n1065 = ~n1063 & n1064;
  assign n1066 = ~n1058 & ~n1065;
  assign n1067 = n316 & n1066;
  assign n1068 = ~n175 & ~n785;
  assign o_10_ = n1067 | ~n1068;
  assign n1070 = ~i_7_ & i_9_;
  assign n1071 = n565 & n1070;
  assign n1072 = ~n126 & n1071;
  assign n1073 = ~n272 & n400;
  assign n1074 = n91 & n564;
  assign n1075 = n1073 & n1074;
  assign n1076 = ~n818 & ~n1075;
  assign n1077 = ~n1072 & n1076;
  assign n1078 = ~i_7_ & n1043;
  assign n1079 = n392 & n1078;
  assign n1080 = n1068 & ~n1079;
  assign n1081 = ~n181 & n1080;
  assign o_11_ = ~n1077 | ~n1081;
  assign n1083 = i_5_ & ~i_7_;
  assign n1084 = ~i_0_ & n1083;
  assign n1085 = i_8_ & n1084;
  assign n1086 = ~i_40_ & n1085;
  assign n1087 = ~i_32_ & n1086;
  assign o_12_ = ~n338 & n1087;
  assign n1089 = ~n412 & ~n460;
  assign n1090 = n454 & ~n1089;
  assign n1091 = ~o_15_ & ~n1090;
  assign o_13_ = n531 | ~n1091;
  assign n1093 = ~i_13_ & n1091;
  assign o_14_ = o_13_ & ~n1093;
  assign n1095 = n177 & n547;
  assign n1096 = n793 & n1095;
  assign n1097 = i_40_ & n346;
  assign n1098 = ~n196 & ~n1097;
  assign n1099 = n151 & ~n1098;
  assign n1100 = i_0_ & n158;
  assign n1101 = ~n151 & ~n434;
  assign n1102 = n1100 & ~n1101;
  assign n1103 = ~n84 & ~n1102;
  assign n1104 = n195 & ~n1103;
  assign n1105 = n188 & n306;
  assign n1106 = n206 & n209;
  assign n1107 = n549 & n1106;
  assign n1108 = n203 & n1107;
  assign n1109 = ~n1105 & ~n1108;
  assign n1110 = ~n1104 & n1109;
  assign n1111 = ~n1099 & n1110;
  assign o_16_ = n1096 | ~n1111;
  assign n1113 = ~n492 & ~n587;
  assign n1114 = n126 & ~n1113;
  assign n1115 = n123 & n1114;
  assign n1116 = n276 & n865;
  assign n1117 = i_39_ & n618;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1115 & n1118;
  assign n1120 = n90 & ~n1119;
  assign n1121 = ~n388 & ~n535;
  assign n1122 = n537 & ~n1121;
  assign n1123 = ~i_5_ & n1122;
  assign n1124 = n644 & ~n1123;
  assign n1125 = ~n1120 & n1124;
  assign n1126 = ~n160 & n1125;
  assign n1127 = i_36_ & n677;
  assign n1128 = ~i_38_ & n681;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = n575 & ~n955;
  assign n1131 = n698 & ~n1130;
  assign n1132 = i_39_ & n350;
  assign n1133 = n242 & n1132;
  assign n1134 = n243 & n1133;
  assign n1135 = ~n1131 & ~n1134;
  assign n1136 = n1129 & n1135;
  assign n1137 = n237 & ~n275;
  assign n1138 = ~i_35_ & n667;
  assign n1139 = ~n1137 & n1138;
  assign n1140 = ~n116 & ~n251;
  assign n1141 = n169 & ~n400;
  assign n1142 = i_15_ & n1141;
  assign n1143 = ~n1140 & n1142;
  assign n1144 = ~n1139 & ~n1143;
  assign n1145 = n665 & ~n1144;
  assign n1146 = ~n715 & ~n1145;
  assign n1147 = n123 & ~n1146;
  assign n1148 = ~n297 & n690;
  assign n1149 = n117 & n638;
  assign n1150 = n203 & n578;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1148 & n1151;
  assign n1153 = ~n1147 & n1152;
  assign n1154 = n1136 & n1153;
  assign o_17_ = ~n1126 | ~n1154;
  assign n1156 = ~i_39_ & n198;
  assign n1157 = ~n274 & ~n355;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = n178 & n1100;
  assign n1160 = ~i_11_ & n96;
  assign n1161 = ~n350 & n389;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1159 & n1162;
  assign n1164 = ~n1158 & n1163;
  assign n1165 = n195 & ~n1164;
  assign n1166 = n427 & ~n876;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n178 & ~n475;
  assign n1169 = n94 & ~n1168;
  assign n1170 = ~n360 & ~n1169;
  assign n1171 = n316 & ~n1170;
  assign n1172 = ~n175 & ~n1171;
  assign n1173 = ~n784 & n1172;
  assign n1174 = n350 & ~n1098;
  assign n1175 = ~n746 & ~n1174;
  assign n1176 = n1173 & n1175;
  assign n1177 = n1167 & n1176;
  assign n1178 = ~n151 & ~n675;
  assign n1179 = n346 & ~n1178;
  assign n1180 = i_40_ & ~n418;
  assign n1181 = ~n208 & ~n1180;
  assign n1182 = n995 & n1181;
  assign n1183 = i_32_ & n788;
  assign n1184 = n708 & n1106;
  assign n1185 = n692 & n1184;
  assign n1186 = ~n1183 & ~n1185;
  assign n1187 = ~n1182 & n1186;
  assign n1188 = ~n1179 & n1187;
  assign n1189 = ~n150 & ~n345;
  assign n1190 = ~i_31_ & n510;
  assign n1191 = n121 & n1190;
  assign n1192 = ~n274 & ~n537;
  assign n1193 = n1191 & n1192;
  assign n1194 = ~n171 & ~n1193;
  assign n1195 = ~n1189 & ~n1194;
  assign n1196 = n1188 & ~n1195;
  assign n1197 = n1177 & n1196;
  assign n1198 = n103 & n515;
  assign n1199 = ~n1113 & n1198;
  assign n1200 = ~i_7_ & n1199;
  assign n1201 = n83 & n303;
  assign n1202 = ~i_35_ & n504;
  assign n1203 = i_38_ & n736;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = n177 & ~n1204;
  assign n1206 = ~n1201 & ~n1205;
  assign n1207 = ~n1200 & n1206;
  assign n1208 = n273 & n274;
  assign n1209 = ~n1132 & ~n1208;
  assign n1210 = i_9_ & ~n1209;
  assign n1211 = n150 & n297;
  assign n1212 = ~n89 & ~n229;
  assign n1213 = ~n300 & n1089;
  assign n1214 = n1212 & ~n1213;
  assign n1215 = ~n955 & ~n1214;
  assign n1216 = ~n1211 & n1215;
  assign n1217 = ~n1210 & n1216;
  assign n1218 = n1191 & ~n1217;
  assign n1219 = n1207 & ~n1218;
  assign n1220 = n943 & n1219;
  assign o_18_ = ~n1197 | ~n1220;
  assign n1222 = ~n172 & n300;
  assign n1223 = n170 & n1222;
  assign n1224 = ~n916 & ~n1223;
  assign n1225 = ~i_2_ & n301;
  assign n1226 = n901 & n1225;
  assign n1227 = ~n1224 & n1226;
  assign n1228 = n414 & n437;
  assign n1229 = i_40_ & n1132;
  assign n1230 = n336 & n1229;
  assign n1231 = ~n97 & ~n434;
  assign n1232 = n882 & ~n1231;
  assign n1233 = i_35_ & n1232;
  assign n1234 = ~n1230 & ~n1233;
  assign n1235 = i_6_ & ~i_32_;
  assign n1236 = ~n1234 & n1235;
  assign n1237 = ~n1228 & ~n1236;
  assign n1238 = ~n1090 & n1237;
  assign n1239 = ~i_7_ & ~n1238;
  assign n1240 = n216 & n297;
  assign n1241 = ~n195 & ~n995;
  assign n1242 = n1240 & ~n1241;
  assign n1243 = ~n1239 & ~n1242;
  assign o_19_ = n1227 | ~n1243;
  assign n1245 = n335 & n414;
  assign n1246 = ~n1032 & ~n1245;
  assign n1247 = n372 & n389;
  assign n1248 = n479 & n549;
  assign n1249 = ~i_36_ & n1248;
  assign n1250 = ~n309 & ~n1249;
  assign n1251 = n169 & n419;
  assign n1252 = ~n413 & ~n1251;
  assign n1253 = n1250 & n1252;
  assign n1254 = i_9_ & n118;
  assign n1255 = ~i_40_ & ~n1254;
  assign n1256 = ~n267 & ~n1255;
  assign n1257 = n1253 & ~n1256;
  assign n1258 = ~n1247 & n1257;
  assign n1259 = n103 & ~n1258;
  assign n1260 = n1246 & ~n1259;
  assign n1261 = ~i_15_ & n339;
  assign n1262 = ~n1260 & n1261;
  assign n1263 = i_14_ & ~n1073;
  assign n1264 = n780 & ~n1263;
  assign n1265 = n403 & n863;
  assign n1266 = ~n267 & n512;
  assign n1267 = ~n126 & n1266;
  assign n1268 = ~n1265 & ~n1267;
  assign n1269 = i_9_ & ~i_12_;
  assign n1270 = ~n1268 & n1269;
  assign n1271 = ~n190 & ~n405;
  assign n1272 = ~n1270 & n1271;
  assign n1273 = ~n1264 & n1272;
  assign n1274 = ~i_7_ & ~n1273;
  assign n1275 = n234 & n274;
  assign n1276 = ~n152 & ~n1275;
  assign n1277 = n1084 & ~n1276;
  assign n1278 = n218 & ~n479;
  assign n1279 = ~n135 & ~n1278;
  assign n1280 = n1253 & n1279;
  assign n1281 = n306 & ~n1280;
  assign n1282 = ~n1277 & ~n1281;
  assign n1283 = n192 & ~n1282;
  assign n1284 = n240 & n1222;
  assign n1285 = ~n916 & ~n1284;
  assign n1286 = ~n148 & n1285;
  assign n1287 = n1084 & ~n1286;
  assign n1288 = ~i_32_ & n1083;
  assign n1289 = n509 & n1288;
  assign n1290 = n84 & n1289;
  assign n1291 = n78 & n218;
  assign n1292 = i_33_ & n1291;
  assign n1293 = n1246 & ~n1292;
  assign n1294 = n1288 & ~n1293;
  assign n1295 = ~n1290 & ~n1294;
  assign n1296 = ~n1287 & n1295;
  assign n1297 = ~i_11_ & n1070;
  assign n1298 = ~n1268 & n1297;
  assign n1299 = n77 & n415;
  assign n1300 = ~n280 & ~n1299;
  assign n1301 = n306 & ~n1300;
  assign n1302 = ~n117 & ~n251;
  assign n1303 = n274 & n809;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n403 & n1083;
  assign n1306 = ~n810 & ~n1305;
  assign n1307 = ~n1304 & ~n1306;
  assign n1308 = n863 & n1289;
  assign n1309 = n402 & n1305;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1307 & n1310;
  assign n1312 = ~n1301 & n1311;
  assign n1313 = ~n1298 & n1312;
  assign n1314 = n1296 & n1313;
  assign n1315 = ~n1283 & n1314;
  assign n1316 = ~n1274 & n1315;
  assign o_20_ = n1262 | ~n1316;
  assign n1318 = n78 & n145;
  assign n1319 = n251 & n1318;
  assign n1320 = ~n735 & ~n793;
  assign n1321 = n134 & ~n1320;
  assign n1322 = ~n1319 & ~n1321;
  assign n1323 = ~i_6_ & ~n1322;
  assign n1324 = i_32_ & ~n169;
  assign n1325 = n202 & n549;
  assign n1326 = ~i_0_ & n1325;
  assign n1327 = ~n1324 & ~n1326;
  assign n1328 = ~i_34_ & ~n1327;
  assign n1329 = i_33_ & ~n176;
  assign n1330 = ~n1202 & n1329;
  assign n1331 = ~n77 & ~n1330;
  assign n1332 = ~n1328 & ~n1331;
  assign n1333 = ~n147 & ~n153;
  assign n1334 = n176 & n1222;
  assign n1335 = n318 & n547;
  assign n1336 = ~n333 & ~n1335;
  assign n1337 = ~n1334 & n1336;
  assign n1338 = n1333 & n1337;
  assign n1339 = ~i_0_ & ~i_5_;
  assign n1340 = ~n1338 & n1339;
  assign n1341 = n1332 & ~n1340;
  assign n1342 = ~n1323 & n1341;
  assign o_21_ = ~o_15_ & ~n1342;
  assign n1344 = ~i_7_ & ~n1216;
  assign n1345 = n273 & n1070;
  assign n1346 = n430 & n1345;
  assign n1347 = ~n1344 & ~n1346;
  assign n1348 = n1190 & ~n1347;
  assign n1349 = n1296 & ~n1348;
  assign n1350 = ~n216 & ~n434;
  assign n1351 = n515 & ~n1350;
  assign n1352 = n510 & ~n1351;
  assign n1353 = i_37_ & n192;
  assign n1354 = ~i_0_ & n1353;
  assign n1355 = ~i_35_ & ~n179;
  assign n1356 = i_35_ & ~n547;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = n1354 & n1357;
  assign n1359 = ~n1352 & ~n1358;
  assign n1360 = n1083 & ~n1359;
  assign n1361 = ~n1183 & ~n1360;
  assign o_22_ = ~n1349 | ~n1361;
  assign n1363 = i_37_ & ~n158;
  assign n1364 = ~n341 & ~n1363;
  assign n1365 = n372 & ~n1364;
  assign n1366 = ~n172 & n390;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n168 & ~n1367;
  assign n1369 = i_35_ & ~n418;
  assign n1370 = ~n274 & n1369;
  assign n1371 = ~n653 & ~n1370;
  assign n1372 = n192 & ~n1371;
  assign n1373 = ~n172 & n1372;
  assign n1374 = ~n1368 & ~n1373;
  assign n1375 = ~i_0_ & i_5_;
  assign n1376 = n300 & n1375;
  assign n1377 = n178 & ~n355;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~i_36_ & ~n1378;
  assign n1380 = ~n504 & ~n1379;
  assign n1381 = n149 & ~n1380;
  assign n1382 = ~n96 & n1157;
  assign n1383 = n194 & ~n1382;
  assign n1384 = ~i_9_ & n116;
  assign n1385 = ~i_31_ & ~n1384;
  assign n1386 = ~i_5_ & n1385;
  assign n1387 = n403 & ~n1386;
  assign n1388 = ~n1383 & ~n1387;
  assign n1389 = ~n1381 & n1388;
  assign n1390 = n302 & n683;
  assign n1391 = ~n280 & ~n360;
  assign n1392 = ~n1390 & n1391;
  assign n1393 = n250 & n792;
  assign n1394 = ~n676 & ~n1393;
  assign n1395 = n1392 & n1394;
  assign n1396 = n1389 & n1395;
  assign n1397 = n1374 & n1396;
  assign n1398 = n318 & n341;
  assign n1399 = n411 & ~n1212;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n77 & ~n1400;
  assign n1402 = ~n969 & ~n1354;
  assign n1403 = i_5_ & ~n1402;
  assign n1404 = i_0_ & n194;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1401 & n1405;
  assign n1407 = i_38_ & ~n1406;
  assign n1408 = n96 & ~n1212;
  assign n1409 = ~i_38_ & n305;
  assign n1410 = ~n229 & ~n1409;
  assign n1411 = n234 & ~n1410;
  assign n1412 = ~n1408 & ~n1411;
  assign n1413 = n969 & ~n1412;
  assign n1414 = ~n570 & ~n624;
  assign n1415 = ~o_15_ & n1414;
  assign n1416 = ~n1413 & n1415;
  assign n1417 = ~n691 & n1416;
  assign n1418 = ~n449 & n577;
  assign n1419 = n465 & ~n547;
  assign n1420 = n302 & n350;
  assign n1421 = ~n502 & ~n1420;
  assign n1422 = ~n863 & n1421;
  assign n1423 = ~n1419 & n1422;
  assign n1424 = n79 & ~n1423;
  assign n1425 = ~n1418 & ~n1424;
  assign n1426 = n1417 & n1425;
  assign n1427 = ~n1407 & n1426;
  assign o_23_ = ~n1397 | ~n1427;
  assign n1429 = n289 & ~n563;
  assign n1430 = i_40_ & n830;
  assign n1431 = n670 & n1059;
  assign n1432 = n214 & n1431;
  assign n1433 = ~n1430 & ~n1432;
  assign n1434 = ~n1429 & n1433;
  assign n1435 = n90 & n111;
  assign n1436 = n339 & n1435;
  assign n1437 = n105 & n1436;
  assign n1438 = ~n322 & ~n1437;
  assign n1439 = ~i_21_ & n325;
  assign n1440 = n1438 & ~n1439;
  assign n1441 = n257 & n1440;
  assign n1442 = n1434 & n1441;
  assign n1443 = n137 & n1431;
  assign n1444 = ~n357 & ~n1443;
  assign n1445 = ~n299 & n1444;
  assign n1446 = n266 & n1445;
  assign n1447 = i_40_ & n476;
  assign n1448 = n911 & n1447;
  assign n1449 = n925 & ~n1130;
  assign n1450 = n276 & ~n620;
  assign n1451 = n119 & n1450;
  assign n1452 = ~n1449 & ~n1451;
  assign n1453 = ~n1448 & n1452;
  assign n1454 = n1446 & n1453;
  assign n1455 = n121 & n1122;
  assign n1456 = n1454 & ~n1455;
  assign n1457 = ~n768 & n1456;
  assign n1458 = n1442 & n1457;
  assign n1459 = ~n161 & ~n271;
  assign n1460 = ~n172 & ~n355;
  assign n1461 = n904 & n1460;
  assign o_32_ = n346 & n1211;
  assign n1463 = ~n917 & ~o_32_;
  assign n1464 = ~n1461 & n1463;
  assign n1465 = n224 & n1464;
  assign n1466 = n1459 & n1465;
  assign o_24_ = ~n1458 | ~n1466;
  assign n1468 = n902 & ~n1224;
  assign o_28_ = n200 | n1468;
  assign n1470 = ~n222 & ~o_28_;
  assign o_25_ = ~n1458 | ~n1470;
  assign n1472 = ~i_39_ & n211;
  assign n1473 = ~n768 & ~n1472;
  assign o_26_ = ~n1459 | ~n1473;
  assign n1475 = ~n222 & n1442;
  assign o_27_ = ~n1454 | ~n1475;
  assign n1477 = n92 & n376;
  assign n1478 = ~n973 & ~n1477;
  assign n1479 = n821 & ~n1478;
  assign n1480 = ~n357 & ~n1479;
  assign o_29_ = n1455 | ~n1480;
  assign n1482 = n111 & n165;
  assign n1483 = n105 & n1482;
  assign n1484 = ~n315 & n1249;
  assign n1485 = i_35_ & n924;
  assign n1486 = ~n575 & n1485;
  assign n1487 = n621 & n1275;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1484 & n1488;
  assign n1490 = n103 & ~n1489;
  assign n1491 = ~n1483 & ~n1490;
  assign n1492 = n329 & ~n1491;
  assign n1493 = ~n200 & ~n1448;
  assign o_30_ = n1492 | ~n1493;
  assign n1495 = ~n264 & n1470;
  assign n1496 = n820 & n1040;
  assign n1497 = n1482 & n1496;
  assign n1498 = n316 & n1116;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n299 & n1499;
  assign o_31_ = ~n1495 | ~n1500;
  assign n1502 = n169 & ~n948;
  assign n1503 = n905 & n1502;
  assign n1504 = n202 & n460;
  assign n1505 = n445 & n1248;
  assign n1506 = n469 & n549;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1504 & n1507;
  assign n1509 = ~n1028 & n1508;
  assign n1510 = ~n1503 & n1509;
  assign n1511 = n192 & ~n1510;
  assign n1512 = n185 & n619;
  assign n1513 = i_32_ & ~i_33_;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = n666 & n905;
  assign n1516 = n1514 & ~n1515;
  assign n1517 = ~o_13_ & n1516;
  assign n1518 = n435 & n1240;
  assign n1519 = n572 & ~n1518;
  assign n1520 = n1517 & n1519;
  assign n1521 = ~n1511 & n1520;
  assign n1522 = ~i_5_ & n400;
  assign n1523 = ~n513 & n1522;
  assign n1524 = n564 & n1523;
  assign n1525 = ~n1040 & n1391;
  assign n1526 = n445 & ~n1525;
  assign n1527 = n475 & n1318;
  assign n1528 = n178 & ~n1320;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = i_33_ & n1235;
  assign n1531 = ~n1529 & n1530;
  assign n1532 = n242 & ~n948;
  assign n1533 = ~n859 & ~n1532;
  assign n1534 = n407 & ~n1533;
  assign n1535 = ~n1531 & ~n1534;
  assign n1536 = ~n1526 & n1535;
  assign n1537 = ~n1524 & n1536;
  assign n1538 = n1050 & n1537;
  assign n1539 = ~i_5_ & i_9_;
  assign n1540 = n228 & n863;
  assign n1541 = ~n273 & n1540;
  assign n1542 = n251 & n510;
  assign n1543 = ~i_40_ & n272;
  assign n1544 = ~n1542 & n1543;
  assign n1545 = ~n126 & ~n1140;
  assign n1546 = ~n513 & n1545;
  assign n1547 = ~n1544 & n1546;
  assign n1548 = n242 & n1547;
  assign n1549 = ~n1133 & ~n1548;
  assign n1550 = ~n1541 & n1549;
  assign n1551 = n1539 & ~n1550;
  assign n1552 = n573 & ~n575;
  assign n1553 = n189 & ~n305;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1027 & ~n1248;
  assign n1556 = n1022 & ~n1555;
  assign n1557 = n78 & n955;
  assign n1558 = ~n374 & ~n1557;
  assign n1559 = n409 & ~n1558;
  assign n1560 = ~n1556 & ~n1559;
  assign n1561 = n1554 & n1560;
  assign n1562 = ~n338 & n1225;
  assign n1563 = n549 & n882;
  assign n1564 = i_0_ & n205;
  assign n1565 = n1563 & n1564;
  assign n1566 = i_35_ & n1565;
  assign n1567 = ~n1562 & ~n1566;
  assign n1568 = n632 & ~n1567;
  assign n1569 = n1561 & ~n1568;
  assign n1570 = ~n1551 & n1569;
  assign n1571 = n1538 & n1570;
  assign o_33_ = ~n1521 | ~n1571;
  assign n1573 = i_36_ & n117;
  assign n1574 = ~n152 & ~n1573;
  assign n1575 = n1100 & ~n1574;
  assign n1576 = ~n516 & ~n1575;
  assign n1577 = n132 & ~n1576;
  assign n1578 = n169 & ~n251;
  assign n1579 = ~n220 & ~n1578;
  assign n1580 = ~i_34_ & ~n1579;
  assign n1581 = n250 & ~n514;
  assign n1582 = ~n415 & ~n1581;
  assign n1583 = ~n1580 & n1582;
  assign n1584 = ~n1291 & n1583;
  assign n1585 = i_5_ & ~n1584;
  assign n1586 = n193 & n863;
  assign n1587 = ~n946 & ~n1502;
  assign n1588 = n918 & ~n1587;
  assign n1589 = i_5_ & ~n401;
  assign n1590 = n1141 & n1589;
  assign n1591 = ~n1506 & ~n1590;
  assign n1592 = ~n1588 & n1591;
  assign n1593 = ~n1586 & n1592;
  assign n1594 = ~i_34_ & ~n1593;
  assign n1595 = ~n1585 & ~n1594;
  assign n1596 = ~n1577 & n1595;
  assign n1597 = ~i_34_ & ~n1276;
  assign n1598 = ~n146 & ~n333;
  assign n1599 = ~n1597 & n1598;
  assign n1600 = n169 & n1222;
  assign n1601 = n1599 & ~n1600;
  assign n1602 = n1375 & ~n1601;
  assign n1603 = n1596 & ~n1602;
  assign n1604 = n77 & ~n1603;
  assign n1605 = ~n1302 & n1318;
  assign n1606 = n134 & n793;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n1530 & ~n1607;
  assign n1609 = n251 & ~n513;
  assign n1610 = ~n434 & ~n1609;
  assign n1611 = n242 & ~n1610;
  assign n1612 = ~n402 & n1611;
  assign n1613 = n170 & n1211;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = ~n1608 & n1614;
  assign n1616 = ~n272 & n1540;
  assign n1617 = ~i_15_ & ~i_31_;
  assign n1618 = n235 & n1617;
  assign n1619 = n969 & n1618;
  assign n1620 = ~n1616 & ~n1619;
  assign n1621 = i_9_ & ~n1620;
  assign n1622 = ~n190 & n1091;
  assign n1623 = ~n1621 & n1622;
  assign n1624 = n1615 & n1623;
  assign n1625 = ~n803 & n947;
  assign n1626 = n510 & ~n1625;
  assign n1627 = n431 & n509;
  assign n1628 = ~n1542 & ~n1627;
  assign n1629 = ~n1626 & n1628;
  assign n1630 = n1617 & ~n1629;
  assign n1631 = n172 & ~n334;
  assign n1632 = n1562 & ~n1631;
  assign n1633 = i_37_ & n1565;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = n204 & ~n1634;
  assign n1636 = ~n1630 & ~n1635;
  assign n1637 = ~i_32_ & ~n1636;
  assign n1638 = n1624 & ~n1637;
  assign o_34_ = n1604 | ~n1638;
endmodule


