// Benchmark "t481" written by ABC on Tue May 16 16:07:52 2017

module t481 ( 
    v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9,
    \v16.0   );
  input  v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7,
    v8, v9;
  output \v16.0 ;
  wire n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132;
  assign n18 = v10 & v9;
  assign n19 = ~v12 & v15;
  assign n20 = v13 & n19;
  assign n21 = ~v5 & ~v8;
  assign n22 = v7 & n21;
  assign n23 = ~v3 & n22;
  assign n24 = v2 & n23;
  assign n25 = v0 & n24;
  assign n26 = n20 & n25;
  assign n27 = ~v11 & n26;
  assign n28 = n18 & n27;
  assign n29 = ~v1 & n23;
  assign n30 = v2 & n29;
  assign n31 = n20 & n30;
  assign n32 = ~v11 & n31;
  assign n33 = n18 & n32;
  assign n34 = v5 & v6;
  assign n35 = v0 & v2;
  assign n36 = ~v3 & n35;
  assign n37 = ~v4 & n36;
  assign n38 = ~v8 & v9;
  assign n39 = ~v11 & n38;
  assign n40 = v10 & n39;
  assign n41 = v15 & n40;
  assign n42 = ~v12 & n41;
  assign n43 = v13 & n42;
  assign n44 = n37 & n43;
  assign n45 = ~v7 & n44;
  assign n46 = n34 & n45;
  assign n47 = ~v1 & v2;
  assign n48 = ~v3 & n47;
  assign n49 = ~v4 & n48;
  assign n50 = ~v7 & n49;
  assign n51 = v6 & n50;
  assign n52 = v5 & n51;
  assign n53 = n43 & n52;
  assign n54 = ~n46 & ~n53;
  assign n55 = ~n33 & n54;
  assign n56 = ~n28 & n55;
  assign n57 = ~v6 & ~v8;
  assign n58 = v4 & n57;
  assign n59 = ~v3 & n58;
  assign n60 = v2 & n59;
  assign n61 = v0 & n60;
  assign n62 = n20 & n61;
  assign n63 = ~v11 & n62;
  assign n64 = n18 & n63;
  assign n65 = ~v1 & n59;
  assign n66 = v2 & n65;
  assign n67 = n20 & n66;
  assign n68 = ~v11 & n67;
  assign n69 = n18 & n68;
  assign n70 = ~v6 & n21;
  assign n71 = ~v3 & n70;
  assign n72 = v2 & n71;
  assign n73 = v0 & n72;
  assign n74 = n20 & n73;
  assign n75 = ~v11 & n74;
  assign n76 = n18 & n75;
  assign n77 = ~v1 & n71;
  assign n78 = v2 & n77;
  assign n79 = n20 & n78;
  assign n80 = ~v11 & n79;
  assign n81 = n18 & n80;
  assign n82 = ~n76 & ~n81;
  assign n83 = ~n69 & n82;
  assign n84 = ~n64 & n83;
  assign n85 = ~v0 & v1;
  assign n86 = ~v4 & n85;
  assign n87 = v3 & n86;
  assign n88 = ~v14 & n40;
  assign n89 = ~v12 & n88;
  assign n90 = v13 & n89;
  assign n91 = n87 & n90;
  assign n92 = ~v7 & n91;
  assign n93 = n34 & n92;
  assign n94 = ~v12 & v13;
  assign n95 = ~v2 & n85;
  assign n96 = ~v4 & n95;
  assign n97 = ~v7 & n96;
  assign n98 = v6 & n97;
  assign n99 = v5 & n98;
  assign n100 = n40 & n99;
  assign n101 = ~v14 & n100;
  assign n102 = n94 & n101;
  assign n103 = ~v12 & ~v14;
  assign n104 = v13 & n103;
  assign n105 = ~v2 & n70;
  assign n106 = ~v0 & n105;
  assign n107 = v1 & n106;
  assign n108 = n104 & n107;
  assign n109 = ~v11 & n108;
  assign n110 = n18 & n109;
  assign n111 = ~v11 & v9;
  assign n112 = v10 & n111;
  assign n113 = ~v14 & n112;
  assign n114 = ~v12 & n113;
  assign n115 = v13 & n114;
  assign n116 = v7 & ~v8;
  assign n117 = v4 & n116;
  assign n118 = v3 & n117;
  assign n119 = ~v0 & n118;
  assign n120 = v1 & n119;
  assign n121 = n115 & n120;
  assign n122 = v15 & n112;
  assign n123 = ~v12 & n122;
  assign n124 = v13 & n123;
  assign n125 = ~v3 & n117;
  assign n126 = v2 & n125;
  assign n127 = v0 & n126;
  assign n128 = n124 & n127;
  assign n129 = ~v1 & n125;
  assign n130 = v2 & n129;
  assign n131 = n124 & n130;
  assign n132 = ~v2 & n117;
  assign n133 = ~v0 & n132;
  assign n134 = v1 & n133;
  assign n135 = n115 & n134;
  assign n136 = ~n131 & ~n135;
  assign n137 = ~n128 & n136;
  assign n138 = ~n121 & n137;
  assign n139 = ~n110 & n138;
  assign n140 = ~n102 & n139;
  assign n141 = ~n93 & n140;
  assign n142 = ~v1 & ~v3;
  assign n143 = v2 & n142;
  assign n144 = n115 & n143;
  assign n145 = n58 & n144;
  assign n146 = v2 & ~v3;
  assign n147 = v0 & n146;
  assign n148 = ~v8 & n147;
  assign n149 = ~v5 & n148;
  assign n150 = ~v6 & n149;
  assign n151 = n115 & n150;
  assign n152 = n70 & n144;
  assign n153 = n22 & n115;
  assign n154 = v3 & n153;
  assign n155 = n85 & n154;
  assign n156 = ~n152 & ~n155;
  assign n157 = ~n151 & n156;
  assign n158 = ~n145 & n157;
  assign n159 = ~v0 & ~v2;
  assign n160 = v1 & n159;
  assign n161 = n115 & n160;
  assign n162 = n22 & n161;
  assign n163 = n58 & n115;
  assign n164 = v3 & n163;
  assign n165 = n85 & n164;
  assign n166 = n58 & n161;
  assign n167 = n70 & n115;
  assign n168 = v3 & n167;
  assign n169 = n85 & n168;
  assign n170 = ~n166 & ~n169;
  assign n171 = ~n165 & n170;
  assign n172 = ~n162 & n171;
  assign n173 = n115 & n130;
  assign n174 = v7 & n149;
  assign n175 = n115 & n174;
  assign n176 = n115 & n127;
  assign n177 = n30 & n104;
  assign n178 = ~v11 & n177;
  assign n179 = n18 & n178;
  assign n180 = n37 & n90;
  assign n181 = ~v7 & n180;
  assign n182 = n34 & n181;
  assign n183 = n40 & n52;
  assign n184 = ~v14 & n183;
  assign n185 = n94 & n184;
  assign n186 = n61 & n104;
  assign n187 = ~v11 & n186;
  assign n188 = n18 & n187;
  assign n189 = ~n185 & ~n188;
  assign n190 = ~n182 & n189;
  assign n191 = ~n179 & n190;
  assign n192 = ~n176 & n191;
  assign n193 = ~n175 & n192;
  assign n194 = ~n173 & n193;
  assign n195 = n172 & n194;
  assign n196 = n158 & n195;
  assign n197 = n141 & n196;
  assign n198 = n84 & n197;
  assign n199 = n56 & n198;
  assign n200 = n43 & n99;
  assign n201 = ~v0 & v3;
  assign n202 = v1 & n201;
  assign n203 = ~v8 & n202;
  assign n204 = v7 & n203;
  assign n205 = v4 & n204;
  assign n206 = n20 & n205;
  assign n207 = ~v11 & n206;
  assign n208 = n18 & n207;
  assign n209 = ~v8 & n160;
  assign n210 = v7 & n209;
  assign n211 = v4 & n210;
  assign n212 = n20 & n211;
  assign n213 = ~v11 & n212;
  assign n214 = n18 & n213;
  assign n215 = ~v10 & ~v12;
  assign n216 = v8 & n215;
  assign n217 = v7 & n147;
  assign n218 = v4 & n217;
  assign n219 = n216 & n218;
  assign n220 = ~v14 & n219;
  assign n221 = v13 & n220;
  assign n222 = ~n214 & ~n221;
  assign n223 = ~n208 & n222;
  assign n224 = ~n200 & n223;
  assign n225 = v7 & n143;
  assign n226 = v4 & n225;
  assign n227 = n216 & n226;
  assign n228 = ~v14 & n227;
  assign n229 = v13 & n228;
  assign n230 = ~v14 & n216;
  assign n231 = v13 & n230;
  assign n232 = n147 & n231;
  assign n233 = ~v5 & n232;
  assign n234 = v7 & n233;
  assign n235 = n143 & n231;
  assign n236 = ~v5 & n235;
  assign n237 = v7 & n236;
  assign n238 = ~v4 & v6;
  assign n239 = v5 & n238;
  assign n240 = ~v10 & ~v7;
  assign n241 = v8 & n240;
  assign n242 = ~v14 & n241;
  assign n243 = ~v12 & n242;
  assign n244 = v13 & n243;
  assign n245 = n239 & n244;
  assign n246 = ~v3 & n245;
  assign n247 = n35 & n246;
  assign n248 = ~n237 & ~n247;
  assign n249 = ~n234 & n248;
  assign n250 = ~n229 & n249;
  assign n251 = ~v2 & n22;
  assign n252 = ~v0 & n251;
  assign n253 = v1 & n252;
  assign n254 = n20 & n253;
  assign n255 = ~v11 & n254;
  assign n256 = n18 & n255;
  assign n257 = v3 & n58;
  assign n258 = ~v0 & n257;
  assign n259 = v1 & n258;
  assign n260 = n20 & n259;
  assign n261 = ~v11 & n260;
  assign n262 = n18 & n261;
  assign n263 = v3 & n22;
  assign n264 = ~v0 & n263;
  assign n265 = v1 & n264;
  assign n266 = n20 & n265;
  assign n267 = ~v11 & n266;
  assign n268 = n18 & n267;
  assign n269 = n124 & n160;
  assign n270 = n58 & n269;
  assign n271 = n70 & n124;
  assign n272 = v3 & n271;
  assign n273 = n85 & n272;
  assign n274 = n70 & n269;
  assign n275 = ~v7 & n87;
  assign n276 = v6 & n275;
  assign n277 = v5 & n276;
  assign n278 = n40 & n277;
  assign n279 = v15 & n278;
  assign n280 = n94 & n279;
  assign n281 = ~n274 & ~n280;
  assign n282 = ~n273 & n281;
  assign n283 = ~n270 & n282;
  assign n284 = ~n268 & n283;
  assign n285 = ~n262 & n284;
  assign n286 = ~n256 & n285;
  assign n287 = ~v6 & n36;
  assign n288 = v4 & n287;
  assign n289 = n216 & n288;
  assign n290 = ~v14 & n289;
  assign n291 = v13 & n290;
  assign n292 = v4 & ~v6;
  assign n293 = ~v3 & n292;
  assign n294 = ~v1 & n293;
  assign n295 = v2 & n294;
  assign n296 = n216 & n295;
  assign n297 = ~v14 & n296;
  assign n298 = v13 & n297;
  assign n299 = ~v3 & n239;
  assign n300 = ~v1 & n299;
  assign n301 = v2 & n300;
  assign n302 = n241 & n301;
  assign n303 = n104 & n302;
  assign n304 = ~n298 & ~n303;
  assign n305 = ~n291 & n304;
  assign n306 = ~v5 & n36;
  assign n307 = ~v6 & n306;
  assign n308 = n216 & n307;
  assign n309 = ~v14 & n308;
  assign n310 = v13 & n309;
  assign n311 = ~v5 & n48;
  assign n312 = ~v6 & n311;
  assign n313 = n216 & n312;
  assign n314 = ~v14 & n313;
  assign n315 = v13 & n314;
  assign n316 = ~v5 & n202;
  assign n317 = v7 & n316;
  assign n318 = n216 & n317;
  assign n319 = ~v14 & n318;
  assign n320 = v13 & n319;
  assign n321 = ~v5 & v7;
  assign n322 = ~v2 & n321;
  assign n323 = ~v0 & n322;
  assign n324 = v1 & n323;
  assign n325 = n216 & n324;
  assign n326 = ~v14 & n325;
  assign n327 = v13 & n326;
  assign n328 = ~n320 & ~n327;
  assign n329 = ~n315 & n328;
  assign n330 = ~n310 & n329;
  assign n331 = ~v6 & n202;
  assign n332 = v4 & n331;
  assign n333 = n216 & n332;
  assign n334 = ~v14 & n333;
  assign n335 = v13 & n334;
  assign n336 = ~v2 & n292;
  assign n337 = ~v0 & n336;
  assign n338 = v1 & n337;
  assign n339 = n216 & n338;
  assign n340 = ~v14 & n339;
  assign n341 = v13 & n340;
  assign n342 = ~v6 & n316;
  assign n343 = n216 & n342;
  assign n344 = ~v14 & n343;
  assign n345 = v13 & n344;
  assign n346 = ~v5 & n95;
  assign n347 = ~v6 & n346;
  assign n348 = n216 & n347;
  assign n349 = ~v14 & n348;
  assign n350 = v13 & n349;
  assign n351 = ~n345 & ~n350;
  assign n352 = ~n341 & n351;
  assign n353 = ~n335 & n352;
  assign n354 = v3 & n239;
  assign n355 = ~v0 & n354;
  assign n356 = v1 & n355;
  assign n357 = n241 & n356;
  assign n358 = n104 & n357;
  assign n359 = ~v2 & n239;
  assign n360 = ~v0 & n359;
  assign n361 = v1 & n360;
  assign n362 = n241 & n361;
  assign n363 = n104 & n362;
  assign n364 = v4 & v7;
  assign n365 = v3 & n364;
  assign n366 = ~v0 & n365;
  assign n367 = v1 & n366;
  assign n368 = n216 & n367;
  assign n369 = ~v14 & n368;
  assign n370 = v13 & n369;
  assign n371 = v11 & v8;
  assign n372 = ~v12 & n371;
  assign n373 = ~v14 & n372;
  assign n374 = v13 & n373;
  assign n375 = n147 & n374;
  assign n376 = v7 & n375;
  assign n377 = v4 & n376;
  assign n378 = ~n370 & ~n377;
  assign n379 = ~n363 & n378;
  assign n380 = ~n358 & n379;
  assign n381 = n353 & n380;
  assign n382 = n330 & n381;
  assign n383 = n305 & n382;
  assign n384 = n286 & n383;
  assign n385 = n250 & n384;
  assign n386 = n224 & n385;
  assign n387 = ~v12 & ~v9;
  assign n388 = v11 & n387;
  assign n389 = v13 & n388;
  assign n390 = v15 & n389;
  assign n391 = n147 & n390;
  assign n392 = ~v5 & n391;
  assign n393 = v7 & n392;
  assign n394 = n143 & n390;
  assign n395 = ~v5 & n394;
  assign n396 = v7 & n395;
  assign n397 = v11 & ~v7;
  assign n398 = ~v9 & n397;
  assign n399 = v15 & n398;
  assign n400 = ~v12 & n399;
  assign n401 = v13 & n400;
  assign n402 = n239 & n401;
  assign n403 = ~v3 & n402;
  assign n404 = n35 & n403;
  assign n405 = n47 & n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n396 & n406;
  assign n408 = ~n393 & n407;
  assign n409 = ~v6 & n391;
  assign n410 = v4 & n409;
  assign n411 = ~v6 & n394;
  assign n412 = v4 & n411;
  assign n413 = ~v6 & n392;
  assign n414 = ~v6 & n395;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~n412 & n415;
  assign n417 = ~n410 & n416;
  assign n418 = v11 & n104;
  assign n419 = ~v7 & n418;
  assign n420 = v8 & n419;
  assign n421 = n202 & n420;
  assign n422 = n239 & n421;
  assign n423 = v6 & n160;
  assign n424 = ~v4 & n423;
  assign n425 = v5 & n424;
  assign n426 = n420 & n425;
  assign n427 = ~v12 & v8;
  assign n428 = v11 & n427;
  assign n429 = ~v5 & ~v6;
  assign n430 = ~v2 & n429;
  assign n431 = ~v0 & n430;
  assign n432 = v1 & n431;
  assign n433 = n428 & n432;
  assign n434 = ~v14 & n433;
  assign n435 = v13 & n434;
  assign n436 = n202 & n374;
  assign n437 = v7 & n436;
  assign n438 = v4 & n437;
  assign n439 = n160 & n374;
  assign n440 = v7 & n439;
  assign n441 = v4 & n440;
  assign n442 = v13 & v15;
  assign n443 = ~v12 & n442;
  assign n444 = ~v9 & n443;
  assign n445 = v11 & n444;
  assign n446 = n147 & n445;
  assign n447 = v7 & n446;
  assign n448 = v4 & n447;
  assign n449 = n143 & n445;
  assign n450 = v7 & n449;
  assign n451 = v4 & n450;
  assign n452 = ~n448 & ~n451;
  assign n453 = ~n441 & n452;
  assign n454 = ~n438 & n453;
  assign n455 = ~n435 & n454;
  assign n456 = ~n426 & n455;
  assign n457 = ~n422 & n456;
  assign n458 = n143 & n374;
  assign n459 = ~v6 & n458;
  assign n460 = v4 & n459;
  assign n461 = n307 & n428;
  assign n462 = ~v14 & n461;
  assign n463 = v13 & n462;
  assign n464 = ~v5 & n458;
  assign n465 = ~v6 & n464;
  assign n466 = ~v5 & n436;
  assign n467 = v7 & n466;
  assign n468 = ~n465 & ~n467;
  assign n469 = ~n463 & n468;
  assign n470 = ~n460 & n469;
  assign n471 = ~v5 & n439;
  assign n472 = v7 & n471;
  assign n473 = ~v6 & n436;
  assign n474 = v4 & n473;
  assign n475 = ~v6 & n439;
  assign n476 = v4 & n475;
  assign n477 = n342 & n428;
  assign n478 = ~v14 & n477;
  assign n479 = v13 & n478;
  assign n480 = ~n476 & ~n479;
  assign n481 = ~n474 & n480;
  assign n482 = ~n472 & n481;
  assign n483 = ~v2 & n364;
  assign n484 = ~v0 & n483;
  assign n485 = v1 & n484;
  assign n486 = n216 & n485;
  assign n487 = ~v14 & n486;
  assign n488 = v13 & n487;
  assign n489 = ~v5 & n375;
  assign n490 = v7 & n489;
  assign n491 = v7 & n458;
  assign n492 = v4 & n491;
  assign n493 = ~v5 & n143;
  assign n494 = v7 & n493;
  assign n495 = n428 & n494;
  assign n496 = ~v14 & n495;
  assign n497 = v13 & n496;
  assign n498 = n239 & n420;
  assign n499 = ~v3 & n498;
  assign n500 = n35 & n499;
  assign n501 = v6 & n143;
  assign n502 = ~v4 & n501;
  assign n503 = v5 & n502;
  assign n504 = n420 & n503;
  assign n505 = v2 & n293;
  assign n506 = v0 & n505;
  assign n507 = n428 & n506;
  assign n508 = ~v14 & n507;
  assign n509 = v13 & n508;
  assign n510 = ~n504 & ~n509;
  assign n511 = ~n500 & n510;
  assign n512 = ~n497 & n511;
  assign n513 = ~n492 & n512;
  assign n514 = ~n490 & n513;
  assign n515 = ~n488 & n514;
  assign n516 = n482 & n515;
  assign n517 = n470 & n516;
  assign n518 = n457 & n517;
  assign n519 = n417 & n518;
  assign n520 = n408 & n519;
  assign n521 = ~v10 & n387;
  assign n522 = v13 & n521;
  assign n523 = v15 & n522;
  assign n524 = n202 & n523;
  assign n525 = ~v6 & n524;
  assign n526 = v4 & n525;
  assign n527 = n160 & n523;
  assign n528 = ~v6 & n527;
  assign n529 = v4 & n528;
  assign n530 = ~v5 & n524;
  assign n531 = ~v6 & n530;
  assign n532 = ~v5 & n527;
  assign n533 = ~v6 & n532;
  assign n534 = ~n531 & ~n533;
  assign n535 = ~n529 & n534;
  assign n536 = ~n526 & n535;
  assign n537 = ~v9 & n240;
  assign n538 = v15 & n537;
  assign n539 = ~v12 & n538;
  assign n540 = v13 & n539;
  assign n541 = n202 & n540;
  assign n542 = n239 & n541;
  assign n543 = n239 & n540;
  assign n544 = ~v2 & n543;
  assign n545 = n85 & n544;
  assign n546 = v7 & n524;
  assign n547 = v4 & n546;
  assign n548 = v13 & n216;
  assign n549 = v15 & n548;
  assign n550 = n147 & n549;
  assign n551 = v7 & n550;
  assign n552 = v4 & n551;
  assign n553 = ~n547 & ~n552;
  assign n554 = ~n545 & n553;
  assign n555 = ~n542 & n554;
  assign n556 = n147 & n523;
  assign n557 = ~v6 & n556;
  assign n558 = v4 & n557;
  assign n559 = n143 & n523;
  assign n560 = ~v6 & n559;
  assign n561 = v4 & n560;
  assign n562 = ~v3 & n543;
  assign n563 = n47 & n562;
  assign n564 = n307 & n521;
  assign n565 = v13 & n564;
  assign n566 = v15 & n565;
  assign n567 = n312 & n521;
  assign n568 = v13 & n567;
  assign n569 = v15 & n568;
  assign n570 = n317 & n521;
  assign n571 = v13 & n570;
  assign n572 = v15 & n571;
  assign n573 = ~v10 & n444;
  assign n574 = n160 & n573;
  assign n575 = ~v5 & n574;
  assign n576 = v7 & n575;
  assign n577 = ~n572 & ~n576;
  assign n578 = ~n569 & n577;
  assign n579 = ~n566 & n578;
  assign n580 = ~n563 & n579;
  assign n581 = ~n561 & n580;
  assign n582 = ~n558 & n581;
  assign n583 = n160 & n445;
  assign n584 = ~v5 & n583;
  assign n585 = v7 & n584;
  assign n586 = n332 & n388;
  assign n587 = v13 & n586;
  assign n588 = v15 & n587;
  assign n589 = n317 & n388;
  assign n590 = v13 & n589;
  assign n591 = v15 & n590;
  assign n592 = ~n588 & ~n591;
  assign n593 = ~n585 & n592;
  assign n594 = ~v6 & n583;
  assign n595 = v4 & n594;
  assign n596 = n342 & n388;
  assign n597 = v13 & n596;
  assign n598 = v15 & n597;
  assign n599 = n347 & n388;
  assign n600 = v13 & n599;
  assign n601 = v15 & n600;
  assign n602 = ~v7 & ~v9;
  assign n603 = n20 & n356;
  assign n604 = v11 & n603;
  assign n605 = n602 & n604;
  assign n606 = ~n601 & ~n605;
  assign n607 = ~n598 & n606;
  assign n608 = ~n595 & n607;
  assign n609 = n20 & n361;
  assign n610 = v11 & n609;
  assign n611 = n602 & n610;
  assign n612 = n202 & n445;
  assign n613 = v7 & n612;
  assign n614 = v4 & n613;
  assign n615 = v7 & n583;
  assign n616 = v4 & n615;
  assign n617 = n147 & n573;
  assign n618 = v7 & n617;
  assign n619 = v4 & n618;
  assign n620 = ~n616 & ~n619;
  assign n621 = ~n614 & n620;
  assign n622 = ~n611 & n621;
  assign n623 = n143 & n573;
  assign n624 = v7 & n623;
  assign n625 = v4 & n624;
  assign n626 = v7 & n306;
  assign n627 = n521 & n626;
  assign n628 = v13 & n627;
  assign n629 = v15 & n628;
  assign n630 = ~v5 & n623;
  assign n631 = v7 & n630;
  assign n632 = ~v4 & v5;
  assign n633 = ~v10 & n20;
  assign n634 = ~v7 & n633;
  assign n635 = ~v9 & n634;
  assign n636 = n147 & n635;
  assign n637 = v6 & n636;
  assign n638 = n632 & n637;
  assign n639 = ~n631 & ~n638;
  assign n640 = ~n629 & n639;
  assign n641 = ~n625 & n640;
  assign n642 = n622 & n641;
  assign n643 = n608 & n642;
  assign n644 = n593 & n643;
  assign n645 = n582 & n644;
  assign n646 = n555 & n645;
  assign n647 = n536 & n646;
  assign n648 = n520 & n647;
  assign n649 = n386 & n648;
  assign n650 = n199 & n649;
  assign n651 = v13 & n428;
  assign n652 = v15 & n651;
  assign n653 = n147 & n652;
  assign n654 = ~v5 & n653;
  assign n655 = v7 & n654;
  assign n656 = v13 & n495;
  assign n657 = v15 & n656;
  assign n658 = v8 & n397;
  assign n659 = n147 & n239;
  assign n660 = n658 & n659;
  assign n661 = n20 & n660;
  assign n662 = n503 & n658;
  assign n663 = n20 & n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = ~n657 & n664;
  assign n666 = ~n655 & n665;
  assign n667 = ~v6 & n653;
  assign n668 = v4 & n667;
  assign n669 = ~v6 & n143;
  assign n670 = v4 & n669;
  assign n671 = n428 & n670;
  assign n672 = v13 & n671;
  assign n673 = v15 & n672;
  assign n674 = ~v6 & n654;
  assign n675 = n143 & n652;
  assign n676 = ~v5 & n675;
  assign n677 = ~v6 & n676;
  assign n678 = ~n674 & ~n677;
  assign n679 = ~n673 & n678;
  assign n680 = ~n668 & n679;
  assign n681 = v15 & n241;
  assign n682 = ~v12 & n681;
  assign n683 = v13 & n682;
  assign n684 = n202 & n683;
  assign n685 = n239 & n684;
  assign n686 = n239 & n683;
  assign n687 = ~v2 & n686;
  assign n688 = n85 & n687;
  assign n689 = n160 & n549;
  assign n690 = ~v5 & n689;
  assign n691 = ~v6 & n690;
  assign n692 = ~v10 & n443;
  assign n693 = v8 & n692;
  assign n694 = n202 & n693;
  assign n695 = v7 & n694;
  assign n696 = v4 & n695;
  assign n697 = v13 & n372;
  assign n698 = v15 & n697;
  assign n699 = n147 & n698;
  assign n700 = v7 & n699;
  assign n701 = v4 & n700;
  assign n702 = n143 & n698;
  assign n703 = v7 & n702;
  assign n704 = v4 & n703;
  assign n705 = n160 & n693;
  assign n706 = v7 & n705;
  assign n707 = v4 & n706;
  assign n708 = ~n704 & ~n707;
  assign n709 = ~n701 & n708;
  assign n710 = ~n696 & n709;
  assign n711 = ~n691 & n710;
  assign n712 = ~n688 & n711;
  assign n713 = ~n685 & n712;
  assign n714 = v7 & n574;
  assign n715 = v4 & n714;
  assign n716 = n216 & n626;
  assign n717 = v13 & n716;
  assign n718 = v15 & n717;
  assign n719 = n143 & n693;
  assign n720 = v7 & n719;
  assign n721 = v4 & n720;
  assign n722 = ~n718 & ~n721;
  assign n723 = ~n715 & n722;
  assign n724 = ~v5 & n719;
  assign n725 = v7 & n724;
  assign n726 = v2 & n299;
  assign n727 = v0 & n726;
  assign n728 = n241 & n727;
  assign n729 = v15 & n728;
  assign n730 = n94 & n729;
  assign n731 = v15 & n302;
  assign n732 = n94 & n731;
  assign n733 = v13 & n289;
  assign n734 = v15 & n733;
  assign n735 = ~n732 & ~n734;
  assign n736 = ~n730 & n735;
  assign n737 = ~n725 & n736;
  assign n738 = ~v6 & n719;
  assign n739 = v4 & n738;
  assign n740 = v13 & n308;
  assign n741 = v15 & n740;
  assign n742 = v13 & n313;
  assign n743 = v15 & n742;
  assign n744 = v13 & n318;
  assign n745 = v15 & n744;
  assign n746 = ~n743 & ~n745;
  assign n747 = ~n741 & n746;
  assign n748 = ~n739 & n747;
  assign n749 = ~v5 & n705;
  assign n750 = v7 & n749;
  assign n751 = v13 & n333;
  assign n752 = v15 & n751;
  assign n753 = ~v6 & n705;
  assign n754 = v4 & n753;
  assign n755 = v13 & n343;
  assign n756 = v15 & n755;
  assign n757 = ~n754 & ~n756;
  assign n758 = ~n752 & n757;
  assign n759 = ~n750 & n758;
  assign n760 = n748 & n759;
  assign n761 = n737 & n760;
  assign n762 = n723 & n761;
  assign n763 = n713 & n762;
  assign n764 = n680 & n763;
  assign n765 = n666 & n764;
  assign n766 = ~v13 & ~v15;
  assign n767 = v14 & n766;
  assign n768 = n259 & n767;
  assign n769 = ~v11 & n768;
  assign n770 = n18 & n769;
  assign n771 = ~v2 & n58;
  assign n772 = ~v0 & n771;
  assign n773 = v1 & n772;
  assign n774 = n767 & n773;
  assign n775 = ~v11 & n774;
  assign n776 = n18 & n775;
  assign n777 = v3 & n70;
  assign n778 = ~v0 & n777;
  assign n779 = v1 & n778;
  assign n780 = n767 & n779;
  assign n781 = ~v11 & n780;
  assign n782 = n18 & n781;
  assign n783 = n107 & n767;
  assign n784 = ~v11 & n783;
  assign n785 = n18 & n784;
  assign n786 = ~n782 & ~n785;
  assign n787 = ~n776 & n786;
  assign n788 = ~n770 & n787;
  assign n789 = ~v15 & n40;
  assign n790 = ~v13 & n789;
  assign n791 = v14 & n790;
  assign n792 = n87 & n791;
  assign n793 = ~v7 & n792;
  assign n794 = n34 & n793;
  assign n795 = ~v13 & v14;
  assign n796 = ~v15 & n100;
  assign n797 = n795 & n796;
  assign n798 = ~v11 & n767;
  assign n799 = v9 & n798;
  assign n800 = v10 & n799;
  assign n801 = n202 & n800;
  assign n802 = ~v8 & n801;
  assign n803 = n364 & n802;
  assign n804 = v14 & ~v15;
  assign n805 = v12 & n804;
  assign n806 = v7 & n148;
  assign n807 = v4 & n806;
  assign n808 = n805 & n807;
  assign n809 = ~v11 & n808;
  assign n810 = n18 & n809;
  assign n811 = ~n803 & ~n810;
  assign n812 = ~n797 & n811;
  assign n813 = ~n794 & n812;
  assign n814 = n61 & n767;
  assign n815 = ~v11 & n814;
  assign n816 = n18 & n815;
  assign n817 = n66 & n767;
  assign n818 = ~v11 & n817;
  assign n819 = n18 & n818;
  assign n820 = ~v15 & n183;
  assign n821 = n795 & n820;
  assign n822 = ~v15 & n112;
  assign n823 = ~v13 & n822;
  assign n824 = v14 & n823;
  assign n825 = n150 & n824;
  assign n826 = n143 & n824;
  assign n827 = n70 & n826;
  assign n828 = n22 & n824;
  assign n829 = v3 & n828;
  assign n830 = n85 & n829;
  assign n831 = n160 & n824;
  assign n832 = n22 & n831;
  assign n833 = ~n830 & ~n832;
  assign n834 = ~n827 & n833;
  assign n835 = ~n825 & n834;
  assign n836 = ~n821 & n835;
  assign n837 = ~n819 & n836;
  assign n838 = ~n816 & n837;
  assign n839 = n160 & n698;
  assign n840 = ~v5 & n839;
  assign n841 = v7 & n840;
  assign n842 = n332 & n428;
  assign n843 = v13 & n842;
  assign n844 = v15 & n843;
  assign n845 = n317 & n428;
  assign n846 = v13 & n845;
  assign n847 = v15 & n846;
  assign n848 = ~n844 & ~n847;
  assign n849 = ~n841 & n848;
  assign n850 = ~v6 & n839;
  assign n851 = v4 & n850;
  assign n852 = v13 & n477;
  assign n853 = v15 & n852;
  assign n854 = n347 & n428;
  assign n855 = v13 & n854;
  assign n856 = v15 & n855;
  assign n857 = v15 & n658;
  assign n858 = ~v12 & n857;
  assign n859 = v13 & n858;
  assign n860 = n356 & n859;
  assign n861 = ~n856 & ~n860;
  assign n862 = ~n853 & n861;
  assign n863 = ~n851 & n862;
  assign n864 = n361 & n859;
  assign n865 = n202 & n698;
  assign n866 = v7 & n865;
  assign n867 = v4 & n866;
  assign n868 = v7 & n839;
  assign n869 = v4 & n868;
  assign n870 = n127 & n824;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n867 & n871;
  assign n873 = ~n864 & n872;
  assign n874 = n130 & n824;
  assign n875 = n174 & n824;
  assign n876 = n22 & n826;
  assign n877 = v6 & ~v7;
  assign n878 = v5 & n877;
  assign n879 = n37 & n791;
  assign n880 = n878 & n879;
  assign n881 = ~n876 & ~n880;
  assign n882 = ~n875 & n881;
  assign n883 = ~n874 & n882;
  assign n884 = n873 & n883;
  assign n885 = n863 & n884;
  assign n886 = n849 & n885;
  assign n887 = n838 & n886;
  assign n888 = n813 & n887;
  assign n889 = n788 & n888;
  assign n890 = n66 & n805;
  assign n891 = ~v11 & n890;
  assign n892 = n18 & n891;
  assign n893 = n73 & n805;
  assign n894 = ~v11 & n893;
  assign n895 = n18 & n894;
  assign n896 = n78 & n805;
  assign n897 = ~v11 & n896;
  assign n898 = n18 & n897;
  assign n899 = n265 & n805;
  assign n900 = ~v11 & n899;
  assign n901 = n18 & n900;
  assign n902 = ~n898 & ~n901;
  assign n903 = ~n895 & n902;
  assign n904 = ~n892 & n903;
  assign n905 = n253 & n805;
  assign n906 = ~v11 & n905;
  assign n907 = n18 & n906;
  assign n908 = n259 & n805;
  assign n909 = ~v11 & n908;
  assign n910 = n18 & n909;
  assign n911 = n773 & n805;
  assign n912 = ~v11 & n911;
  assign n913 = n18 & n912;
  assign n914 = n779 & n805;
  assign n915 = ~v11 & n914;
  assign n916 = n18 & n915;
  assign n917 = ~n913 & ~n916;
  assign n918 = ~n910 & n917;
  assign n919 = ~n907 & n918;
  assign n920 = n211 & n767;
  assign n921 = ~v11 & n920;
  assign n922 = n18 & n921;
  assign n923 = n25 & n805;
  assign n924 = ~v11 & n923;
  assign n925 = n18 & n924;
  assign n926 = ~v8 & n143;
  assign n927 = v7 & n926;
  assign n928 = v4 & n927;
  assign n929 = n805 & n928;
  assign n930 = ~v11 & n929;
  assign n931 = n18 & n930;
  assign n932 = v14 & n822;
  assign n933 = v12 & n932;
  assign n934 = n143 & n933;
  assign n935 = n22 & n934;
  assign n936 = v14 & n789;
  assign n937 = v12 & n936;
  assign n938 = n37 & n937;
  assign n939 = n878 & n938;
  assign n940 = n49 & n937;
  assign n941 = n878 & n940;
  assign n942 = ~v6 & n148;
  assign n943 = v4 & n942;
  assign n944 = n933 & n943;
  assign n945 = ~n941 & ~n944;
  assign n946 = ~n939 & n945;
  assign n947 = ~n935 & n946;
  assign n948 = ~n931 & n947;
  assign n949 = ~n925 & n948;
  assign n950 = ~n922 & n949;
  assign n951 = n388 & n626;
  assign n952 = ~v14 & n951;
  assign n953 = v13 & n952;
  assign n954 = ~v3 & n321;
  assign n955 = ~v1 & n954;
  assign n956 = v2 & n955;
  assign n957 = n388 & n956;
  assign n958 = ~v14 & n957;
  assign n959 = v13 & n958;
  assign n960 = n104 & n727;
  assign n961 = v11 & n960;
  assign n962 = n602 & n961;
  assign n963 = n104 & n301;
  assign n964 = v11 & n963;
  assign n965 = n602 & n964;
  assign n966 = ~n962 & ~n965;
  assign n967 = ~n959 & n966;
  assign n968 = ~n953 & n967;
  assign n969 = n288 & n388;
  assign n970 = ~v14 & n969;
  assign n971 = v13 & n970;
  assign n972 = n295 & n388;
  assign n973 = ~v14 & n972;
  assign n974 = v13 & n973;
  assign n975 = n307 & n388;
  assign n976 = ~v14 & n975;
  assign n977 = v13 & n976;
  assign n978 = n312 & n388;
  assign n979 = ~v14 & n978;
  assign n980 = v13 & n979;
  assign n981 = ~n977 & ~n980;
  assign n982 = ~n974 & n981;
  assign n983 = ~n971 & n982;
  assign n984 = n87 & n937;
  assign n985 = n878 & n984;
  assign n986 = n96 & n937;
  assign n987 = n878 & n986;
  assign n988 = n160 & n933;
  assign n989 = n70 & n988;
  assign n990 = n205 & n805;
  assign n991 = ~v11 & n990;
  assign n992 = n18 & n991;
  assign n993 = n211 & n805;
  assign n994 = ~v11 & n993;
  assign n995 = n18 & n994;
  assign n996 = n218 & n388;
  assign n997 = ~v14 & n996;
  assign n998 = v13 & n997;
  assign n999 = n226 & n388;
  assign n1000 = ~v14 & n999;
  assign n1001 = v13 & n1000;
  assign n1002 = ~n998 & ~n1001;
  assign n1003 = ~n995 & n1002;
  assign n1004 = ~n992 & n1003;
  assign n1005 = ~n989 & n1004;
  assign n1006 = ~n987 & n1005;
  assign n1007 = ~n985 & n1006;
  assign n1008 = n983 & n1007;
  assign n1009 = n968 & n1008;
  assign n1010 = n950 & n1009;
  assign n1011 = n919 & n1010;
  assign n1012 = n904 & n1011;
  assign n1013 = ~v14 & n398;
  assign n1014 = ~v12 & n1013;
  assign n1015 = v13 & n1014;
  assign n1016 = n239 & n1015;
  assign n1017 = ~v2 & n1016;
  assign n1018 = n85 & n1017;
  assign n1019 = v3 & n85;
  assign n1020 = v7 & n1019;
  assign n1021 = v4 & n1020;
  assign n1022 = n388 & n1021;
  assign n1023 = ~v14 & n1022;
  assign n1024 = v13 & n1023;
  assign n1025 = ~v13 & ~v9;
  assign n1026 = v11 & n1025;
  assign n1027 = n218 & n1026;
  assign n1028 = ~v15 & n1027;
  assign n1029 = v14 & n1028;
  assign n1030 = n226 & n1026;
  assign n1031 = ~v15 & n1030;
  assign n1032 = v14 & n1031;
  assign n1033 = ~n1029 & ~n1032;
  assign n1034 = ~n1024 & n1033;
  assign n1035 = ~n1018 & n1034;
  assign n1036 = v7 & n160;
  assign n1037 = v4 & n1036;
  assign n1038 = n388 & n1037;
  assign n1039 = ~v14 & n1038;
  assign n1040 = v13 & n1039;
  assign n1041 = ~v15 & n1026;
  assign n1042 = v14 & n1041;
  assign n1043 = n147 & n1042;
  assign n1044 = ~v5 & n1043;
  assign n1045 = v7 & n1044;
  assign n1046 = n143 & n1042;
  assign n1047 = ~v5 & n1046;
  assign n1048 = v7 & n1047;
  assign n1049 = ~v15 & n398;
  assign n1050 = ~v13 & n1049;
  assign n1051 = v14 & n1050;
  assign n1052 = n239 & n1051;
  assign n1053 = ~v3 & n1052;
  assign n1054 = n35 & n1053;
  assign n1055 = ~n1048 & ~n1054;
  assign n1056 = ~n1045 & n1055;
  assign n1057 = ~n1040 & n1056;
  assign n1058 = ~v14 & n388;
  assign n1059 = v13 & n1058;
  assign n1060 = n160 & n1059;
  assign n1061 = ~v5 & n1060;
  assign n1062 = v7 & n1061;
  assign n1063 = n202 & n1059;
  assign n1064 = ~v6 & n1063;
  assign n1065 = v4 & n1064;
  assign n1066 = ~v5 & n1063;
  assign n1067 = v7 & n1066;
  assign n1068 = n338 & n388;
  assign n1069 = ~v14 & n1068;
  assign n1070 = v13 & n1069;
  assign n1071 = ~v14 & n596;
  assign n1072 = v13 & n1071;
  assign n1073 = ~v14 & n599;
  assign n1074 = v13 & n1073;
  assign n1075 = n104 & n356;
  assign n1076 = v11 & n1075;
  assign n1077 = n602 & n1076;
  assign n1078 = ~n1074 & ~n1077;
  assign n1079 = ~n1072 & n1078;
  assign n1080 = ~n1070 & n1079;
  assign n1081 = ~n1067 & n1080;
  assign n1082 = ~n1065 & n1081;
  assign n1083 = ~n1062 & n1082;
  assign n1084 = n288 & n1026;
  assign n1085 = ~v15 & n1084;
  assign n1086 = v14 & n1085;
  assign n1087 = n295 & n1026;
  assign n1088 = ~v15 & n1087;
  assign n1089 = v14 & n1088;
  assign n1090 = n301 & n767;
  assign n1091 = v11 & n1090;
  assign n1092 = n602 & n1091;
  assign n1093 = ~n1089 & ~n1092;
  assign n1094 = ~n1086 & n1093;
  assign n1095 = n307 & n1026;
  assign n1096 = ~v15 & n1095;
  assign n1097 = v14 & n1096;
  assign n1098 = n312 & n1026;
  assign n1099 = ~v15 & n1098;
  assign n1100 = v14 & n1099;
  assign n1101 = n317 & n1026;
  assign n1102 = ~v15 & n1101;
  assign n1103 = v14 & n1102;
  assign n1104 = n324 & n1026;
  assign n1105 = ~v15 & n1104;
  assign n1106 = v14 & n1105;
  assign n1107 = ~n1103 & ~n1106;
  assign n1108 = ~n1100 & n1107;
  assign n1109 = ~n1097 & n1108;
  assign n1110 = n332 & n1026;
  assign n1111 = ~v15 & n1110;
  assign n1112 = v14 & n1111;
  assign n1113 = n338 & n1026;
  assign n1114 = ~v15 & n1113;
  assign n1115 = v14 & n1114;
  assign n1116 = n342 & n1026;
  assign n1117 = ~v15 & n1116;
  assign n1118 = v14 & n1117;
  assign n1119 = n347 & n1026;
  assign n1120 = ~v15 & n1119;
  assign n1121 = v14 & n1120;
  assign n1122 = ~n1118 & ~n1121;
  assign n1123 = ~n1115 & n1122;
  assign n1124 = ~n1112 & n1123;
  assign n1125 = n356 & n767;
  assign n1126 = v11 & n1125;
  assign n1127 = n602 & n1126;
  assign n1128 = n361 & n767;
  assign n1129 = v11 & n1128;
  assign n1130 = n602 & n1129;
  assign n1131 = n367 & n1026;
  assign n1132 = ~v15 & n1131;
  assign n1133 = v14 & n1132;
  assign n1134 = n485 & n1026;
  assign n1135 = ~v15 & n1134;
  assign n1136 = v14 & n1135;
  assign n1137 = ~n1133 & ~n1136;
  assign n1138 = ~n1130 & n1137;
  assign n1139 = ~n1127 & n1138;
  assign n1140 = n1124 & n1139;
  assign n1141 = n1109 & n1140;
  assign n1142 = n1094 & n1141;
  assign n1143 = n1083 & n1142;
  assign n1144 = n1057 & n1143;
  assign n1145 = n1035 & n1144;
  assign n1146 = n1012 & n1145;
  assign n1147 = n889 & n1146;
  assign n1148 = n765 & n1147;
  assign n1149 = ~v13 & v8;
  assign n1150 = v11 & n1149;
  assign n1151 = v2 & n954;
  assign n1152 = v0 & n1151;
  assign n1153 = n1150 & n1152;
  assign n1154 = ~v15 & n1153;
  assign n1155 = v14 & n1154;
  assign n1156 = n494 & n1150;
  assign n1157 = ~v15 & n1156;
  assign n1158 = v14 & n1157;
  assign n1159 = v11 & n767;
  assign n1160 = ~v7 & n1159;
  assign n1161 = v8 & n1160;
  assign n1162 = n239 & n1161;
  assign n1163 = ~v3 & n1162;
  assign n1164 = n35 & n1163;
  assign n1165 = n503 & n1161;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = ~n1158 & n1166;
  assign n1168 = ~n1155 & n1167;
  assign n1169 = n506 & n1150;
  assign n1170 = ~v15 & n1169;
  assign n1171 = v14 & n1170;
  assign n1172 = n670 & n1150;
  assign n1173 = ~v15 & n1172;
  assign n1174 = v14 & n1173;
  assign n1175 = ~v3 & n429;
  assign n1176 = v2 & n1175;
  assign n1177 = v0 & n1176;
  assign n1178 = n1150 & n1177;
  assign n1179 = ~v15 & n1178;
  assign n1180 = v14 & n1179;
  assign n1181 = ~v1 & n1175;
  assign n1182 = v2 & n1181;
  assign n1183 = n1150 & n1182;
  assign n1184 = ~v15 & n1183;
  assign n1185 = v14 & n1184;
  assign n1186 = ~n1180 & ~n1185;
  assign n1187 = ~n1174 & n1186;
  assign n1188 = ~n1171 & n1187;
  assign n1189 = ~v15 & n241;
  assign n1190 = ~v13 & n1189;
  assign n1191 = v14 & n1190;
  assign n1192 = n202 & n1191;
  assign n1193 = n239 & n1192;
  assign n1194 = n239 & n1191;
  assign n1195 = ~v2 & n1194;
  assign n1196 = n85 & n1195;
  assign n1197 = ~v10 & ~v13;
  assign n1198 = v8 & n1197;
  assign n1199 = ~v15 & n1198;
  assign n1200 = v14 & n1199;
  assign n1201 = n160 & n1200;
  assign n1202 = ~v5 & n1201;
  assign n1203 = ~v6 & n1202;
  assign n1204 = n367 & n1198;
  assign n1205 = ~v15 & n1204;
  assign n1206 = v14 & n1205;
  assign n1207 = ~v13 & n371;
  assign n1208 = ~v15 & n1207;
  assign n1209 = v14 & n1208;
  assign n1210 = n147 & n1209;
  assign n1211 = v7 & n1210;
  assign n1212 = v4 & n1211;
  assign n1213 = n143 & n1209;
  assign n1214 = v7 & n1213;
  assign n1215 = v4 & n1214;
  assign n1216 = n485 & n1198;
  assign n1217 = ~v15 & n1216;
  assign n1218 = v14 & n1217;
  assign n1219 = ~n1215 & ~n1218;
  assign n1220 = ~n1212 & n1219;
  assign n1221 = ~n1206 & n1220;
  assign n1222 = ~n1203 & n1221;
  assign n1223 = ~n1196 & n1222;
  assign n1224 = ~n1193 & n1223;
  assign n1225 = ~v3 & n364;
  assign n1226 = ~v1 & n1225;
  assign n1227 = v2 & n1226;
  assign n1228 = n1198 & n1227;
  assign n1229 = ~v15 & n1228;
  assign n1230 = v14 & n1229;
  assign n1231 = n626 & n1198;
  assign n1232 = ~v15 & n1231;
  assign n1233 = v14 & n1232;
  assign n1234 = v2 & n1225;
  assign n1235 = v0 & n1234;
  assign n1236 = n1198 & n1235;
  assign n1237 = ~v15 & n1236;
  assign n1238 = v14 & n1237;
  assign n1239 = ~n1233 & ~n1238;
  assign n1240 = ~n1230 & n1239;
  assign n1241 = n956 & n1198;
  assign n1242 = ~v15 & n1241;
  assign n1243 = v14 & n1242;
  assign n1244 = n728 & n767;
  assign n1245 = n302 & n767;
  assign n1246 = n288 & n1198;
  assign n1247 = ~v15 & n1246;
  assign n1248 = v14 & n1247;
  assign n1249 = ~n1245 & ~n1248;
  assign n1250 = ~n1244 & n1249;
  assign n1251 = ~n1243 & n1250;
  assign n1252 = n295 & n1198;
  assign n1253 = ~v15 & n1252;
  assign n1254 = v14 & n1253;
  assign n1255 = n307 & n1198;
  assign n1256 = ~v15 & n1255;
  assign n1257 = v14 & n1256;
  assign n1258 = n312 & n1198;
  assign n1259 = ~v15 & n1258;
  assign n1260 = v14 & n1259;
  assign n1261 = n317 & n1198;
  assign n1262 = ~v15 & n1261;
  assign n1263 = v14 & n1262;
  assign n1264 = ~n1260 & ~n1263;
  assign n1265 = ~n1257 & n1264;
  assign n1266 = ~n1254 & n1265;
  assign n1267 = n324 & n1198;
  assign n1268 = ~v15 & n1267;
  assign n1269 = v14 & n1268;
  assign n1270 = n332 & n1198;
  assign n1271 = ~v15 & n1270;
  assign n1272 = v14 & n1271;
  assign n1273 = n338 & n1198;
  assign n1274 = ~v15 & n1273;
  assign n1275 = v14 & n1274;
  assign n1276 = n342 & n1198;
  assign n1277 = ~v15 & n1276;
  assign n1278 = v14 & n1277;
  assign n1279 = ~n1275 & ~n1278;
  assign n1280 = ~n1272 & n1279;
  assign n1281 = ~n1269 & n1280;
  assign n1282 = n1266 & n1281;
  assign n1283 = n1251 & n1282;
  assign n1284 = n1240 & n1283;
  assign n1285 = n1224 & n1284;
  assign n1286 = n1188 & n1285;
  assign n1287 = n1168 & n1286;
  assign n1288 = v12 & ~v9;
  assign n1289 = v11 & n1288;
  assign n1290 = v3 & n292;
  assign n1291 = ~v0 & n1290;
  assign n1292 = v1 & n1291;
  assign n1293 = n1289 & n1292;
  assign n1294 = ~v15 & n1293;
  assign n1295 = v14 & n1294;
  assign n1296 = ~v6 & n160;
  assign n1297 = v4 & n1296;
  assign n1298 = n1289 & n1297;
  assign n1299 = ~v15 & n1298;
  assign n1300 = v14 & n1299;
  assign n1301 = v3 & n429;
  assign n1302 = ~v0 & n1301;
  assign n1303 = v1 & n1302;
  assign n1304 = n1289 & n1303;
  assign n1305 = ~v15 & n1304;
  assign n1306 = v14 & n1305;
  assign n1307 = n432 & n1289;
  assign n1308 = ~v15 & n1307;
  assign n1309 = v14 & n1308;
  assign n1310 = ~n1306 & ~n1309;
  assign n1311 = ~n1300 & n1310;
  assign n1312 = ~n1295 & n1311;
  assign n1313 = v14 & n1049;
  assign n1314 = v12 & n1313;
  assign n1315 = n202 & n1314;
  assign n1316 = n239 & n1315;
  assign n1317 = n239 & n1314;
  assign n1318 = ~v2 & n1317;
  assign n1319 = n85 & n1318;
  assign n1320 = n1021 & n1289;
  assign n1321 = ~v15 & n1320;
  assign n1322 = v14 & n1321;
  assign n1323 = n1037 & n1289;
  assign n1324 = ~v15 & n1323;
  assign n1325 = v14 & n1324;
  assign n1326 = ~n1322 & ~n1325;
  assign n1327 = ~n1319 & n1326;
  assign n1328 = ~n1316 & n1327;
  assign n1329 = n506 & n1289;
  assign n1330 = ~v15 & n1329;
  assign n1331 = v14 & n1330;
  assign n1332 = n670 & n1289;
  assign n1333 = ~v15 & n1332;
  assign n1334 = v14 & n1333;
  assign n1335 = ~v3 & n1317;
  assign n1336 = n47 & n1335;
  assign n1337 = n307 & n1289;
  assign n1338 = ~v15 & n1337;
  assign n1339 = v14 & n1338;
  assign n1340 = n312 & n1289;
  assign n1341 = ~v15 & n1340;
  assign n1342 = v14 & n1341;
  assign n1343 = ~v15 & n1289;
  assign n1344 = v14 & n1343;
  assign n1345 = n202 & n1344;
  assign n1346 = ~v5 & n1345;
  assign n1347 = v7 & n1346;
  assign n1348 = n160 & n1344;
  assign n1349 = ~v5 & n1348;
  assign n1350 = v7 & n1349;
  assign n1351 = ~n1347 & ~n1350;
  assign n1352 = ~n1342 & n1351;
  assign n1353 = ~n1339 & n1352;
  assign n1354 = ~n1336 & n1353;
  assign n1355 = ~n1334 & n1354;
  assign n1356 = ~n1331 & n1355;
  assign n1357 = ~v15 & n658;
  assign n1358 = ~v13 & n1357;
  assign n1359 = v14 & n1358;
  assign n1360 = n361 & n1359;
  assign n1361 = n202 & n1209;
  assign n1362 = v7 & n1361;
  assign n1363 = v4 & n1362;
  assign n1364 = n160 & n1209;
  assign n1365 = v7 & n1364;
  assign n1366 = v4 & n1365;
  assign n1367 = n147 & n1344;
  assign n1368 = v7 & n1367;
  assign n1369 = v4 & n1368;
  assign n1370 = ~n1366 & ~n1369;
  assign n1371 = ~n1363 & n1370;
  assign n1372 = ~n1360 & n1371;
  assign n1373 = n143 & n1344;
  assign n1374 = v7 & n1373;
  assign n1375 = v4 & n1374;
  assign n1376 = n626 & n1289;
  assign n1377 = ~v15 & n1376;
  assign n1378 = v14 & n1377;
  assign n1379 = ~v5 & n1373;
  assign n1380 = v7 & n1379;
  assign n1381 = n727 & n805;
  assign n1382 = v11 & n1381;
  assign n1383 = n602 & n1382;
  assign n1384 = ~n1380 & ~n1383;
  assign n1385 = ~n1378 & n1384;
  assign n1386 = ~n1375 & n1385;
  assign n1387 = ~v5 & n1364;
  assign n1388 = v7 & n1387;
  assign n1389 = ~v6 & n1361;
  assign n1390 = v4 & n1389;
  assign n1391 = ~v5 & n1361;
  assign n1392 = v7 & n1391;
  assign n1393 = n1150 & n1297;
  assign n1394 = ~v15 & n1393;
  assign n1395 = v14 & n1394;
  assign n1396 = n1150 & n1303;
  assign n1397 = ~v15 & n1396;
  assign n1398 = v14 & n1397;
  assign n1399 = n432 & n1150;
  assign n1400 = ~v15 & n1399;
  assign n1401 = v14 & n1400;
  assign n1402 = n202 & n1161;
  assign n1403 = n239 & n1402;
  assign n1404 = ~n1401 & ~n1403;
  assign n1405 = ~n1398 & n1404;
  assign n1406 = ~n1395 & n1405;
  assign n1407 = ~n1392 & n1406;
  assign n1408 = ~n1390 & n1407;
  assign n1409 = ~n1388 & n1408;
  assign n1410 = n1386 & n1409;
  assign n1411 = n1372 & n1410;
  assign n1412 = n1356 & n1411;
  assign n1413 = n1328 & n1412;
  assign n1414 = n1312 & n1413;
  assign n1415 = ~v10 & n1025;
  assign n1416 = ~v15 & n1415;
  assign n1417 = v14 & n1416;
  assign n1418 = n147 & n1417;
  assign n1419 = ~v5 & n1418;
  assign n1420 = v7 & n1419;
  assign n1421 = n143 & n1417;
  assign n1422 = ~v5 & n1421;
  assign n1423 = v7 & n1422;
  assign n1424 = ~v15 & n537;
  assign n1425 = ~v13 & n1424;
  assign n1426 = v14 & n1425;
  assign n1427 = n239 & n1426;
  assign n1428 = ~v3 & n1427;
  assign n1429 = n35 & n1428;
  assign n1430 = n47 & n1428;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1423 & n1431;
  assign n1433 = ~n1420 & n1432;
  assign n1434 = ~v6 & n1418;
  assign n1435 = v4 & n1434;
  assign n1436 = ~v6 & n1421;
  assign n1437 = v4 & n1436;
  assign n1438 = ~v6 & n1419;
  assign n1439 = ~v6 & n1422;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1437 & n1440;
  assign n1442 = ~n1435 & n1441;
  assign n1443 = ~v14 & n537;
  assign n1444 = ~v12 & n1443;
  assign n1445 = v13 & n1444;
  assign n1446 = n202 & n1445;
  assign n1447 = n239 & n1446;
  assign n1448 = n239 & n1445;
  assign n1449 = ~v2 & n1448;
  assign n1450 = n85 & n1449;
  assign n1451 = ~v14 & n521;
  assign n1452 = v13 & n1451;
  assign n1453 = n160 & n1452;
  assign n1454 = ~v5 & n1453;
  assign n1455 = ~v6 & n1454;
  assign n1456 = n367 & n521;
  assign n1457 = ~v14 & n1456;
  assign n1458 = v13 & n1457;
  assign n1459 = n1235 & n1415;
  assign n1460 = ~v15 & n1459;
  assign n1461 = v14 & n1460;
  assign n1462 = n1227 & n1415;
  assign n1463 = ~v15 & n1462;
  assign n1464 = v14 & n1463;
  assign n1465 = n485 & n521;
  assign n1466 = ~v14 & n1465;
  assign n1467 = v13 & n1466;
  assign n1468 = ~n1464 & ~n1467;
  assign n1469 = ~n1461 & n1468;
  assign n1470 = ~n1458 & n1469;
  assign n1471 = ~n1455 & n1470;
  assign n1472 = ~n1450 & n1471;
  assign n1473 = ~n1447 & n1472;
  assign n1474 = n521 & n1227;
  assign n1475 = ~v14 & n1474;
  assign n1476 = v13 & n1475;
  assign n1477 = ~v14 & n627;
  assign n1478 = v13 & n1477;
  assign n1479 = n521 & n1235;
  assign n1480 = ~v14 & n1479;
  assign n1481 = v13 & n1480;
  assign n1482 = ~n1478 & ~n1481;
  assign n1483 = ~n1476 & n1482;
  assign n1484 = n521 & n956;
  assign n1485 = ~v14 & n1484;
  assign n1486 = v13 & n1485;
  assign n1487 = n537 & n727;
  assign n1488 = n104 & n1487;
  assign n1489 = n301 & n537;
  assign n1490 = n104 & n1489;
  assign n1491 = n288 & n521;
  assign n1492 = ~v14 & n1491;
  assign n1493 = v13 & n1492;
  assign n1494 = ~n1490 & ~n1493;
  assign n1495 = ~n1488 & n1494;
  assign n1496 = ~n1486 & n1495;
  assign n1497 = n295 & n521;
  assign n1498 = ~v14 & n1497;
  assign n1499 = v13 & n1498;
  assign n1500 = ~v14 & n564;
  assign n1501 = v13 & n1500;
  assign n1502 = ~v14 & n567;
  assign n1503 = v13 & n1502;
  assign n1504 = ~v14 & n570;
  assign n1505 = v13 & n1504;
  assign n1506 = ~n1503 & ~n1505;
  assign n1507 = ~n1501 & n1506;
  assign n1508 = ~n1499 & n1507;
  assign n1509 = n324 & n521;
  assign n1510 = ~v14 & n1509;
  assign n1511 = v13 & n1510;
  assign n1512 = n332 & n521;
  assign n1513 = ~v14 & n1512;
  assign n1514 = v13 & n1513;
  assign n1515 = n338 & n521;
  assign n1516 = ~v14 & n1515;
  assign n1517 = v13 & n1516;
  assign n1518 = n342 & n521;
  assign n1519 = ~v14 & n1518;
  assign n1520 = v13 & n1519;
  assign n1521 = ~n1517 & ~n1520;
  assign n1522 = ~n1514 & n1521;
  assign n1523 = ~n1511 & n1522;
  assign n1524 = n1508 & n1523;
  assign n1525 = n1496 & n1524;
  assign n1526 = n1483 & n1525;
  assign n1527 = n1473 & n1526;
  assign n1528 = n1442 & n1527;
  assign n1529 = n1433 & n1528;
  assign n1530 = ~v10 & ~v9;
  assign n1531 = v12 & n1530;
  assign n1532 = ~v15 & n1531;
  assign n1533 = v14 & n1532;
  assign n1534 = n202 & n1533;
  assign n1535 = ~v6 & n1534;
  assign n1536 = v4 & n1535;
  assign n1537 = n160 & n1533;
  assign n1538 = ~v6 & n1537;
  assign n1539 = v4 & n1538;
  assign n1540 = ~v5 & n1534;
  assign n1541 = ~v6 & n1540;
  assign n1542 = ~v5 & n1537;
  assign n1543 = ~v6 & n1542;
  assign n1544 = ~n1541 & ~n1543;
  assign n1545 = ~n1539 & n1544;
  assign n1546 = ~n1536 & n1545;
  assign n1547 = v14 & n1424;
  assign n1548 = v12 & n1547;
  assign n1549 = n202 & n1548;
  assign n1550 = n239 & n1549;
  assign n1551 = n239 & n1548;
  assign n1552 = ~v2 & n1551;
  assign n1553 = n85 & n1552;
  assign n1554 = v7 & n1534;
  assign n1555 = v4 & n1554;
  assign n1556 = ~v10 & v12;
  assign n1557 = v8 & n1556;
  assign n1558 = n218 & n1557;
  assign n1559 = ~v15 & n1558;
  assign n1560 = v14 & n1559;
  assign n1561 = ~n1555 & ~n1560;
  assign n1562 = ~n1553 & n1561;
  assign n1563 = ~n1550 & n1562;
  assign n1564 = n147 & n1533;
  assign n1565 = ~v6 & n1564;
  assign n1566 = v4 & n1565;
  assign n1567 = n143 & n1533;
  assign n1568 = ~v6 & n1567;
  assign n1569 = v4 & n1568;
  assign n1570 = ~v3 & n1551;
  assign n1571 = n47 & n1570;
  assign n1572 = ~v10 & n1288;
  assign n1573 = n307 & n1572;
  assign n1574 = ~v15 & n1573;
  assign n1575 = v14 & n1574;
  assign n1576 = n312 & n1572;
  assign n1577 = ~v15 & n1576;
  assign n1578 = v14 & n1577;
  assign n1579 = n317 & n1572;
  assign n1580 = ~v15 & n1579;
  assign n1581 = v14 & n1580;
  assign n1582 = n324 & n1572;
  assign n1583 = ~v15 & n1582;
  assign n1584 = v14 & n1583;
  assign n1585 = ~n1581 & ~n1584;
  assign n1586 = ~n1578 & n1585;
  assign n1587 = ~n1575 & n1586;
  assign n1588 = ~n1571 & n1587;
  assign n1589 = ~n1569 & n1588;
  assign n1590 = ~n1566 & n1589;
  assign n1591 = n324 & n1415;
  assign n1592 = ~v15 & n1591;
  assign n1593 = v14 & n1592;
  assign n1594 = n332 & n1415;
  assign n1595 = ~v15 & n1594;
  assign n1596 = v14 & n1595;
  assign n1597 = n317 & n1415;
  assign n1598 = ~v15 & n1597;
  assign n1599 = v14 & n1598;
  assign n1600 = ~n1596 & ~n1599;
  assign n1601 = ~n1593 & n1600;
  assign n1602 = n338 & n1415;
  assign n1603 = ~v15 & n1602;
  assign n1604 = v14 & n1603;
  assign n1605 = n342 & n1415;
  assign n1606 = ~v15 & n1605;
  assign n1607 = v14 & n1606;
  assign n1608 = n347 & n1415;
  assign n1609 = ~v15 & n1608;
  assign n1610 = v14 & n1609;
  assign n1611 = n356 & n537;
  assign n1612 = n767 & n1611;
  assign n1613 = ~n1610 & ~n1612;
  assign n1614 = ~n1607 & n1613;
  assign n1615 = ~n1604 & n1614;
  assign n1616 = n361 & n537;
  assign n1617 = n767 & n1616;
  assign n1618 = n367 & n1415;
  assign n1619 = ~v15 & n1618;
  assign n1620 = v14 & n1619;
  assign n1621 = n1235 & n1572;
  assign n1622 = ~v15 & n1621;
  assign n1623 = v14 & n1622;
  assign n1624 = n1227 & n1572;
  assign n1625 = ~v15 & n1624;
  assign n1626 = v14 & n1625;
  assign n1627 = ~n1623 & ~n1626;
  assign n1628 = ~n1620 & n1627;
  assign n1629 = ~n1617 & n1628;
  assign n1630 = n485 & n1415;
  assign n1631 = ~v15 & n1630;
  assign n1632 = v14 & n1631;
  assign n1633 = n626 & n1572;
  assign n1634 = ~v15 & n1633;
  assign n1635 = v14 & n1634;
  assign n1636 = n956 & n1572;
  assign n1637 = ~v15 & n1636;
  assign n1638 = v14 & n1637;
  assign n1639 = ~v10 & n805;
  assign n1640 = ~v7 & n1639;
  assign n1641 = ~v9 & n1640;
  assign n1642 = n147 & n1641;
  assign n1643 = v6 & n1642;
  assign n1644 = n632 & n1643;
  assign n1645 = ~n1638 & ~n1644;
  assign n1646 = ~n1635 & n1645;
  assign n1647 = ~n1632 & n1646;
  assign n1648 = n1629 & n1647;
  assign n1649 = n1615 & n1648;
  assign n1650 = n1601 & n1649;
  assign n1651 = n1590 & n1650;
  assign n1652 = n1563 & n1651;
  assign n1653 = n1546 & n1652;
  assign n1654 = n1529 & n1653;
  assign n1655 = n1414 & n1654;
  assign n1656 = n1287 & n1655;
  assign n1657 = v12 & v8;
  assign n1658 = v11 & n1657;
  assign n1659 = n1152 & n1658;
  assign n1660 = ~v15 & n1659;
  assign n1661 = v14 & n1660;
  assign n1662 = n494 & n1658;
  assign n1663 = ~v15 & n1662;
  assign n1664 = v14 & n1663;
  assign n1665 = n660 & n805;
  assign n1666 = v12 & v14;
  assign n1667 = ~v15 & n662;
  assign n1668 = n1666 & n1667;
  assign n1669 = ~n1665 & ~n1668;
  assign n1670 = ~n1664 & n1669;
  assign n1671 = ~n1661 & n1670;
  assign n1672 = n506 & n1658;
  assign n1673 = ~v15 & n1672;
  assign n1674 = v14 & n1673;
  assign n1675 = n670 & n1658;
  assign n1676 = ~v15 & n1675;
  assign n1677 = v14 & n1676;
  assign n1678 = n1177 & n1658;
  assign n1679 = ~v15 & n1678;
  assign n1680 = v14 & n1679;
  assign n1681 = n1182 & n1658;
  assign n1682 = ~v15 & n1681;
  assign n1683 = v14 & n1682;
  assign n1684 = ~n1680 & ~n1683;
  assign n1685 = ~n1677 & n1684;
  assign n1686 = ~n1674 & n1685;
  assign n1687 = v14 & n1189;
  assign n1688 = v12 & n1687;
  assign n1689 = n202 & n1688;
  assign n1690 = n239 & n1689;
  assign n1691 = n239 & n1688;
  assign n1692 = ~v2 & n1691;
  assign n1693 = n85 & n1692;
  assign n1694 = n432 & n1557;
  assign n1695 = ~v15 & n1694;
  assign n1696 = v14 & n1695;
  assign n1697 = ~v15 & n1557;
  assign n1698 = v14 & n1697;
  assign n1699 = n202 & n1698;
  assign n1700 = v7 & n1699;
  assign n1701 = v4 & n1700;
  assign n1702 = ~v15 & n1658;
  assign n1703 = v14 & n1702;
  assign n1704 = n147 & n1703;
  assign n1705 = v7 & n1704;
  assign n1706 = v4 & n1705;
  assign n1707 = n143 & n1703;
  assign n1708 = v7 & n1707;
  assign n1709 = v4 & n1708;
  assign n1710 = n160 & n1698;
  assign n1711 = v7 & n1710;
  assign n1712 = v4 & n1711;
  assign n1713 = ~n1709 & ~n1712;
  assign n1714 = ~n1706 & n1713;
  assign n1715 = ~n1701 & n1714;
  assign n1716 = ~n1696 & n1715;
  assign n1717 = ~n1693 & n1716;
  assign n1718 = ~n1690 & n1717;
  assign n1719 = n143 & n1698;
  assign n1720 = ~v6 & n1719;
  assign n1721 = v4 & n1720;
  assign n1722 = n307 & n1557;
  assign n1723 = ~v15 & n1722;
  assign n1724 = v14 & n1723;
  assign n1725 = n312 & n1557;
  assign n1726 = ~v15 & n1725;
  assign n1727 = v14 & n1726;
  assign n1728 = ~v5 & n1699;
  assign n1729 = v7 & n1728;
  assign n1730 = ~n1727 & ~n1729;
  assign n1731 = ~n1724 & n1730;
  assign n1732 = ~n1721 & n1731;
  assign n1733 = ~v5 & n1710;
  assign n1734 = v7 & n1733;
  assign n1735 = ~v6 & n1699;
  assign n1736 = v4 & n1735;
  assign n1737 = ~v6 & n1710;
  assign n1738 = v4 & n1737;
  assign n1739 = n342 & n1557;
  assign n1740 = ~v15 & n1739;
  assign n1741 = v14 & n1740;
  assign n1742 = ~n1738 & ~n1741;
  assign n1743 = ~n1736 & n1742;
  assign n1744 = ~n1734 & n1743;
  assign n1745 = n485 & n1572;
  assign n1746 = ~v15 & n1745;
  assign n1747 = v14 & n1746;
  assign n1748 = n626 & n1557;
  assign n1749 = ~v15 & n1748;
  assign n1750 = v14 & n1749;
  assign n1751 = v7 & n1719;
  assign n1752 = v4 & n1751;
  assign n1753 = n494 & n1557;
  assign n1754 = ~v15 & n1753;
  assign n1755 = v14 & n1754;
  assign n1756 = ~v3 & n1691;
  assign n1757 = n35 & n1756;
  assign n1758 = n47 & n1756;
  assign n1759 = n506 & n1557;
  assign n1760 = ~v15 & n1759;
  assign n1761 = v14 & n1760;
  assign n1762 = ~n1758 & ~n1761;
  assign n1763 = ~n1757 & n1762;
  assign n1764 = ~n1755 & n1763;
  assign n1765 = ~n1752 & n1764;
  assign n1766 = ~n1750 & n1765;
  assign n1767 = ~n1747 & n1766;
  assign n1768 = n1744 & n1767;
  assign n1769 = n1732 & n1768;
  assign n1770 = n1718 & n1769;
  assign n1771 = n1686 & n1770;
  assign n1772 = n1671 & n1771;
  assign n1773 = ~v4 & v7;
  assign n1774 = v5 & n1773;
  assign n1775 = v11 & n1774;
  assign n1776 = ~v8 & n1775;
  assign n1777 = v9 & n1776;
  assign n1778 = ~v11 & n1774;
  assign n1779 = v8 & n1778;
  assign n1780 = v10 & n1779;
  assign n1781 = ~v13 & n1774;
  assign n1782 = v15 & n1781;
  assign n1783 = ~v14 & n1781;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1780 & n1784;
  assign n1786 = ~n1777 & n1785;
  assign n1787 = ~v9 & n1778;
  assign n1788 = v10 & n1787;
  assign n1789 = ~v10 & n1774;
  assign n1790 = ~v8 & n1789;
  assign n1791 = v9 & n1790;
  assign n1792 = ~v6 & n632;
  assign n1793 = ~v14 & n1792;
  assign n1794 = v12 & n1793;
  assign n1795 = ~v12 & n1792;
  assign n1796 = ~v15 & n1795;
  assign n1797 = v13 & n1796;
  assign n1798 = v14 & n1797;
  assign n1799 = ~n1794 & ~n1798;
  assign n1800 = ~n1791 & n1799;
  assign n1801 = ~n1788 & n1800;
  assign n1802 = ~v0 & v2;
  assign n1803 = v1 & n1802;
  assign n1804 = ~v14 & n1803;
  assign n1805 = ~v3 & n1804;
  assign n1806 = ~v13 & n1805;
  assign n1807 = ~v3 & n85;
  assign n1808 = v2 & n1807;
  assign n1809 = ~v11 & n1808;
  assign n1810 = ~v9 & n1809;
  assign n1811 = v10 & n1810;
  assign n1812 = v15 & n1803;
  assign n1813 = ~v3 & n1812;
  assign n1814 = ~v13 & n1813;
  assign n1815 = ~v10 & n1808;
  assign n1816 = ~v8 & n1815;
  assign n1817 = v9 & n1816;
  assign n1818 = v7 & n632;
  assign n1819 = ~v14 & n1818;
  assign n1820 = v12 & n1819;
  assign n1821 = ~v12 & n632;
  assign n1822 = v7 & n1821;
  assign n1823 = ~v15 & n1822;
  assign n1824 = v13 & n1823;
  assign n1825 = v14 & n1824;
  assign n1826 = v15 & n1818;
  assign n1827 = v12 & n1826;
  assign n1828 = ~n1825 & ~n1827;
  assign n1829 = ~n1820 & n1828;
  assign n1830 = ~n1817 & n1829;
  assign n1831 = ~n1814 & n1830;
  assign n1832 = ~n1811 & n1831;
  assign n1833 = ~n1806 & n1832;
  assign n1834 = v14 & n1357;
  assign n1835 = v12 & n1834;
  assign n1836 = n361 & n1835;
  assign n1837 = n202 & n1703;
  assign n1838 = v7 & n1837;
  assign n1839 = v4 & n1838;
  assign n1840 = n160 & n1703;
  assign n1841 = v7 & n1840;
  assign n1842 = v4 & n1841;
  assign n1843 = ~v14 & ~v3;
  assign n1844 = v12 & n1843;
  assign n1845 = v2 & n1844;
  assign n1846 = ~v0 & n1845;
  assign n1847 = v1 & n1846;
  assign n1848 = ~n1842 & ~n1847;
  assign n1849 = ~n1839 & n1848;
  assign n1850 = ~n1836 & n1849;
  assign n1851 = ~v15 & n94;
  assign n1852 = v14 & n1851;
  assign n1853 = n1808 & n1852;
  assign n1854 = v12 & n1813;
  assign n1855 = v11 & n1808;
  assign n1856 = ~v8 & n1855;
  assign n1857 = v9 & n1856;
  assign n1858 = v8 & n1809;
  assign n1859 = v10 & n1858;
  assign n1860 = ~n1857 & ~n1859;
  assign n1861 = ~n1854 & n1860;
  assign n1862 = ~n1853 & n1861;
  assign n1863 = ~v5 & n1840;
  assign n1864 = v7 & n1863;
  assign n1865 = ~v6 & n1837;
  assign n1866 = v4 & n1865;
  assign n1867 = ~v5 & n1837;
  assign n1868 = v7 & n1867;
  assign n1869 = n1297 & n1658;
  assign n1870 = ~v15 & n1869;
  assign n1871 = v14 & n1870;
  assign n1872 = n1303 & n1658;
  assign n1873 = ~v15 & n1872;
  assign n1874 = v14 & n1873;
  assign n1875 = n432 & n1658;
  assign n1876 = ~v15 & n1875;
  assign n1877 = v14 & n1876;
  assign n1878 = n202 & n239;
  assign n1879 = n658 & n1878;
  assign n1880 = n805 & n1879;
  assign n1881 = ~n1877 & ~n1880;
  assign n1882 = ~n1874 & n1881;
  assign n1883 = ~n1871 & n1882;
  assign n1884 = ~n1868 & n1883;
  assign n1885 = ~n1866 & n1884;
  assign n1886 = ~n1864 & n1885;
  assign n1887 = n1862 & n1886;
  assign n1888 = n1850 & n1887;
  assign n1889 = n1833 & n1888;
  assign n1890 = n1801 & n1889;
  assign n1891 = n1786 & n1890;
  assign n1892 = v0 & v3;
  assign n1893 = ~v13 & n1892;
  assign n1894 = ~v14 & n1893;
  assign n1895 = ~v9 & n1892;
  assign n1896 = ~v11 & n1895;
  assign n1897 = v10 & n1896;
  assign n1898 = ~v8 & n1892;
  assign n1899 = ~v10 & n1898;
  assign n1900 = v9 & n1899;
  assign n1901 = ~v1 & v3;
  assign n1902 = ~v14 & n1901;
  assign n1903 = v12 & n1902;
  assign n1904 = ~n1900 & ~n1903;
  assign n1905 = ~n1897 & n1904;
  assign n1906 = ~n1894 & n1905;
  assign n1907 = v13 & ~v15;
  assign n1908 = v14 & n1907;
  assign n1909 = ~v12 & n1908;
  assign n1910 = ~v1 & n1909;
  assign n1911 = v3 & n1910;
  assign n1912 = v15 & n1901;
  assign n1913 = v12 & n1912;
  assign n1914 = v11 & v9;
  assign n1915 = ~v8 & n1914;
  assign n1916 = ~v1 & n1915;
  assign n1917 = v3 & n1916;
  assign n1918 = ~v1 & v8;
  assign n1919 = v3 & n1918;
  assign n1920 = ~v11 & n1919;
  assign n1921 = v10 & n1920;
  assign n1922 = ~n1917 & ~n1921;
  assign n1923 = ~n1913 & n1922;
  assign n1924 = ~n1911 & n1923;
  assign n1925 = ~v14 & n1892;
  assign n1926 = v12 & n1925;
  assign n1927 = ~v12 & v0;
  assign n1928 = v3 & n1927;
  assign n1929 = ~v15 & n1928;
  assign n1930 = v13 & n1929;
  assign n1931 = v14 & n1930;
  assign n1932 = ~v5 & ~v7;
  assign n1933 = v6 & n1932;
  assign n1934 = ~v10 & n1933;
  assign n1935 = ~v8 & n1934;
  assign n1936 = v9 & n1935;
  assign n1937 = v15 & n1892;
  assign n1938 = v12 & n1937;
  assign n1939 = v0 & ~v8;
  assign n1940 = v3 & n1939;
  assign n1941 = v9 & n1940;
  assign n1942 = v11 & n1941;
  assign n1943 = v10 & ~v11;
  assign n1944 = v8 & n1943;
  assign n1945 = v0 & n1944;
  assign n1946 = v3 & n1945;
  assign n1947 = v15 & n1893;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~n1942 & n1948;
  assign n1950 = ~n1938 & n1949;
  assign n1951 = ~n1936 & n1950;
  assign n1952 = ~n1931 & n1951;
  assign n1953 = ~n1926 & n1952;
  assign n1954 = ~v14 & n1933;
  assign n1955 = v12 & n1954;
  assign n1956 = ~v5 & v6;
  assign n1957 = ~v7 & n1956;
  assign n1958 = ~v12 & n1957;
  assign n1959 = ~v15 & n1958;
  assign n1960 = v13 & n1959;
  assign n1961 = v14 & n1960;
  assign n1962 = v15 & n1933;
  assign n1963 = v12 & n1962;
  assign n1964 = v11 & n1933;
  assign n1965 = ~v8 & n1964;
  assign n1966 = v9 & n1965;
  assign n1967 = ~n1963 & ~n1966;
  assign n1968 = ~n1961 & n1967;
  assign n1969 = ~n1955 & n1968;
  assign n1970 = ~v11 & n1933;
  assign n1971 = v8 & n1970;
  assign n1972 = v10 & n1971;
  assign n1973 = ~v13 & n1933;
  assign n1974 = v15 & n1973;
  assign n1975 = ~v13 & ~v14;
  assign n1976 = ~v7 & n1975;
  assign n1977 = ~v5 & n1976;
  assign n1978 = v6 & n1977;
  assign n1979 = ~v9 & n1970;
  assign n1980 = v10 & n1979;
  assign n1981 = ~n1978 & ~n1980;
  assign n1982 = ~n1974 & n1981;
  assign n1983 = ~n1972 & n1982;
  assign n1984 = ~v4 & ~v6;
  assign n1985 = v5 & n1984;
  assign n1986 = v11 & n1985;
  assign n1987 = ~v8 & n1986;
  assign n1988 = v9 & n1987;
  assign n1989 = ~v11 & n1985;
  assign n1990 = v8 & n1989;
  assign n1991 = v10 & n1990;
  assign n1992 = v15 & n1985;
  assign n1993 = v12 & n1992;
  assign n1994 = ~v13 & n1792;
  assign n1995 = v15 & n1994;
  assign n1996 = ~v14 & n1994;
  assign n1997 = ~v9 & n1989;
  assign n1998 = v10 & n1997;
  assign n1999 = ~v10 & n1985;
  assign n2000 = ~v8 & n1999;
  assign n2001 = v9 & n2000;
  assign n2002 = ~n1998 & ~n2001;
  assign n2003 = ~n1996 & n2002;
  assign n2004 = ~n1995 & n2003;
  assign n2005 = ~n1993 & n2004;
  assign n2006 = ~n1991 & n2005;
  assign n2007 = ~n1988 & n2006;
  assign n2008 = n1983 & n2007;
  assign n2009 = n1969 & n2008;
  assign n2010 = n1953 & n2009;
  assign n2011 = n1924 & n2010;
  assign n2012 = n1906 & n2011;
  assign n2013 = v4 & ~v7;
  assign n2014 = v6 & n2013;
  assign n2015 = v11 & n2014;
  assign n2016 = ~v8 & n2015;
  assign n2017 = v9 & n2016;
  assign n2018 = ~v11 & n2014;
  assign n2019 = v8 & n2018;
  assign n2020 = v10 & n2019;
  assign n2021 = v4 & v6;
  assign n2022 = ~v7 & n2021;
  assign n2023 = ~v13 & n2022;
  assign n2024 = v15 & n2023;
  assign n2025 = ~v14 & n2023;
  assign n2026 = ~n2024 & ~n2025;
  assign n2027 = ~n2020 & n2026;
  assign n2028 = ~n2017 & n2027;
  assign n2029 = ~v9 & n2018;
  assign n2030 = v10 & n2029;
  assign n2031 = ~v10 & n2014;
  assign n2032 = ~v8 & n2031;
  assign n2033 = v9 & n2032;
  assign n2034 = v0 & ~v2;
  assign n2035 = ~v14 & n2034;
  assign n2036 = v12 & n2035;
  assign n2037 = ~v2 & n1909;
  assign n2038 = v0 & n2037;
  assign n2039 = ~n2036 & ~n2038;
  assign n2040 = ~n2033 & n2039;
  assign n2041 = ~n2030 & n2040;
  assign n2042 = ~v13 & n1901;
  assign n2043 = ~v14 & n2042;
  assign n2044 = ~v9 & n1943;
  assign n2045 = ~v1 & n2044;
  assign n2046 = v3 & n2045;
  assign n2047 = v15 & n2042;
  assign n2048 = ~v1 & ~v8;
  assign n2049 = v3 & n2048;
  assign n2050 = ~v10 & n2049;
  assign n2051 = v9 & n2050;
  assign n2052 = v12 & ~v14;
  assign n2053 = ~v7 & n2052;
  assign n2054 = v4 & n2053;
  assign n2055 = v6 & n2054;
  assign n2056 = ~v12 & n2022;
  assign n2057 = ~v15 & n2056;
  assign n2058 = v13 & n2057;
  assign n2059 = v14 & n2058;
  assign n2060 = v15 & n2014;
  assign n2061 = v12 & n2060;
  assign n2062 = ~n2059 & ~n2061;
  assign n2063 = ~n2055 & n2062;
  assign n2064 = ~n2051 & n2063;
  assign n2065 = ~n2047 & n2064;
  assign n2066 = ~n2046 & n2065;
  assign n2067 = ~n2043 & n2066;
  assign n2068 = v15 & n2034;
  assign n2069 = v12 & n2068;
  assign n2070 = ~v2 & ~v8;
  assign n2071 = v0 & n2070;
  assign n2072 = v9 & n2071;
  assign n2073 = v11 & n2072;
  assign n2074 = ~v2 & n1944;
  assign n2075 = v0 & n2074;
  assign n2076 = ~v13 & n2034;
  assign n2077 = v15 & n2076;
  assign n2078 = ~n2075 & ~n2077;
  assign n2079 = ~n2073 & n2078;
  assign n2080 = ~n2069 & n2079;
  assign n2081 = ~v14 & n2076;
  assign n2082 = ~v2 & ~v9;
  assign n2083 = v0 & n2082;
  assign n2084 = ~v11 & n2083;
  assign n2085 = v10 & n2084;
  assign n2086 = ~v10 & n2071;
  assign n2087 = v9 & n2086;
  assign n2088 = ~v1 & ~v2;
  assign n2089 = ~v14 & n2088;
  assign n2090 = v12 & n2089;
  assign n2091 = ~n2087 & ~n2090;
  assign n2092 = ~n2085 & n2091;
  assign n2093 = ~n2081 & n2092;
  assign n2094 = ~v12 & ~v1;
  assign n2095 = ~v2 & n2094;
  assign n2096 = ~v15 & n2095;
  assign n2097 = v13 & n2096;
  assign n2098 = v14 & n2097;
  assign n2099 = v15 & n2088;
  assign n2100 = v12 & n2099;
  assign n2101 = ~v2 & n2048;
  assign n2102 = v9 & n2101;
  assign n2103 = v11 & n2102;
  assign n2104 = v8 & n2088;
  assign n2105 = ~v11 & n2104;
  assign n2106 = v10 & n2105;
  assign n2107 = ~n2103 & ~n2106;
  assign n2108 = ~n2100 & n2107;
  assign n2109 = ~n2098 & n2108;
  assign n2110 = ~v13 & n2088;
  assign n2111 = v15 & n2110;
  assign n2112 = ~v14 & n2110;
  assign n2113 = ~v1 & ~v9;
  assign n2114 = ~v2 & n2113;
  assign n2115 = ~v11 & n2114;
  assign n2116 = v10 & n2115;
  assign n2117 = ~v10 & n2101;
  assign n2118 = v9 & n2117;
  assign n2119 = ~n2116 & ~n2118;
  assign n2120 = ~n2112 & n2119;
  assign n2121 = ~n2111 & n2120;
  assign n2122 = n2109 & n2121;
  assign n2123 = n2093 & n2122;
  assign n2124 = n2080 & n2123;
  assign n2125 = n2067 & n2124;
  assign n2126 = n2041 & n2125;
  assign n2127 = n2028 & n2126;
  assign n2128 = n2012 & n2127;
  assign n2129 = n1891 & n2128;
  assign n2130 = n1772 & n2129;
  assign n2131 = n1656 & n2130;
  assign n2132 = n1148 & n2131;
  assign \v16.0  = ~n650 | ~n2132;
endmodule


