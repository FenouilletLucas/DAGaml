// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:52 2016

module TOP ( clock, 
    Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746, Pg6745,
    Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116, Pg115,
    Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, Pg72, Pg64,
    Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, PCLK,
    Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919, Pg34917,
    Pg34915, Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436, Pg34435,
    Pg34425, Pg34383, Pg34240, Pg34239, Pg34238, Pg34237, Pg34236, Pg34235,
    Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, Pg33959, Pg33950, Pg33949,
    Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874, Pg33659,
    Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429, Pg32185,
    Pg31863, Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656, Pg31521,
    Pg30332, Pg30331, Pg30330, Pg30329, Pg30327, Pg29221, Pg29220, Pg29219,
    Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, Pg29213, Pg29212, Pg29211,
    Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877, Pg26876,
    Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586, Pg25585,
    Pg25584, Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114, Pg24185,
    Pg24184, Pg24183, Pg24182, Pg24181, Pg24180, Pg24179, Pg24178, Pg24177,
    Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, Pg24171, Pg24170, Pg24169,
    Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162, Pg24161,
    Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002, Pg21727,
    Pg21698, Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899, Pg20763,
    Pg20654, Pg20652, Pg20557, Pg20049, Pg19357, Pg19334, Pg18881, Pg18101,
    Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, Pg18095, Pg18094, Pg18092,
    Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764, Pg17760,
    Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685, Pg17678,
    Pg17674, Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580, Pg17577,
    Pg17519, Pg17423, Pg17404, Pg17400, Pg17320, Pg17316, Pg17291, Pg16955,
    Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, Pg16722, Pg16718, Pg16693,
    Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828, Pg14779,
    Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635, Pg14597,
    Pg14518, Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167, Pg14147,
    Pg14125, Pg14096, Pg13966, Pg13926, Pg13906, Pg13895, Pg13881, Pg13865,
    Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, Pg13049, Pg13039, Pg12923,
    Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350, Pg12300,
    Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388, Pg11349,
    Pg10527, Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741, Pg9682,
    Pg9680, Pg9617, Pg9615, Pg9555, Pg9553, Pg9497, Pg9251, Pg9048, Pg9019,
    Pg8920, Pg8919, Pg8918, Pg8917, Pg8916, Pg8915, Pg8870, Pg8839, Pg8789,
    Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, Pg8783, Pg8719, Pg8475, Pg8416,
    Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, Pg8291, Pg8283, Pg8279,
    Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, Pg7540, Pg7260,
    Pg7257, Pg7245, Pg7243  );
  input  clock;
  input  Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746,
    Pg6745, Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116,
    Pg115, Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, Pg72,
    Pg64, Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, PCLK;
  output Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919,
    Pg34917, Pg34915, Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436,
    Pg34435, Pg34425, Pg34383, Pg34240, Pg34239, Pg34238, Pg34237, Pg34236,
    Pg34235, Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, Pg33959, Pg33950,
    Pg33949, Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874,
    Pg33659, Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429,
    Pg32185, Pg31863, Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656,
    Pg31521, Pg30332, Pg30331, Pg30330, Pg30329, Pg30327, Pg29221, Pg29220,
    Pg29219, Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, Pg29213, Pg29212,
    Pg29211, Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877,
    Pg26876, Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586,
    Pg25585, Pg25584, Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114,
    Pg24185, Pg24184, Pg24183, Pg24182, Pg24181, Pg24180, Pg24179, Pg24178,
    Pg24177, Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, Pg24171, Pg24170,
    Pg24169, Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162,
    Pg24161, Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002,
    Pg21727, Pg21698, Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899,
    Pg20763, Pg20654, Pg20652, Pg20557, Pg20049, Pg19357, Pg19334, Pg18881,
    Pg18101, Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, Pg18095, Pg18094,
    Pg18092, Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764,
    Pg17760, Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685,
    Pg17678, Pg17674, Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580,
    Pg17577, Pg17519, Pg17423, Pg17404, Pg17400, Pg17320, Pg17316, Pg17291,
    Pg16955, Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, Pg16722, Pg16718,
    Pg16693, Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828,
    Pg14779, Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635,
    Pg14597, Pg14518, Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167,
    Pg14147, Pg14125, Pg14096, Pg13966, Pg13926, Pg13906, Pg13895, Pg13881,
    Pg13865, Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, Pg13049, Pg13039,
    Pg12923, Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350,
    Pg12300, Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388,
    Pg11349, Pg10527, Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741,
    Pg9682, Pg9680, Pg9617, Pg9615, Pg9555, Pg9553, Pg9497, Pg9251, Pg9048,
    Pg9019, Pg8920, Pg8919, Pg8918, Pg8917, Pg8916, Pg8915, Pg8870, Pg8839,
    Pg8789, Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, Pg8783, Pg8719, Pg8475,
    Pg8416, Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, Pg8291, Pg8283,
    Pg8279, Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, Pg7540,
    Pg7260, Pg7257, Pg7245, Pg7243;
  reg Ng5057, Ng2771, Ng1882, Ng2299, Ng4040, Ng2547, Ng559, Ng3243, Ng452,
    Ng3542, Ng5232, Ng5813, Ng2907, Ng1744, Ng5909, Ng1802, Ng3554, Ng6219,
    Ng807, Ng6031, Ng847, Ng976, Ng4172, Ng4372, Ng3512, Ng749, Ng3490,
    Pg12350, Ng4235, Ng1600, Ng1714, Pg14451, Ng3155, Ng2236, Ng4555,
    Ng3698, Ng1736, Ng1968, Ng4621, Ng5607, Ng2657, Pg12300, Ng490, Ng311,
    Ng772, Ng5587, Ng6177, Ng6377, Ng3167, Ng5615, Ng4567, Ng3457, Ng6287,
    Pg7946, Ng2563, Ng4776, Ng4593, Ng6199, Ng2295, Ng1384, Ng1339, Ng5180,
    Ng2844, Ng1024, Ng5591, Ng3598, Ng4264, Ng767, Ng5853, Pg13865, Ng2089,
    Ng4933, Ng4521, Ng5507, Pg16656, Ng6291, Ng294, Ng5559, Pg9617, Pg9741,
    Ng3813, Ng562, Ng608, Ng1205, Ng3909, Ng6259, Ng5905, Ng921, Ng2955,
    Ng203, Ng1099, Ng4878, Ng5204, Pg17604, Ng3606, Ng1926, Ng6215, Ng3586,
    Ng291, Ng4674, Ng3570, Pg9048, Pg17607, Ng1862, Ng676, Ng843, Ng4332,
    Ng4153, Pg17711, Ng6336, Ng622, Ng3506, Ng4558, Pg17685, Ng3111,
    \[4430] , Ng26936, Ng939, Ng278, Ng4492, Ng4864, Ng1036, \[4427] ,
    Ng1178, Ng3239, Ng718, Ng6195, Ng1135, Ng6395, \[4415] , Ng554, Ng496,
    Ng3853, Ng5134, Pg17404, Pg8344, Ng2485, Ng925, Ng48, Ng5555, Pg14096,
    Ng1798, Ng4076, Ng2941, Ng3905, Ng763, Ng6255, Ng4375, Ng4871, Ng4722,
    Ng590, Pg13099, Ng1632, Pg12238, Ng3100, Ng1495, Ng1437, Ng6154,
    Ng1579, Ng5567, Ng1752, Ng1917, Ng744, Ng4737, \[4661] , Ng6267,
    Pg16659, Ng1442, Ng5965, Ng4477, Pg10500, Ng4643, Ng5264, Pg14779,
    Ng2610, Ng5160, Ng5933, Ng1454, Ng753, Ng1296, Ng3151, Ng2980, Ng6727,
    Ng3530, Ng4104, Ng1532, Pg9251, Ng2177, Ng52, Ng4754, Ng1189, Ng2287,
    Ng4273, Ng1389, Ng1706, Ng5835, Ng1171, Ng4269, Ng2399, Ng4983, Ng5611,
    Pg16627, Ng4572, Ng3143, Ng2898, Ng3343, Ng3235, Ng4543, Ng3566,
    Ng4534, Ng4961, Ng4927, Ng2259, Ng2819, Pg7257, Ng5802, Ng2852, Ng417,
    Ng681, Ng437, Ng351, Ng5901, Ng2886, Ng3494, Ng5511, Ng3518, Ng1604,
    Ng5092, Ng4831, Ng4382, Ng6386, Ng479, Ng3965, Ng4749, Ng2008, Ng736,
    Ng3933, Ng222, Ng3050, Ng1052, Pg17580, Ng2122, Ng2465, Ng5889, Ng4495,
    Pg8719, Ng4653, Ng3179, Ng1728, Ng2433, Ng3835, Ng6187, Ng4917, Ng1070,
    Ng822, Pg17715, Ng914, Ng5339, Ng4164, Ng969, Ng2807, Ng4054, Ng6191,
    Ng5077, Ng5523, Ng3680, Ng6637, Ng174, Ng1682, Ng355, Ng1087, Ng1105,
    Ng2342, Ng6307, Ng3802, Ng6159, Ng2255, Ng2815, Ng911, Ng43, Pg16775,
    Ng1748, Ng5551, Ng3558, Ng5499, Ng2960, Ng3901, Ng4888, Ng6251,
    Pg17649, Ng1373, Pg8215, Ng157, Ng2783, Ng4281, Ng3574, Ng2112, Ng1283,
    Ng433, Ng4297, Pg14738, Pg13272, Ng758, Ng4639, Ng6537, Ng5543, Pg8475,
    Ng5961, Ng6243, Ng632, Pg12919, Ng3889, Ng3476, Ng1664, Ng1246, Ng6629,
    Ng246, Ng4049, Pg7260, Ng2932, Ng4575, Ng4098, Ng4498, Ng528, Ng16,
    Ng3139, \[4432] , Ng4584, Ng142, Pg17639, Ng5831, Ng239, Ng1216,
    Ng2848, Ng5022, Pg16955, Ng1030, Pg13881, Ng3231, Pg9817, Ng1430,
    Ng4452, Ng2241, Ng1564, Pg9680, Ng6148, Ng6649, Ng110, Pg14147, Ng225,
    Ng4486, Ng4504, Ng5873, Ng5037, Ng2319, Ng5495, Pg11770, Ng5208,
    Ng5579, Ng5869, Ng1589, Ng5752, Ng6279, Ng5917, Ng2975, Ng6167,
    Pg13966, Ng2599, Ng1448, Pg14125, Ng2370, Ng5164, Ng1333, Ng153,
    Ng6549, Ng4087, Ng4801, Ng2984, Ng3961, Ng962, Ng101, Pg8918, Ng6625,
    Ng51, Ng1018, Pg17320, Ng4045, Ng1467, Ng2461, Ng2756, Ng5990, Ng1256,
    Ng5029, Ng6519, Ng1816, Ng4369, Ng4578, Ng4459, Ng3831, Ng2514, Ng3288,
    Ng2403, Ng2145, Ng1700, Ng513, Ng2841, Ng5297, Ng2763, Ng4793, Ng952,
    Ng1263, Ng1950, Ng5138, Ng2307, Ng5109, Pg8398, Ng4664, Ng2223, Ng5808,
    Ng6645, Ng2016, Ng3873, Pg13926, Ng2315, Ng2811, Ng5957, Ng2047,
    Ng3869, Pg17760, Ng5575, Ng46, Ng3752, Ng3917, Pg8783, Ng1585, Ng4388,
    Ng6275, Ng6311, Pg8916, Ng1041, Ng2595, Ng2537, \[4426] , Ng4430,
    Ng4564, Ng4826, Ng6239, Ng232, Ng5268, Ng6545, Ng2417, Ng1772, Ng5052,
    Pg9615, Ng1890, Ng2629, Ng572, Ng2130, Ng4108, Ng4308, Ng475, Ng990,
    Ng45, Pg12184, Ng3990, Ng5881, Ng1992, Ng3171, Ng812, Ng832, Ng5897,
    Ng4571, Pg13895, Ng4455, Ng2902, Ng333, Ng168, Ng2823, Ng3684, Ng3639,
    Pg14597, Ng3338, Ng5406, Ng269, Ng401, Ng6040, Ng441, Pg9553, Ng3808,
    Ng10384, Ng3957, Ng4093, Ng1760, Pg12422, Ng160, Ng2279, Ng3498, Ng586,
    Pg14201, Ng2619, Ng1183, Ng1608, Pg8785, Pg17577, Ng1779, Ng2652,
    Ng2193, Ng2393, Ng661, Ng4950, Ng5535, Ng2834, Ng1361, Ng6235, Ng1146,
    Ng2625, Ng150, Ng1696, Ng6555, Pg14189, Ng3881, Ng6621, Ng3470, Ng3897,
    Ng518, Ng538, Ng2606, Ng1472, Ng542, Ng5188, Ng5689, Pg13259, Ng405,
    Ng5216, Ng6494, Ng4669, Ng996, Ng4531, Ng2860, Ng4743, Ng6593, Pg8291,
    Ng4411, Ng1413, Ng26960, Pg13039, Ng6641, Ng1936, Ng55, Ng504, Ng2587,
    Ng4480, Ng2311, Ng3602, Ng5571, Ng3578, Pg9555, Ng5827, Ng3582, Ng6271,
    Ng4688, Ng2380, Ng5196, Ng3227, Ng2020, Pg14518, Pg17316, Ng6541,
    Ng3203, Ng1668, Ng4760, Ng262, Ng1840, Ng5467, Ng460, Ng6209, \[4436] ,
    Pg14662, Ng655, Ng3502, Ng2204, Ng5256, Ng4608, Ng794, Pg13906, Ng4423,
    Ng3689, Ng5685, Ng703, Ng862, Ng3247, Ng2040, Ng4146, Ng4633, Pg7916,
    Ng4732, Pg9497, Ng5817, Ng2351, Ng2648, Ng6736, Ng4944, Ng4072, Pg7540,
    Ng4443, Ng3466, Ng4116, Ng5041, Ng4434, Ng3827, Ng6500, Pg17813,
    Ng3133, Ng3333, Ng979, Ng4681, Ng298, Ng2667, Pg8789, Ng1894, Ng2988,
    Ng3538, Ng301, Ng341, Ng827, Pg17291, Ng2555, Ng5011, Ng199, Ng6523,
    Ng1526, Ng4601, Ng854, Ng1484, Ng4922, Ng5080, Ng5863, Ng4581, Ng2518,
    Ng2567, Ng568, Ng3263, Ng6613, Ng6044, Ng6444, Ng2965, Ng5857, Ng1616,
    Ng890, Pg17646, Ng3562, Pg10122, Ng1404, Ng3817, Ng93, Ng4501, Ng287,
    Ng2724, Ng4704, Ng22, Ng2878, Ng5220, Ng617, Pg12368, Ng316, Ng1277,
    Ng6513, Ng336, Ng2882, Ng933, Ng1906, Ng305, Ng8, Ng2799, Pg14167,
    Pg17787, Ng4912, Ng4157, Ng2541, Ng2153, Ng550, Ng255, Ng1945, Ng5240,
    Ng1478, Ng3863, Ng1959, Ng3480, Ng6653, Pg17764, Ng2864, Ng4894,
    Pg17678, Ng3857, Pg16693, Ng499, Ng1002, Ng776, Ng1236, Ng4646, Ng2476,
    Ng1657, Ng2375, Ng63, Pg17739, Ng358, Ng896, Ng283, Ng3161, Ng2384,
    Pg14828, Ng4616, Ng4561, Ng2024, Ng3451, Ng2795, Ng613, Ng4527, Ng1844,
    Ng5937, Ng4546, Ng2523, Pg11349, Ng2643, Ng1489, Pg8358, Ng2551,
    Ng5156, \[4421] , Pg8279, Pg8839, Ng1955, Ng6049, Ng2273, Pg14749,
    Ng4771, Ng6098, Ng3147, Ng3347, Ng2269, Ng191, Ng2712, Ng626, Ng2729,
    Ng5357, Ng4991, Pg17819, Ng4709, Ng2927, Ng4340, Ng5929, Ng4907,
    Pg16874, Ng4035, Ng2946, Ng918, Ng4082, Pg9743, Ng2036, Ng577, Ng1620,
    Ng2831, Ng667, Ng930, Ng3937, Ng817, Ng1249, Ng837, Pg16924, Ng599,
    Ng5475, Ng739, Ng5949, Ng6682, Ng904, Ng2873, Ng1854, Ng5084, Ng5603,
    Pg8870, Ng2495, Ng2437, Ng2102, Ng2208, Ng2579, Ng4064, Ng4899, Ng2719,
    Ng4785, Ng5583, Ng781, Ng6173, Pg17743, Ng2917, Ng686, Ng1252, Ng671,
    Ng2265, Ng6283, Pg14705, Pg17519, Pg8784, Ng5527, Ng4489, Ng1974,
    Ng1270, Ng4966, Ng6227, Ng3929, Ng5503, Ng4242, Ng5925, Ng1124, Ng4955,
    Ng5224, Ng2012, Ng6203, Ng5120, Pg17674, Ng2389, Ng4438, Ng2429,
    Ng2787, Ng1287, Ng2675, \[4507] , Ng4836, Ng1199, Pg19357, Ng5547,
    Ng2138, Pg16744, Ng2338, Pg8919, Ng6247, Ng2791, Ng3949, Ng1291,
    Ng5945, Ng5244, Ng2759, Ng6741, Ng785, Ng1259, Ng3484, Ng209, Ng6609,
    Ng5517, Ng2449, Ng2575, Ng65, Ng2715, Ng936, Ng2098, Ng4462, Ng604,
    Ng6589, Ng1886, Pg17845, Pg17871, Ng429, Ng1870, Ng4249, Ng1825,
    Ng1008, Ng4392, Ng3546, Ng5236, Ng1768, Ng4854, Ng3925, Ng6509, Ng732,
    Ng2504, Ng1322, Ng4520, Pg8917, Ng2185, Ng37, Ng4031, Ng2070, \[4658] ,
    Ng4176, Pg11418, Ng4405, Ng872, Ng6181, Ng6381, Ng4765, Ng5563, Ng1395,
    Ng1913, Ng2331, Ng6263, Ng50, Ng3945, Ng347, Ng4473, Ng1266, Ng5489,
    Ng714, Ng2748, Ng5471, Ng4540, Ng6723, Ng6605, Ng2445, Ng2173, Pg9019,
    Ng2491, Ng4849, Ng2169, Ng2283, Ng6585, \[4428] , Ng2407, Ng2868,
    Ng2767, Ng1783, Pg16718, Ng1312, Ng5212, Ng4245, Ng645, Ng4291,
    \[4435] , Ng182, Ng1129, Ng2227, Pg8788, Ng2246, Ng1830, Ng3590, Ng392,
    Ng1592, Ng6505, Ng1221, Ng5921, \[4431] , Ng146, Ng218, Ng1932, Ng1624,
    Ng5062, Ng5462, Ng2689, Ng6573, Ng1677, Ng2028, Ng2671, Pg10527,
    Pg7243, Ng1848, \[4434] , Ng5485, Ng2741, Pg11678, Ng2638, Ng4122,
    Ng4322, Ng5941, Ng2108, Pg13068, Ng25, Ng1644, Ng595, Ng2217, Ng1319,
    Ng2066, Ng1152, Ng5252, Ng2165, Ng2571, Ng5176, Pg14673, Ng1211,
    Ng2827, Pg14217, Ng4859, Ng424, Ng1274, Pg17423, Ng85, Ng2803, Ng1821,
    Ng2509, Ng5073, Ng1280, \[4651] , Pg13085, Ng6633, Ng5124, Pg17400,
    Ng6303, Ng5069, Ng2994, Ng650, Ng1636, Ng3921, Ng2093, Ng6732, Ng1306,
    Ng1061, Ng3462, Ng2181, Ng956, Ng1756, Ng5849, Ng4112, Ng2685, Ng2197,
    Ng2421, Ng1046, Ng482, Ng4401, Ng1514, Ng329, Ng6565, Ng2950, Ng1345,
    Ng6533, Pg14421, Ng4727, Pg12470, Ng1536, Ng3941, Ng370, Ng5694,
    Ng1858, Ng446, Ng3219, Ng1811, Ng6601, Ng2441, Ng1874, Ng4349, Ng6581,
    Ng6597, Ng3610, Ng2890, Ng1978, Ng1612, Ng112, Ng2856, Ng1982, Pg17722,
    Ng5228, Ng4119, Ng6390, Ng1542, Ng4258, Ng4818, Ng5033, Ng4717, Ng1554,
    Ng3849, Pg17778, Ng3199, Ng5845, Ng4975, Ng790, Ng5913, Ng1902, Ng6163,
    Ng4125, Ng4821, Ng4939, Pg19334, Ng3207, Ng4483, Ng3259, Ng5142,
    Ng5248, Ng2126, Ng3694, Ng5481, Ng1964, Ng5097, Ng3215, Pg16748, Ng111,
    Ng4427, Ng2779, Pg8786, Pg7245, Ng1720, Ng1367, Ng5112, Ng4145, Ng2161,
    Ng376, Ng2361, Pg11447, Ng582, Ng2051, Ng1193, Ng2327, Ng907, Ng947,
    Ng1834, Ng3594, Ng2999, Ng2303, Pg17688, Ng699, Ng723, Ng5703, Ng546,
    Ng2472, Ng5953, Pg8277, Ng1740, Ng3550, Ng3845, Ng2116, Pg14635,
    Ng3195, Ng3913, Pg10306, Ng1687, Ng2681, Ng2533, Ng324, Ng2697, Ng4417,
    Ng6561, Ng1141, Pg12923, Ng2413, Ng1710, Ng6527, Ng3255, Ng1691,
    Ng2936, Ng5644, Ng5152, Ng5352, Pg8915, Ng2775, Ng2922, Ng1111, Ng5893,
    Pg16603, Ng6617, Ng2060, Ng4512, Ng5599, Ng3401, Ng4366, Pg16722,
    \[4433] , Ng3129, Ng3329, Ng5170, Ng26959, Ng5821, Ng6299, Pg8416,
    Ng2079, Ng4698, Ng3703, Ng1559, Ng943, Ng411, Pg9682, Ng3953, Ng2704,
    Ng6035, Ng1300, Ng4057, Ng5200, Ng4843, Ng5046, Ng2250, Ng26885,
    Ng4549, Ng2453, Ng5841, Pg14694, Ng2912, Ng2357, Pg8920, Ng164, Ng4253,
    Ng5016, Ng3119, Ng1351, Ng1648, Ng6972, Ng5115, Ng3352, Ng6657, Ng4552,
    Ng3893, Ng3211, Pg13049, Pg16624, Ng5595, Ng3614, Ng2894, Ng3125,
    Pg16686, Ng3821, Ng4141, Ng6974, Ng5272, Ng2735, Ng728, Ng6295, Ng2661,
    Ng1988, Ng5128, Ng1548, Ng3106, Ng4659, Ng4358, Ng1792, Ng2084, Ng3187,
    Ng4311, Ng2583, Ng3003, Ng1094, Ng3841, Ng4284, Ng3191, Ng4239, Ng4180,
    Ng691, Ng534, Ng385, Ng2004, Ng2527, Ng5456, Ng4420, Ng5148, Ng4507,
    Ng5348, Ng3223, Ng2970, Ng5698, Ng5260, Ng1521, Ng3522, Ng3115, Ng3251,
    Pg12832, Ng4628, Ng1996, Pg8342, Ng4515, Pg8787, Ng4300, Ng1724,
    Ng1379, Pg11388, Ng1878, Ng5619, Ng71, \[4437] ;
  wire n4125_1, n4126, n4127, n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143_1, n4144,
    n4145, n4146, n4147, n4148_1, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160, n4161_1, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
    n4175_1, n4176, n4177, n4178, n4179_1, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188_1, n4189, n4190, n4191, n4192,
    n4193_1, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207_1, n4208, n4209, n4210, n4211, n4212,
    n4213, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232_1, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240_1, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250_1, n4251, n4253, n4254,
    n4255_1, n4256, n4257, n4258, n4259, n4260_1, n4261, n4262, n4263,
    n4264_1, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
    n4273_1, n4274, n4275, n4276, n4277, n4278_1, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370_1, n4371, n4373, n4374,
    n4375_1, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390_1, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4408_1, n4409, n4410, n4411, n4412, n4413_1, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423_1, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438_1, n4439, n4440, n4441, n4442, n4443, n4445,
    n4446, n4447, n4448_1, n4449, n4450, n4451, n4452, n4453_1, n4454,
    n4455, n4456, n4457_1, n4458, n4459, n4460, n4461_1, n4462, n4463,
    n4464, n4465, n4466_1, n4467, n4468, n4469, n4470, n4471_1, n4472,
    n4473, n4474, n4475, n4476_1, n4478, n4479, n4480, n4481_1, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488, n4491, n4492, n4493_1, n4494,
    n4495, n4496_1, n4497, n4498, n4499, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4521, n4522, n4523, n4524, n4525_1, n4526,
    n4527, n4528, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545_1, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4554, n4555_1, n4556, n4557, n4558,
    n4560_1, n4561, n4562, n4563, n4565_1, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575_1, n4577, n4578, n4579_1,
    n4580, n4581, n4582, n4583_1, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598_1, n4599,
    n4600, n4602, n4604, n4605, n4606, n4607, n4608_1, n4609, n4610, n4611,
    n4612, n4613_1, n4614, n4615, n4616, n4617, n4618_1, n4619, n4620,
    n4621, n4624, n4625, n4626, n4627, n4628_1, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
    n4643, n4644, n4645_1, n4646, n4647, n4648, n4649_1, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657, n4658_1, n4659, n4660, n4661,
    n4662, n4663, n4665, n4666, n4667, n4668_1, n4669, n4670, n4672, n4674,
    n4675, n4676, n4677, n4678_1, n4679, n4680, n4682, n4683_1, n4684,
    n4685, n4686, n4687, n4688_1, n4689, n4690, n4692, n4693_1, n4695,
    n4697, n4698_1, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708_1, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
    n4718_1, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
    n4728_1, n4729, n4730, n4731, n4732_1, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4741, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4760, n4761,
    n4762_1, n4763, n4764, n4765, n4766, n4767, n4768, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788_1, n4789, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798_1, n4799, n4800, n4801, n4802, n4803_1,
    n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4820, n4822, n4823, n4824, n4825,
    n4826, n4828_1, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843_1, n4844, n4845, n4846,
    n4847_1, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865_1, n4866, n4867,
    n4868, n4869_1, n4870, n4871, n4873, n4874_1, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4889, n4890, n4891_1, n4892, n4893, n4894, n4895, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905_1, n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920_1, n4921,
    n4922, n4923, n4924, n4925_1, n4926, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974_1,
    n4975, n4976, n4977, n4978, n4979_1, n4980, n4981, n4982, n4983, n4984,
    n4985, n4986, n4987, n4988_1, n4989, n4990, n4992, n4993_1, n4994,
    n4995, n4996, n4997, n4998, n4999, n5001, n5002, n5003_1, n5004, n5005,
    n5006, n5007, n5008_1, n5009, n5010, n5011, n5012, n5014, n5015, n5016,
    n5017_1, n5018, n5019, n5020, n5021, n5022_1, n5024, n5025, n5026,
    n5027_1, n5028, n5029, n5031, n5032_1, n5033, n5034, n5035, n5036,
    n5037_1, n5038, n5039, n5041, n5042_1, n5043, n5044, n5045, n5046,
    n5047, n5048, n5050, n5051, n5052, n5054, n5055, n5057, n5058, n5059,
    n5060, n5061_1, n5062, n5063, n5064, n5065_1, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5077, n5078, n5079,
    n5080_1, n5081, n5082, n5083, n5084, n5085, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5095, n5096, n5097, n5098, n5099_1, n5100, n5101,
    n5103, n5104_1, n5105, n5106, n5107, n5108_1, n5109, n5110, n5111,
    n5112_1, n5114, n5115, n5116, n5117_1, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127_1, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
    n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5150, n5151, n5152,
    n5153, n5155, n5156, n5157_1, n5158, n5159, n5160, n5161_1, n5163,
    n5165, n5166_1, n5167, n5168, n5169, n5170, n5171_1, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191_1, n5192, n5193,
    n5194, n5195, n5196, n5197, n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5208, n5209, n5210, n5211, n5213, n5214, n5215, n5217,
    n5218, n5219, n5220, n5221, n5222, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
    n5251, n5252, n5253, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270_1, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279_1, n5280, n5282,
    n5283, n5284, n5285, n5286, n5288, n5289_1, n5290, n5291, n5292, n5293,
    n5294_1, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314_1, n5315,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5326, n5327,
    n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5341, n5342, n5343, n5344, n5345, n5346, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5365, n5366, n5368, n5369, n5370, n5371,
    n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5395, n5396, n5397, n5399, n5400, n5401, n5402, n5403, n5404, n5406,
    n5407, n5408, n5409, n5410, n5411, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432_1, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447_1,
    n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457_1,
    n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
    n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525, n5527, n5528, n5529, n5530,
    n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542_1, n5543, n5544, n5545, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5584, n5585,
    n5586, n5587, n5588, n5589, n5591, n5592, n5594_1, n5595, n5596, n5597,
    n5598, n5599, n5600, n5602, n5603, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624_1, n5625, n5627, n5628, n5629_1,
    n5630, n5631, n5632, n5634, n5635, n5636, n5637, n5638, n5639_1, n5640,
    n5641, n5643, n5645, n5646, n5647, n5649, n5650, n5651, n5652, n5655,
    n5656, n5657, n5658, n5659_1, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5668, n5669, n5670, n5671, n5672_1, n5673, n5674, n5675, n5676,
    n5677, n5678, n5680, n5681, n5684, n5685, n5686, n5687, n5688, n5689,
    n5691_1, n5692, n5693, n5694, n5695, n5696_1, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711_1, n5712, n5713, n5714, n5715, n5716, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5727, n5728, n5730, n5731, n5732, n5734,
    n5735, n5736, n5737, n5738, n5739_1, n5740, n5741, n5742, n5743, n5744,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759_1, n5760, n5762, n5763, n5764_1, n5766,
    n5767, n5768, n5769_1, n5770, n5771, n5772, n5773_1, n5775, n5776,
    n5777, n5778, n5779, n5780, n5782_1, n5783, n5784, n5785, n5786,
    n5787_1, n5788, n5790, n5791, n5792_1, n5793, n5795, n5796, n5797_1,
    n5798, n5799, n5800, n5801, n5802_1, n5803, n5804, n5805, n5807_1,
    n5808, n5809, n5811, n5812, n5813, n5814, n5815, n5817, n5818, n5820,
    n5821, n5822_1, n5823, n5824, n5825, n5826_1, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834_1, n5836, n5837, n5838, n5839_1, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5848, n5849, n5850, n5852,
    n5853, n5854, n5855, n5856_1, n5857, n5859, n5860, n5861, n5862, n5864,
    n5866, n5867, n5868, n5869, n5870, n5871, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889_1, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
    n5898, n5899_1, n5900, n5901, n5902, n5903, n5905, n5906, n5907, n5908,
    n5909_1, n5911, n5912, n5913, n5914_1, n5915, n5916, n5917, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929_1,
    n5931, n5932, n5933, n5934_1, n5935, n5936, n5937, n5938, n5939, n5940,
    n5942_1, n5943, n5944, n5945, n5946, n5947, n5948, n5950, n5952, n5953,
    n5955, n5956, n5957, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967_1, n5968, n5969, n5970, n5971, n5972_1, n5973, n5974,
    n5975, n5976_1, n5977, n5978, n5979, n5982, n5983, n5984, n5986, n5988,
    n5989, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009_1, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6018_1, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027, n6028_1, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037, n6038_1, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053_1, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067_1, n6068, n6069, n6070, n6071,
    n6072, n6074, n6075, n6076, n6077, n6078, n6079, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087_1, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6099, n6100, n6101_1, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110_1, n6111, n6113, n6114, n6115, n6116, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6127, n6128, n6129,
    n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138_1, n6139, n6142,
    n6143_1, n6144, n6145, n6148_1, n6149, n6150, n6151, n6152, n6153_1,
    n6154, n6155, n6156, n6158, n6159, n6160, n6161_1, n6162, n6163, n6164,
    n6165, n6166_1, n6167, n6168, n6169, n6170_1, n6172, n6173, n6174,
    n6175_1, n6176, n6177, n6178, n6179, n6180_1, n6182, n6183, n6184_1,
    n6185, n6186, n6187, n6188, n6189_1, n6190, n6191, n6192, n6193_1,
    n6194, n6195, n6197_1, n6198, n6199, n6200, n6201, n6202_1, n6203,
    n6204, n6205, n6206, n6208, n6209, n6210, n6211, n6213, n6214, n6215,
    n6216, n6217_1, n6218, n6219, n6221, n6222_1, n6223, n6224, n6226,
    n6227_1, n6228, n6229, n6230, n6231_1, n6232, n6233, n6236_1, n6239,
    n6240, n6242, n6243, n6244, n6245, n6247, n6248, n6249, n6250, n6251,
    n6252, n6253, n6254, n6255, n6256, n6258, n6259, n6260, n6261, n6262,
    n6264, n6265, n6266_1, n6267, n6268, n6270, n6271_1, n6272, n6273,
    n6274, n6275, n6276_1, n6277, n6278, n6279, n6280_1, n6281, n6283,
    n6284, n6285_1, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6294_1, n6295, n6296, n6297, n6298_1, n6299, n6300, n6301, n6302,
    n6303_1, n6304, n6305, n6306, n6307_1, n6308, n6309, n6310, n6311_1,
    n6312, n6313, n6314, n6315, n6316_1, n6317, n6318, n6319, n6320,
    n6321_1, n6322, n6323, n6324, n6325, n6326_1, n6327, n6328, n6329,
    n6330, n6331_1, n6332, n6333, n6334, n6335, n6336_1, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344, n6345_1, n6346, n6347, n6348,
    n6349, n6350_1, n6351, n6352, n6353, n6354, n6355_1, n6357, n6358,
    n6359, n6360_1, n6361, n6362, n6364, n6365_1, n6366, n6367, n6368,
    n6369, n6370_1, n6372, n6373, n6374_1, n6376, n6377_1, n6378, n6379,
    n6381_1, n6382, n6385, n6386, n6387, n6388, n6389, n6390, n6391_1,
    n6392, n6394, n6395, n6397, n6398, n6399, n6400_1, n6402, n6403,
    n6404_1, n6405, n6406, n6408, n6409_1, n6411, n6412, n6413, n6414_1,
    n6415, n6416, n6417, n6419, n6420, n6421, n6422, n6423_1, n6426, n6427,
    n6428_1, n6429, n6430, n6431, n6432, n6433_1, n6435, n6436, n6437,
    n6438_1, n6439, n6440, n6441, n6442, n6443_1, n6444, n6445, n6447,
    n6448_1, n6449, n6451, n6452, n6453_1, n6456, n6457, n6458_1, n6460,
    n6461, n6462, n6463_1, n6464, n6465, n6466, n6467, n6469, n6471, n6472,
    n6473_1, n6475, n6476, n6477, n6478_1, n6479, n6480, n6481, n6482,
    n6483_1, n6485, n6486, n6487, n6488_1, n6489, n6492, n6493_1, n6494,
    n6495, n6496, n6497, n6498_1, n6499, n6500, n6501, n6502, n6503_1,
    n6504, n6505, n6506, n6507, n6508_1, n6509, n6510, n6512, n6513_1,
    n6514, n6515, n6516, n6517, n6518_1, n6519, n6520, n6522, n6523_1,
    n6524, n6525, n6526, n6528, n6529, n6530, n6531, n6532_1, n6533, n6534,
    n6536, n6537_1, n6538, n6539, n6540, n6541, n6542_1, n6543, n6545,
    n6546, n6547_1, n6548, n6549, n6550, n6552_1, n6553, n6555, n6556_1,
    n6557, n6558, n6559, n6560, n6561_1, n6562, n6563, n6564, n6565, n6567,
    n6568, n6569, n6570, n6571_1, n6572, n6573, n6574, n6575, n6576_1,
    n6577, n6578, n6579, n6580, n6581_1, n6582, n6584, n6585, n6586_1,
    n6588, n6589, n6591_1, n6592, n6593, n6594, n6595, n6596_1, n6597,
    n6598, n6600, n6601_1, n6602, n6603, n6604, n6605, n6607, n6608, n6609,
    n6610, n6611_1, n6612, n6613, n6614, n6615, n6616_1, n6617, n6618,
    n6619, n6620, n6621_1, n6622, n6623, n6624, n6625_1, n6626, n6627,
    n6628, n6629, n6630_1, n6631, n6632, n6633, n6634, n6635_1, n6636,
    n6637, n6638, n6640, n6641, n6642, n6643_1, n6644, n6645, n6647_1,
    n6648, n6650, n6651, n6652_1, n6653, n6654, n6655, n6656, n6658, n6659,
    n6660, n6661, n6662_1, n6663, n6664, n6666_1, n6667, n6668, n6670,
    n6671_1, n6672, n6673, n6674, n6675, n6677, n6678, n6679, n6680,
    n6681_1, n6682, n6683, n6684, n6685, n6686, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
    n6702, n6704, n6705, n6707, n6708, n6709, n6710, n6711, n6712, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6735, n6736,
    n6738, n6739, n6740, n6741, n6742, n6744, n6745, n6747, n6748, n6750,
    n6751, n6752, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6762,
    n6763, n6764, n6766, n6767, n6768, n6769, n6770, n6771, n6773, n6774,
    n6775, n6777, n6778, n6780, n6781, n6782, n6783, n6785, n6786, n6787,
    n6788, n6789, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
    n6870, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6880, n6881,
    n6882, n6883, n6884, n6885, n6887, n6888, n6889, n6890, n6892, n6893,
    n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6927, n6928, n6929, n6930, n6932, n6933, n6934, n6935, n6936, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6969, n6970, n6971,
    n6972, n6973, n6974, n6976, n6977, n6978, n6980, n6982, n6983, n6984,
    n6985, n6987, n6988, n6990, n6991, n6992, n6994, n6995, n6996, n6997,
    n6998, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7023, n7024, n7025, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7050, n7051, n7052, n7053, n7055,
    n7056, n7057, n7058, n7059, n7060, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7091, n7092, n7093, n7094, n7095, n7096, n7098, n7100, n7101,
    n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7111, n7112, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7126, n7127, n7128, n7129, n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7149, n7150, n7151, n7152, n7153, n7154, n7156, n7157, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7178, n7179, n7180, n7181, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189, n7191, n7192, n7193, n7194,
    n7195, n7196, n7198, n7199, n7200, n7201, n7202, n7203, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7213, n7214, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7224, n7225, n7226, n7227, n7228, n7229,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7284,
    n7285, n7286, n7287, n7288, n7289, n7291, n7292, n7293, n7294, n7295,
    n7296, n7298, n7299, n7300, n7302, n7303, n7304, n7305, n7307, n7308,
    n7309, n7310, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7321,
    n7322, n7323, n7324, n7325, n7326, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7344,
    n7345, n7346, n7347, n7348, n7349, n7351, n7352, n7354, n7355, n7356,
    n7357, n7358, n7359, n7361, n7362, n7363, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7378, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386, n7388, n7389, n7390, n7391,
    n7392, n7393, n7394, n7395, n7397, n7399, n7400, n7401, n7402, n7403,
    n7404, n7406, n7407, n7408, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7444, n7446, n7447,
    n7448, n7449, n7451, n7452, n7453, n7455, n7456, n7457, n7458, n7459,
    n7461, n7462, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
    n7472, n7473, n7475, n7476, n7477, n7478, n7479, n7481, n7482, n7483,
    n7484, n7486, n7487, n7488, n7489, n7490, n7491, n7493, n7494, n7495,
    n7496, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
    n7508, n7509, n7510, n7512, n7513, n7514, n7515, n7516, n7518, n7519,
    n7520, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7530, n7531,
    n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7546, n7547, n7548, n7549, n7550, n7551, n7553, n7554,
    n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7565, n7566,
    n7567, n7568, n7570, n7572, n7573, n7574, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7597, n7598, n7599, n7600, n7601,
    n7602, n7603, n7604, n7606, n7607, n7609, n7610, n7611, n7612, n7613,
    n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7632, n7633, n7635, n7637, n7638,
    n7639, n7640, n7641, n7643, n7644, n7645, n7646, n7647, n7648, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656, n7658, n7659, n7660, n7662,
    n7663, n7664, n7665, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
    n7674, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
    n7708, n7709, n7710, n7711, n7713, n7714, n7715, n7717, n7718, n7719,
    n7720, n7721, n7723, n7724, n7725, n7726, n7727, n7729, n7730, n7731,
    n7732, n7733, n7734, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
    n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7761, n7762, n7763, n7764, n7766,
    n7767, n7768, n7769, n7770, n7772, n7773, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7807, n7808, n7809, n7810, n7811,
    n7812, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
    n7857, n7858, n7860, n7862, n7863, n7864, n7865, n7866, n7867, n7869,
    n7870, n7871, n7872, n7873, n7874, n7876, n7877, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7891, n7892,
    n7893, n7894, n7895, n7896, n7898, n7899, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7910, n7911, n7912, n7913, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7924, n7925, n7926, n7927,
    n7928, n7929, n7931, n7932, n7934, n7935, n7937, n7938, n7939, n7940,
    n7941, n7942, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
    n7952, n7953, n7954, n7955, n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7973, n7974,
    n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7996, n7997,
    n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8006, n8007, n8008,
    n8009, n8010, n8011, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8029, n8030, n8031,
    n8032, n8033, n8034, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
    n8044, n8045, n8046, n8047, n8048, n8049, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8063, n8064, n8066,
    n8067, n8068, n8069, n8070, n8071, n8073, n8074, n8075, n8076, n8077,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8087, n8088, n8089,
    n8091, n8092, n8093, n8094, n8095, n8096, n8098, n8099, n8100, n8101,
    n8103, n8104, n8105, n8106, n8107, n8108, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8119, n8120, n8121, n8122, n8123, n8124,
    n8126, n8127, n8129, n8130, n8131, n8132, n8134, n8136, n8137, n8138,
    n8140, n8141, n8142, n8143, n8144, n8145, n8147, n8148, n8149, n8150,
    n8152, n8153, n8154, n8155, n8156, n8157, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8168, n8169, n8170, n8171, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8181, n8182, n8184, n8185, n8186, n8187,
    n8188, n8189, n8191, n8192, n8193, n8194, n8196, n8197, n8198, n8199,
    n8202, n8203, n8204, n8205, n8207, n8208, n8209, n8210, n8213, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8224, n8225, n8226,
    n8227, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8237, n8238,
    n8239, n8240, n8242, n8243, n8244, n8245, n8246, n8247, n8249, n8250,
    n8251, n8252, n8253, n8254, n8256, n8257, n8258, n8259, n8260, n8261,
    n8263, n8264, n8265, n8266, n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8284,
    n8285, n8287, n8288, n8289, n8290, n8292, n8293, n8294, n8295, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8306, n8307, n8308,
    n8310, n8311, n8312, n8313, n8314, n8316, n8317, n8318, n8319, n8321,
    n8322, n8324, n8325, n8326, n8327, n8328, n8329, n8331, n8332, n8334,
    n8335, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8410, n8411, n8412, n8414, n8415, n8416, n8417,
    n8418, n8419, n8421, n8422, n8423, n8424, n8425, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8438, n8439, n8440,
    n8441, n8442, n8444, n8445, n8446, n8447, n8448, n8450, n8451, n8453,
    n8454, n8455, n8457, n8458, n8459, n8460, n8462, n8463, n8464, n8465,
    n8466, n8467, n8469, n8470, n8471, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8493, n8494, n8495, n8496, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8506, n8507, n8508, n8509, n8511, n8512,
    n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
    n8524, n8525, n8527, n8529, n8530, n8531, n8533, n8535, n8536, n8537,
    n8538, n8540, n8541, n8542, n8543, n8544, n8545, n8547, n8548, n8549,
    n8550, n8551, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8565, n8566, n8567, n8568, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8581, n8582, n8583,
    n8584, n8587, n8588, n8589, n8590, n8592, n8593, n8594, n8595, n8596,
    n8597, n8599, n8600, n8601, n8602, n8603, n8605, n8606, n8607, n8608,
    n8609, n8610, n8612, n8613, n8615, n8617, n8618, n8619, n8620, n8621,
    n8622, n8623, n8624, n8625, n8626, n8627, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8637, n8638, n8639, n8641, n8642, n8644, n8645,
    n8646, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8656, n8657,
    n8659, n8660, n8661, n8662, n8663, n8664, n8666, n8667, n8668, n8669,
    n8671, n8673, n8674, n8675, n8676, n8677, n8678, n8680, n8681, n8683,
    n8684, n8685, n8686, n8687, n8688, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8699, n8700, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8722, n8723, n8724, n8725, n8726, n8727,
    n8729, n8730, n8731, n8732, n8734, n8735, n8737, n8738, n8739, n8740,
    n8741, n8743, n8744, n8745, n8746, n8747, n8748, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8758, n8759, n8760, n8761, n8762, n8763,
    n8765, n8766, n8767, n8768, n8769, n8770, n8772, n8773, n8774, n8775,
    n8776, n8777, n8779, n8780, n8782, n8783, n8784, n8785, n8786, n8787,
    n8789, n8790, n8791, n8792, n8793, n8794, n8797, n8798, n8800, n8801,
    n8802, n8803, n8804, n8805, n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8823, n8824,
    n8825, n8827, n8828, n8829, n8830, n8831, n8832, n8834, n8835, n8836,
    n8837, n8838, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8852, n8853, n8854, n8855, n8857, n8858, n8859,
    n8860, n8862, n8863, n8865, n8866, n8867, n8868, n8869, n8871, n8872,
    n8873, n8875, n8876, n8877, n8878, n8880, n8881, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8896, n8897,
    n8898, n8899, n8900, n8901, n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8911, n8912, n8913, n8914, n8916, n8917, n8918, n8919, n8921,
    n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8931, n8932,
    n8933, n8934, n8936, n8937, n8938, n8939, n8940, n8941, n8943, n8944,
    n8945, n8946, n8947, n8948, n8950, n8951, n8953, n8954, n8955, n8956,
    n8957, n8958, n8959, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
    n8968, n8969, n8970, n8971, n8972, n8973, n8975, n8976, n8978, n8979,
    n8980, n8981, n8982, n8983, n8985, n8986, n8987, n8988, n8989, n8991,
    n8992, n8993, n8994, n8995, n8997, n8999, n9000, n9001, n9002, n9003,
    n9004, n9006, n9007, n9008, n9009, n9010, n9011, n9013, n9015, n9016,
    n9017, n9018, n9019, n9020, n9022, n9023, n9024, n9025, n9026, n9027,
    n9028, n9029, n9030, n9031, n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9041, n9042, n9044, n9045, n9047, n9048, n9049, n9050, n9051,
    n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
    n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
    n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
    n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
    n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199, n9202, n9203, n9204, n9205,
    n9207, n9208, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9219, n9220, n9222, n9223, n9224, n9225, n9226, n9227, n9229, n9231,
    n9232, n9234, n9235, n9236, n9237, n9238, n9240, n9241, n9242, n9243,
    n9245, n9246, n9247, n9248, n9250, n9251, n9252, n9253, n9255, n9256,
    n9257, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9275, n9276, n9277, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9309, n9310, n9311,
    n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9320, n9321, n9323,
    n9324, n9325, n9326, n9327, n9328, n9330, n9331, n9332, n9334, n9335,
    n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9345, n9346, n9347,
    n9348, n9350, n9351, n9352, n9353, n9355, n9356, n9357, n9358, n9360,
    n9361, n9362, n9363, n9364, n9365, n9367, n9369, n9370, n9371, n9372,
    n9373, n9375, n9376, n9377, n9378, n9379, n9382, n9383, n9384, n9385,
    n9386, n9387, n9389, n9390, n9391, n9392, n9393, n9394, n9396, n9397,
    n9398, n9399, n9400, n9401, n9403, n9404, n9405, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9416, n9417, n9418, n9419, n9420,
    n9421, n9423, n9424, n9426, n9427, n9428, n9429, n9430, n9432, n9433,
    n9434, n9435, n9436, n9437, n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9451, n9452, n9454, n9455, n9456,
    n9457, n9458, n9459, n9461, n9462, n9463, n9464, n9466, n9468, n9469,
    n9470, n9472, n9473, n9474, n9475, n9477, n9478, n9479, n9480, n9481,
    n9483, n9484, n9485, n9487, n9488, n9489, n9491, n9492, n9493, n9494,
    n9497, n9498, n9499, n9500, n9502, n9503, n9505, n9507, n9508, n9509,
    n9510, n9511, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
    n9522, n9523, n9524, n9526, n9527, n9528, n9529, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
    n9544, n9545, n9546, n9547, n9548, n9549, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9567, n9568, n9569, n9571, n9572, n9573, n9574, n9575, n9577, n9578,
    n9579, n9580, n9581, n9583, n9584, n9585, n9586, n9587, n9588, n9590,
    n9591, n9592, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9607, n9608, n9609, n9610, n9611, n9613, n9614,
    n9615, n9616, n9618, n9619, n9620, n9621, n9624, n9625, n9626, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9636, n9637, n9638, n9639,
    n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9648, n9649, n9650,
    n9652, n9654, n9655, n9656, n9658, n9659, n9660, n9661, n9662, n9664,
    n9665, n9666, n9668, n9669, n9671, n9672, n9673, n9674, n9675, n9676,
    n9678, n9679, n9680, n9681, n9683, n9684, n9685, n9686, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9699, n9700,
    n9701, n9702, n9703, n9704, n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9714, n9715, n9717, n9718, n9719, n9720, n9721, n9722, n9724,
    n9725, n9726, n9727, n9728, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9742, n9743, n9744, n9745, n9747,
    n9748, n9749, n9750, n9751, n9752, n9754, n9755, n9756, n9757, n9758,
    n9760, n9761, n9762, n9764, n9765, n9767, n9768, n9769, n9770, n9772,
    n9773, n9774, n9775, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
    n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9798, n9799, n9800, n9801, n9802, n9804, n9805, n9806,
    n9808, n9810, n9811, n9812, n9813, n9814, n9816, n9817, n9818, n9820,
    n9821, n9822, n9823, n9825, n9826, n9827, n9828, n9830, n9831, n9832,
    n9833, n9834, n9835, n9837, n9838, n9839, n9840, n9841, n9843, n9844,
    n9845, n9846, n9847, n9848, n9849, n9851, n9852, n9853, n9854, n9856,
    n9857, n9858, n9859, n9860, n9861, n9863, n9864, n9865, n9866, n9867,
    n9868, n9870, n9871, n9873, n9874, n9875, n9877, n9878, n9879, n9881,
    n9882, n9883, n9884, n9886, n9887, n9888, n9889, n9892, n9893, n9894,
    n9895, n9896, n9897, n9899, n9900, n9901, n9902, n9904, n9905, n9906,
    n9907, n9908, n9909, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9931, n9932, n9934, n9935, n9936, n9937, n9938, n9940,
    n9941, n9942, n9943, n9944, n9945, n9946, n9948, n9949, n9950, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9962, n9963, n9964,
    n9965, n9967, n9968, n9969, n9970, n9971, n9973, n9974, n9975, n9976,
    n9978, n9979, n9980, n9981, n9982, n9983, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9996, n9997, n9999, n10000, n10001,
    n10002, n10003, n10005, n10006, n10007, n10008, n10009, n10010, n10012,
    n10013, n10014, n10015, n10016, n10017, n10019, n10020, n10021, n10022,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10032, n10033,
    n10034, n10035, n10037, n10038, n10039, n10040, n10042, n10043, n10044,
    n10045, n10046, n10047, n10049, n10050, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10060, n10061, n10062, n10064, n10065, n10066,
    n10067, n10068, n10070, n10071, n10072, n10073, n10074, n10075, n10077,
    n10078, n10079, n10080, n10082, n10083, n10085, n10086, n10087, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095, n10097, n10098, n10099,
    n10100, n10102, n10103, n10104, n10106, n10107, n10109, n10110, n10111,
    n10112, n10113, n10114, n10116, n10117, n10118, n10119, n10121, n10123,
    n10124, n10126, n10127, n10128, n10129, n10131, n10132, n10133, n10135,
    n10137, n10138, n10139, n10141, n10142, n10143, n10144, n10145, n10146,
    n10148, n10149, n10150, n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10168, n10169, n10170, n10171, n10172, n10173, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10188, n10189, n10190, n10191, n10192, n10193, n10195, n10196, n10197,
    n10198, n10199, n10200, n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10211, n10212, n10213, n10215, n10216, n10217, n10218, n10219,
    n10220, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10239, n10240,
    n10241, n10243, n10244, n10245, n10246, n10247, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10258, n10259, n10261, n10262,
    n10263, n10264, n10265, n10267, n10268, n10270, n10271, n10272, n10273,
    n10274, n10275, n10277, n10278, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10292, n10293, n10294,
    n10295, n10296, n10297, n10299, n10300, n10301, n10302, n10304, n10305,
    n10306, n10307, n10308, n10309, n10312, n10313, n10314, n10315, n10316,
    n10317, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10327,
    n10328, n10329, n10330, n10332, n10333, n10334, n10335, n10336, n10337,
    n10339, n10340, n10341, n10342, n10344, n10345, n10346, n10347, n10349,
    n10350, n10351, n10352, n10354, n10355, n10356, n10357, n10358, n10359,
    n10361, n10362, n10363, n10364, n10365, n10366, n10368, n10369, n10370,
    n10372, n10373, n10374, n10375, n10376, n10377, n10379, n10380, n10381,
    n10382, n10383, n10384, n10386, n10387, n10389, n10390, n10391, n10392,
    n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10405, n10406, n10407, n10408, n10409, n10411, n10412, n10413,
    n10414, n10416, n10417, n10418, n10419, n10420, n10421, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10431, n10432, n10434, n10435,
    n10436, n10437, n10438, n10439, n10441, n10442, n10444, n10445, n10446,
    n10447, n10448, n10450, n10451, n10452, n10453, n10454, n10456, n10457,
    n10458, n10460, n10461, n10462, n10463, n10464, n10465, n10467, n10468,
    n10469, n10470, n10471, n10472, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10482, n10483, n10484, n10485, n10486, n10487, n10489,
    n10490, n10491, n10492, n10493, n10494, n10496, n10497, n10498, n10499,
    n10500, n10501, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10541, n10542, n10543, n10544, n10545, n10547, n10548,
    n10550, n10551, n10552, n10553, n10555, n10556, n10558, n10559, n10560,
    n10561, n10562, n10564, n10565, n10566, n10567, n10569, n10570, n10571,
    n10573, n10574, n10575, n10576, n10577, n10578, n10580, n10581, n10582,
    n10583, n10584, n10585, n10587, n10588, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10602, n10603,
    n10604, n10605, n10607, n10608, n10609, n10610, n10611, n10612, n10614,
    n10615, n10616, n10617, n10618, n10619, n10621, n10622, n10623, n10624,
    n10626, n10627, n10628, n10629, n10630, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10641, n10642, n10643, n10644, n10645,
    n10646, n10648, n10649, n10650, n10651, n10652, n10653, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10663, n10664, n10666, n10667,
    n10668, n10669, n10670, n10671, n10673, n10674, n10675, n10676, n10677,
    n10678, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10688,
    n10689, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10702, n10703, n10704, n10705, n10706, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10716, n10717, n10718, n10719,
    n10720, n10722, n10723, n10724, n10725, n10726, n10727, n10729, n10731,
    n10732, n10733, n10734, n10736, n10737, n10739, n10740, n10741, n10742,
    n10744, n10745, n10746, n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10757, n10758, n10759, n10760, n10761, n10762, n10764,
    n10765, n10767, n10768, n10769, n10771, n10772, n10773, n10774, n10775,
    n10777, n10778, n10779, n10780, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10790, n10791, n10792, n10793, n10795, n10796, n10798,
    n10799, n10800, n10801, n10802, n10803, n10805, n10806, n10807, n10808,
    n10809, n10810, n10812, n10813, n10814, n10815, n10816, n10818, n10819,
    n10820, n10821, n10822, n10824, n10825, n10827, n10828, n10829, n10830,
    n10832, n10833, n10834, n10835, n10836, n10837, n10839, n10840, n10841,
    n10843, n10844, n10845, n10846, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10859, n10860, n10861, n10862,
    n10863, n10865, n10866, n10867, n10868, n10869, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
    n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
    n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10946, n10947,
    n10948, n10949, n10950, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10982, n10983, n10984, n10985, n10986,
    n10987, n10989, n10990, n10991, n10992, n10993, n10995, n10996, n10998,
    n10999, n11000, n11001, n11002, n11004, n11005, n11006, n11007, n11009,
    n11010, n11011, n11012, n11013, n11015, n11016, n11017, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
    n11040, n11041, n11042, n11043, n11044, n11045, n11047, n11048, n11049,
    n11050, n11051, n11053, n11054, n11055, n11056, n11057, n11058, n11060,
    n11061, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11075, n11076, n11077, n11078, n11080, n11081,
    n11082, n11083, n11084, n11086, n11087, n11088, n11089, n11090, n11091,
    n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11105, n11106, n11108, n11109, n11110, n11111, n11112,
    n11113, n11115, n11116, n11117, n11118, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11128, n11129, n11131, n11132, n11133, n11135,
    n11136, n11137, n11138, n11140, n11141, n11142, n11143, n11145, n11146,
    n11148, n11149, n11150, n11151, n11152, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11162, n11163, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11177, n11179,
    n11180, n11181, n11182, n11184, n11185, n11186, n11187, n11188, n11189,
    n11191, n11192, n11193, n11194, n11195, n11196, n11198, n11199, n11200,
    n11201, n11202, n11203, n11205, n11207, n11208, n11210, n11211, n11212,
    n11213, n11215, n11216, n11217, n11218, n11219, n11221, n11222, n11223,
    n11224, n11225, n11226, n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11237, n11238, n11240, n11241, n11242, n11243, n11244,
    n11245, n11247, n11248, n11249, n11250, n11251, n11252, n11254, n11255,
    n11257, n11258, n11259, n11260, n11261, n11262, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11272, n11273, n11274, n11275, n11276,
    n11277, n11279, n11280, n11281, n11283, n11284, n11285, n11286, n11288,
    n11289, n11290, n11291, n11292, n11293, n11295, n11296, n11297, n11298,
    n11300, n11301, n11302, n11303, n11305, n11306, n11307, n11308, n11309,
    n11311, n11312, n11313, n11314, n11316, n11318, n11319, n11320, n11322,
    n11323, n11324, n11325, n11327, n11328, n11330, n11331, n11332, n11333,
    n11335, n11336, n11339, n11340, n11341, n11342, n11343, n11345, n11346,
    n11347, n11348, n11350, n11351, n11352, n11353, n11354, n11355, n11357,
    n11358, n11359, n11360, n11361, n11363, n11364, n11366, n11367, n11368,
    n11369, n11370, n11372, n11373, n11374, n11375, n11377, n11378, n11379,
    n11380, n11381, n11382, n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11403, n11404, n11405, n11406, n11407, n11408,
    n11410, n11411, n11412, n11413, n11414, n11415, n11417, n11418, n11419,
    n11420, n11422, n11423, n11424, n11425, n11426, n11428, n11429, n11430,
    n11431, n11432, n11433, n11435, n11436, n11437, n11438, n11439, n11440,
    n11442, n11443, n11444, n11445, n11446, n11447, n11449, n11450, n11452,
    n11453, n11454, n11455, n11456, n11458, n11459, n11460, n11461, n11462,
    n11463, n11465, n11466, n11467, n11469, n11470, n11471, n11472, n11474,
    n11475, n11476, n11477, n11478, n11479, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11489, n11491, n11492, n11493, n11494, n11495,
    n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11505, n11506,
    n11508, n11509, n11510, n11511, n11512, n11514, n11515, n11516, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11527, n11528,
    n11529, n11530, n11531, n11533, n11534, n11535, n11536, n11537, n11539,
    n11540, n11541, n11542, n11544, n11545, n11546, n11547, n11548, n11549,
    n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11559, n11560,
    n11561, n11562, n11563, n11564, n11566, n11568, n11569, n11570, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
    n11583, n11584, n11586, n11587, n11588, n11589, n11590, n11591, n11593,
    n11594, n11595, n11596, n11597, n11598, n11600, n11601, n11602, n11603,
    n11604, n11606, n11607, n11608, n11609, n11610, n11611, n11613, n11614,
    n11615, n11616, n11617, n11618, n11620, n11621, n11623, n11624, n11626,
    n11627, n11628, n11629, n11630, n11631, n11633, n11634, n11635, n11637,
    n11638, n11639, n11640, n11641, n11642, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11653, n11654, n11655, n11656, n11658,
    n11659, n11660, n11662, n11663, n11665, n11666, n11667, n11669, n11670,
    n11671, n11672, n11673, n11675, n11676, n11677, n11678, n11679, n11680,
    n11682, n11683, n11684, n11685, n11687, n11688, n11689, n11690, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11705, n11706, n11707, n11708, n11710, n11711, n11712,
    n11714, n11715, n11716, n11717, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11727, n11728, n11729, n11730, n11733, n11734, n11735,
    n11736, n11738, n11739, n11740, n11741, n11742, n11743, n11745, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753, n11755, n11756, n11757,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11775, n11776, n11777, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11791, n11792, n11793, n11794, n11795, n11796, n11798, n11799,
    n11801, n11802, n11803, n11804, n11806, n11807, n11808, n11809, n11810,
    n11811, n11813, n11814, n11815, n11816, n11817, n11819, n11820, n11821,
    n11822, n11824, n11825, n11826, n11827, n11828, n11829, n11831, n11832,
    n11833, n11834, n11835, n11836, n11838, n11839, n11840, n11841, n11842,
    n11843, n11845, n11846, n11848, n11849, n11851, n11852, n11854, n11855,
    n11856, n11858, n11859, n11861, n11863, n11864, n11866, n11867, n11868,
    n11869, n11870, n11871, n11872, n11873, n11874, n11876, n11877, n11879,
    n11880, n11882, n11883, n11884, n11885, n11886, n11888, n11889, n11890,
    n11891, n11893, n11894, n11895, n11896, n11897, n11898, n11900, n11901,
    n11902, n11903, n11905, n11906, n11908, n11909, n11910, n11911, n11912,
    n11913, n11915, n11916, n11917, n11918, n11919, n11921, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11931, n11932, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11944, n11945,
    n11946, n11947, n11948, n11949, n11951, n11952, n11953, n11954, n11955,
    n11956, n11958, n11959, n11960, n11961, n11962, n11964, n11965, n11966,
    n11968, n11969, n11970, n11971, n11972, n11973, n11975, n11976, n11977,
    n11978, n11979, n11981, n11982, n11983, n11985, n11986, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11996, n11997, n11998, n12001,
    n12002, n12003, n12004, n12006, n12007, n12008, n12009, n12010, n12011,
    n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12032, n12033, n12034, n12035, n12036, n12037, n12039, n12040, n12041,
    n12042, n12043, n12045, n12046, n12047, n12048, n12050, n12051, n12053,
    n12054, n12055, n12056, n12058, n12059, n12060, n12061, n12062, n12063,
    n12065, n12066, n12068, n12069, n12070, n12072, n12073, n12074, n12075,
    n12076, n12077, n12078, n12080, n12081, n12082, n12084, n12085, n12086,
    n12087, n12088, n12089, n12091, n12092, n12093, n12094, n12096, n12097,
    n12098, n12099, n12100, n12101, n12103, n12104, n12105, n12106, n12108,
    n12110, n12111, n12113, n12114, n12115, n12116, n12117, n12118, n12120,
    n12121, n12123, n12124, n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12137, n12138, n12139, n12140, n12142,
    n12143, n12145, n12146, n12147, n12148, n12149, n12150, n12152, n12153,
    n12154, n12155, n12157, n12158, n12159, n12160, n12162, n12163, n12164,
    n12166, n12167, n12168, n12169, n12170, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12180, n12181, n12182, n12183, n12184, n12186,
    n12187, n12188, n12189, n12191, n12192, n12194, n12195, n12196, n12197,
    n12198, n12199, n12201, n12202, n12203, n12204, n12205, n12206, n12208,
    n12209, n12210, n12211, n12212, n12213, n12215, n12216, n12217, n12218,
    n12220, n12221, n12223, n12224, n12226, n12227, n12228, n12229, n12231,
    n12232, n12233, n12234, n12235, n12237, n12238, n12240, n12241, n12242,
    n12243, n12245, n12246, n12247, n12248, n12249, n12251, n12252, n12254,
    n12255, n12256, n12257, n12258, n12259, n12261, n12262, n12263, n12264,
    n12266, n12267, n12269, n12270, n12271, n12272, n12274, n12275, n12276,
    n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12287,
    n12288, n12289, n12290, n12291, n12293, n12294, n12295, n12296, n12297,
    n12299, n12300, n12301, n12302, n12303, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12317, n12318,
    n12319, n12320, n12321, n12322, n12324, n12326, n12327, n12328, n12329,
    n12330, n12331, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
    n12341, n12342, n12344, n12345, n12347, n12348, n12349, n12351, n12352,
    n12353, n12354, n12355, n12356, n12358, n12359, n12361, n12362, n12363,
    n12364, n12365, n12367, n12368, n12370, n12371, n12373, n12374, n12375,
    n12376, n12377, n12378, n12380, n12381, n12382, n12383, n12385, n12386,
    n12387, n12389, n12390, n12392, n12393, n12394, n12395, n12397, n12398,
    n12400, n12401, n12402, n12403, n12404, n12405, n12407, n12408, n12410,
    n12412, n12413, n12414, n12415, n12416, n12417, n12419, n12420, n12421,
    n12422, n12423, n12425, n12426, n12427, n12428, n12430, n12431, n12432,
    n12433, n12434, n12435, n12437, n12438, n12439, n12440, n12441, n12442,
    n12444, n12446, n12447, n12448, n12450, n12451, n12452, n12453, n12455,
    n12456, n12458, n12459, n12460, n12461, n12462, n12464, n12465, n12466,
    n12468, n12469, n12470, n12471, n12472, n12474, n12475, n12476, n12477,
    n12478, n12480, n12481, n12482, n12483, n12484, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12494, n12495, n12496, n12497, n688,
    n693, n698_1, n703_1, n708_1, n713_1, n717_1, n722_1, n727_1, n732_1,
    n737_1, n742_1, n747_1, n752_1, n757_1, n762_1, n767_1, n772_1, n777_1,
    n781, n786_1, n791_1, n796_1, n801_1, n806_1, n811_1, n816_1, n821_1,
    n824, n829_1, n834_1, n838_1, n842_1, n847_1, n852_1, n857_1, n862_1,
    n867_1, n872_1, n877_1, n882_1, n887_1, n891_1, n896_1, n901_1, n906_1,
    n911_1, n915_1, n920_1, n925_1, n930, n935_1, n940_1, n945_1, n949_1,
    n954_1, n959_1, n964_1, n969_1, n974_1, n979_1, n984_1, n989_1, n994_1,
    n999_1, n1004_1, n1009_1, n1014_1, n1019_1, n1023_1, n1027_1, n1032_1,
    n1037_1, n1042_1, n1046_1, n1050_1, n1055_1, n1060, n1065_1, n1069_1,
    n1073_1, n1078_1, n1083_1, n1088_1, n1093_1, n1098, n1103, n1108_1,
    n1113_1, n1118_1, n1123, n1128, n1133_1, n1137, n1141_1, n1146_1,
    n1151_1, n1156_1, n1161, n1166_1, n1171, n1175_1, n1178_1, n1182_1,
    n1187_1, n1192_1, n1197_1, n1202, n1206, n1210, n1215_1, n1220_1,
    n1225, n1229_1, n1233_1, n1238_1, n1243_1, n1248_1, n1253_1, n1258_1,
    n1263_1, n1268_1, n1273_1, n1278_1, n1283_1, n1288_1, n1293_1, n1298_1,
    n1303_1, n1308_1, n1313_1, n1318_1, n1323_1, n1328_1, n1332, n1336_1,
    n1340, n1345_1, n1350_1, n1355_1, n1359_1, n1363_1, n1368_1, n1373_1,
    n1378_1, n1383_1, n1388_1, n1393_1, n1398_1, n1403_1, n1408_1, n1412_1,
    n1416_1, n1421_1, n1424, n1429_1, n1434, n1439_1, n1443, n1448, n1453,
    n1458_1, n1463, n1468_1, n1473, n1478_1, n1482, n1486, n1491_1, n1496,
    n1501_1, n1505_1, n1510_1, n1514_1, n1518_1, n1523_1, n1528, n1533_1,
    n1538, n1543_1, n1548_1, n1553, n1558_1, n1563_1, n1568, n1573,
    n1578_1, n1582_1, n1587_1, n1592_1, n1597_1, n1602_1, n1607_1, n1612_1,
    n1617_1, n1622_1, n1627_1, n1632_1, n1637, n1642_1, n1647_1, n1651_1,
    n1655_1, n1660_1, n1665, n1670_1, n1675_1, n1680, n1685_1, n1690_1,
    n1695_1, n1700_1, n1705, n1710_1, n1715_1, n1718_1, n1723, n1728,
    n1733_1, n1738, n1743_1, n1748, n1753_1, n1758_1, n1763_1, n1768_1,
    n1773_1, n1778, n1783_1, n1788_1, n1793_1, n1798_1, n1803, n1808_1,
    n1813_1, n1817, n1822, n1827_1, n1832_1, n1837_1, n1841_1, n1845_1,
    n1850, n1855_1, n1860_1, n1865_1, n1869_1, n1874, n1879_1, n1884_1,
    n1889_1, n1894, n1899, n1904, n1909_1, n1913_1, n1917, n1921_1, n1926,
    n1931_1, n1936_1, n1941_1, n1946, n1951, n1956_1, n1960_1, n1965_1,
    n1970_1, n1975_1, n1980_1, n1984_1, n1989, n1994_1, n1999_1, n2003_1,
    n2008_1, n2013_1, n2018, n2023_1, n2028, n2032, n2036_1, n2041,
    n2046_1, n2051_1, n2056, n2061, n2066, n2071, n2075_1, n2079_1,
    n2084_1, n2088_1, n2093_1, n2097_1, n2102, n2107_1, n2112, n2117_1,
    n2121_1, n2125, n2128_1, n2132, n2137, n2142_1, n2147_1, n2151_1,
    n2155, n2160_1, n2165, n2170_1, n2174, n2179, n2184, n2189, n2194_1,
    n2199, n2204_1, n2209_1, n2213, n2218_1, n2223_1, n2228_1, n2233_1,
    n2238_1, n2243_1, n2248_1, n2253_1, n2258_1, n2262, n2266_1, n2271_1,
    n2276_1, n2281_1, n2286, n2290_1, n2294_1, n2298, n2302_1, n2307,
    n2310_1, n2314, n2319_1, n2324, n2329_1, n2332_1, n2337, n2342_1,
    n2346_1, n2350, n2355_1, n2360, n2365, n2370_1, n2375, n2380_1,
    n2385_1, n2389, n2394_1, n2399_1, n2404_1, n2409_1, n2414_1, n2419_1,
    n2424_1, n2429, n2433_1, n2437_1, n2442, n2446_1, n2450_1, n2455,
    n2459_1, n2464_1, n2469_1, n2474_1, n2479_1, n2484_1, n2489_1, n2494,
    n2499, n2503_1, n2507_1, n2512, n2517_1, n2522_1, n2526_1, n2531,
    n2536_1, n2541_1, n2546_1, n2551_1, n2556, n2561_1, n2566, n2571_1,
    n2576_1, n2581, n2586_1, n2591_1, n2596, n2601_1, n2606_1, n2611_1,
    n2616_1, n2620_1, n2625_1, n2630_1, n2635_1, n2640_1, n2645_1, n2650_1,
    n2655_1, n2660_1, n2664_1, n2669_1, n2673_1, n2678_1, n2683_1, n2688_1,
    n2693_1, n2698_1, n2702_1, n2706_1, n2711_1, n2716_1, n2721_1, n2726_1,
    n2730_1, n2734_1, n2739_1, n2744_1, n2749, n2753_1, n2756_1, n2761_1,
    n2766_1, n2771_1, n2775_1, n2779_1, n2784_1, n2789_1, n2794_1, n2799_1,
    n2804_1, n2809_1, n2814_1, n2819, n2824_1, n2829_1, n2834_1, n2839_1,
    n2844_1, n2849_1, n2853_1, n2858_1, n2863_1, n2868_1, n2873_1, n2877_1,
    n2882_1, n2886_1, n2891_1, n2896, n2900_1, n2905_1, n2910_1, n2915_1,
    n2920_1, n2925_1, n2930_1, n2935_1, n2938_1, n2942_1, n2947_1, n2952_1,
    n2957_1, n2962_1, n2967_1, n2972_1, n2976_1, n2980_1, n2985, n2990_1,
    n2995_1, n3000_1, n3005_1, n3010_1, n3014_1, n3019_1, n3024_1, n3029_1,
    n3034_1, n3039_1, n3043_1, n3048_1, n3053_1, n3058, n3062_1, n3066,
    n3071_1, n3076, n3080_1, n3083_1, n3087, n3092_1, n3097, n3102,
    n3107_1, n3112, n3117, n3122_1, n3127, n3132_1, n3137_1, n3142, n3147,
    n3152_1, n3157_1, n3162, n3166, n3171_1, n3176_1, n3181_1, n3186,
    n3191, n3196, n3201, n3206, n3211_1, n3216, n3220_1, n3224, n3229_1,
    n3233_1, n3238_1, n3243_1, n3248, n3253_1, n3258, n3263_1, n3268,
    n3271, n3276_1, n3280, n3283_1, n3287_1, n3292_1, n3297, n3302_1,
    n3307, n3312, n3317_1, n3322_1, n3327_1, n3332, n3337_1, n3341_1,
    n3346_1, n3351_1, n3356, n3361_1, n3366, n3371_1, n3376, n3380_1,
    n3383_1, n3387, n3392_1, n3397_1, n3402_1, n3407, n3412_1, n3417_1,
    n3422, n3427_1, n3432, n3436_1, n3440_1, n3445, n3450_1, n3455_1,
    n3460, n3465_1, n3469, n3472, n3477_1, n3481_1, n3486, n3491_1, n3496,
    n3501_1, n3506, n3511_1, n3516_1, n3520_1, n3525_1, n3529_1, n3534_1,
    n3539_1, n3544, n3549, n3554_1, n3559, n3562, n3567_1, n3572_1,
    n3577_1, n3582, n3587_1, n3592, n3596, n3600, n3605, n3609_1, n3614,
    n3619_1, n3624_1, n3628_1, n3632, n3637, n3642_1, n3647_1, n3652_1,
    n3657_1, n3662, n3666, n3671, n3676_1, n3681_1, n3686_1, n3691, n3696,
    n3701, n3706_1, n3711, n3716_1, n3721_1, n3726, n3731_1, n3736_1,
    n3741_1, n3746, n3751, n3756, n3761_1, n3766_1, n3771_1, n3776_1,
    n3780_1, n3784_1, n3789_1, n3793_1, n3798_1, n3803_1, n3808, n3813_1,
    n3818_1, n3823_1, n3828_1, n3833_1, n3838_1, n3843_1, n3848, n3852_1,
    n3857, n3862_1, n3867_1, n3872_1, n3877_1, n3882_1, n3887_1, n3892,
    n3897, n3901_1, n3904_1, n3908, n3913, n3918_1, n3923_1, n3928,
    n3933_1, n3938, n3943_1, n3948_1, n3953_1, n3958, n3963_1, n3968,
    n3972, n3976_1, n3981, n3985_1, n3989, n3993_1, n3997_1, n4002, n4007,
    n4011, n4016, n4021_1, n4026, n4031_1, n4036_1, n4040, n4043, n4048_1,
    n4053, n4058_1, n4063_1, n4067_1, n4071_1, n4076_1, n4081, n4085_1,
    n4090, n4095_1, n4100_1, n4105, n4110_1, n4115_1, n4120_1, n4125,
    n4129_1, n4134_1, n4139_1, n4143, n4148, n4152_1, n4157_1, n4161,
    n4165_1, n4170_1, n4175, n4179, n4183_1, n4188, n4193, n4198_1,
    n4203_1, n4207, n4212_1, n4217_1, n4222_1, n4227_1, n4232, n4236_1,
    n4240, n4245_1, n4250, n4255, n4260, n4264, n4268_1, n4273, n4278,
    n4283_1, n4288_1, n4292_1, n4297_1, n4302_1, n4307_1, n4312_1, n4317_1,
    n4322_1, n4327_1, n4332_1, n4337_1, n4341_1, n4345_1, n4350_1, n4355_1,
    n4360_1, n4365_1, n4370, n4375, n4380_1, n4385_1, n4390, n4394_1,
    n4398_1, n4403_1, n4408, n4413, n4418_1, n4423, n4428_1, n4433_1,
    n4438, n4443_1, n4448, n4453, n4457, n4461, n4466, n4471, n4476, n4481,
    n4486_1, n4490_1, n4493, n4496, n4500, n4505, n4510_1, n4515_1, n4520,
    n4525, n4530_1, n4535_1, n4540_1, n4545, n4550_1, n4555, n4560, n4565,
    n4570_1, n4575, n4579, n4583, n4588_1, n4593_1, n4598, n4603, n4608,
    n4613, n4618, n4623, n4628, n4632_1, n4637_1, n4641_1, n4645, n4649,
    n4653_1, n4658, n4663_1, n4668, n4673_1, n4678, n4683, n4688, n4693,
    n4698, n4703_1, n4708, n4713_1, n4718, n4723_1, n4728, n4732, n4737_1,
    n4742_1, n4747_1, n4752_1, n4757_1, n4762, n4767_1, n4771_1, n4774_1,
    n4778_1, n4783_1, n4788, n4793_1, n4798, n4803, n4808_1, n4813_1,
    n4818_1, n4823_1, n4828, n4833_1, n4838_1, n4843, n4847, n4852_1,
    n4856_1, n4860_1, n4865, n4869, n4874, n4878_1, n4883_1, n4888_1,
    n4891, n4895_1, n4900_1, n4905, n4910_1, n4915_1, n4920, n4925,
    n4930_1, n4935_1, n4940_1, n4945_1, n4949_1, n4954_1, n4959_1, n4964_1,
    n4969_1, n4974, n4979, n4984_1, n4988, n4993, n4998_1, n5003, n5008,
    n5012_1, n5017, n5022, n5027, n5032, n5037, n5042, n5047_1, n5052_1,
    n5057_1, n5061, n5065, n5070_1, n5075_1, n5080, n5084_1, n5089_1,
    n5094_1, n5099, n5104, n5108, n5112, n5117, n5122_1, n5127, n5132_1,
    n5137_1, n5142_1, n5147_1, n5152_1, n5157, n5161, n5166, n5171,
    n5176_1, n5181_1, n5186_1, n5191, n5196_1, n5201_1, n5206_1, n5211_1,
    n5215_1, n5219_1, n5224_1, n5229_1, n5234_1, n5238_1, n5242_1, n5247_1,
    n5252_1, n5257_1, n5262_1, n5266_1, n5270, n5274_1, n5279, n5284_1,
    n5289, n5294, n5299_1, n5304_1, n5309_1, n5314, n5319_1, n5323_1,
    n5327_1, n5332_1, n5336_1, n5340_1, n5345_1, n5350_1, n5354_1, n5357_1,
    n5362_1, n5367_1, n5372_1, n5377_1, n5382_1, n5386_1, n5390_1, n5394_1,
    n5399_1, n5403_1, n5407_1, n5412, n5417_1, n5422_1, n5427_1, n5432,
    n5437_1, n5442_1, n5447, n5452_1, n5457, n5462_1, n5467_1, n5472_1,
    n5477_1, n5482_1, n5487_1, n5492_1, n5497_1, n5502_1, n5507_1, n5512_1,
    n5517_1, n5522_1, n5527_1, n5532_1, n5537_1, n5542, n5546_1, n5550_1,
    n5555_1, n5559_1, n5564_1, n5569_1, n5574, n5579_1, n5584_1, n5589_1,
    n5594, n5599_1, n5604_1, n5609_1, n5614_1, n5619_1, n5624, n5629,
    n5634_1, n5639, n5644_1, n5649_1, n5654_1, n5659, n5663_1, n5667,
    n5672, n5677_1, n5682_1, n5687_1, n5691, n5696, n5701_1, n5706_1,
    n5711, n5715_1, n5719_1, n5724_1, n5729, n5734_1, n5739, n5744_1,
    n5749_1, n5754_1, n5759, n5764, n5769, n5773, n5777_1, n5782, n5787,
    n5792, n5797, n5802, n5807, n5812_1, n5817_1, n5822, n5826, n5829_1,
    n5834, n5839, n5843_1, n5847_1, n5851, n5856, n5860_1, n5865_1,
    n5870_1, n5875_1, n5880_1, n5885_1, n5889, n5894_1, n5899, n5904,
    n5909, n5914, n5919_1, n5924_1, n5929, n5934, n5938_1, n5942, n5947_1,
    n5952_1, n5957_1, n5962_1, n5967, n5972, n5976, n5981, n5986_1, n5991,
    n5995_1, n5999_1, n6004_1, n6009, n6013_1, n6018, n6023_1, n6028,
    n6033_1, n6038, n6043_1, n6048_1, n6053, n6057_1, n6062_1, n6067,
    n6072_1, n6077_1, n6082_1, n6087, n6092_1, n6097_1, n6101, n6105_1,
    n6110, n6115_1, n6120_1, n6124_1, n6128_1, n6133_1, n6138, n6143,
    n6148, n6153, n6157, n6161, n6166, n6170, n6175, n6180, n6184, n6189,
    n6193, n6197, n6202, n6207_1, n6212, n6217, n6222, n6227, n6231, n6236,
    n6241, n6246, n6251_1, n6256_1, n6261_1, n6266, n6271, n6276, n6280,
    n6285, n6290_1, n6294, n6298, n6303, n6307, n6311, n6316, n6321, n6326,
    n6331, n6336, n6341_1, n6345, n6350, n6355, n6360, n6365, n6370, n6374,
    n6377, n6381, n6386_1, n6391, n6396, n6400, n6404, n6409, n6414, n6418,
    n6423, n6428, n6433, n6438, n6443, n6448, n6453, n6458, n6463, n6468,
    n6473, n6478, n6483, n6488, n6493, n6498, n6503, n6508, n6513, n6518,
    n6523, n6527, n6532, n6537, n6542, n6547, n6552, n6556, n6561, n6566,
    n6571, n6576, n6581, n6586, n6591, n6596, n6601, n6606, n6611, n6616,
    n6621, n6625, n6630, n6635, n6639, n6643, n6647, n6652, n6657, n6662,
    n6666, n6671, n6676, n6681;
  assign n4125_1 = ~Pg56 & Pg54;
  assign n4126 = ~Ng55 & n4125_1;
  assign n4127 = ~Pg57 & n4126;
  assign n3828_1 = ~Pg53 & n4127;
  assign n4129 = ~Ng46 & ~Ng8;
  assign n4130 = ~Ng45 & n4129;
  assign n4131 = Ng51 & n4130;
  assign n4132 = ~Ng52 & n4131;
  assign n4133 = ~Ng48 & n4132;
  assign n4134 = ~Ng16 & ~Ng50;
  assign n4135 = n4133 & n4134;
  assign n4136 = Ng794 & n4135;
  assign n4137 = Ng16 & ~Ng50;
  assign n4138 = Ng52 & n4130;
  assign n4139 = ~Ng48 & n4138;
  assign n4140 = Ng51 & n4139;
  assign n4141 = n4137 & n4140;
  assign n4142 = Ng37 & n4141;
  assign n4143_1 = ~Ng52 & Ng46;
  assign n4144 = Ng48 & Ng45;
  assign n4145 = Ng8 & n4144;
  assign n4146 = n4143_1 & n4145;
  assign n4147 = ~Ng51 & n4146;
  assign n4148_1 = n4134 & n4147;
  assign n4149 = Ng2955 & n4148_1;
  assign n4150 = ~Ng16 & Ng50;
  assign n4151 = n4139 & n4150;
  assign n4152 = ~Ng51 & n4151;
  assign n4153 = Ng586 & n4152;
  assign n4154 = ~n4149 & ~n4153;
  assign n4155 = ~n4142 & n4154;
  assign n4156 = ~Ng51 & n4130;
  assign n4157 = ~Ng52 & n4156;
  assign n4158 = ~Ng48 & n4157;
  assign n4159 = n4134 & n4158;
  assign n4160 = Ng534 & n4159;
  assign n4161_1 = n4150 & n4158;
  assign n4162 = Ng613 & n4161_1;
  assign n4163 = ~n4160 & ~n4162;
  assign n4164 = n4133 & n4137;
  assign n4165 = Ng2868 & n4164;
  assign n4166 = Ng51 & n4146;
  assign n4167 = n4150 & n4166;
  assign n4168 = Ng48 & n4134;
  assign n4169 = n4132 & n4168;
  assign n4170 = Ng2882 & n4169;
  assign n4171 = ~n4167 & ~n4170;
  assign n4172 = ~n4165 & n4171;
  assign n4173 = n4163 & n4172;
  assign n4174 = n4155 & n4173;
  assign n4175_1 = n4134 & n4140;
  assign n4176 = ~n4152 & ~n4161_1;
  assign n4177 = ~n4175_1 & n4176;
  assign n4178 = ~n4135 & n4177;
  assign n4179_1 = ~Pg35 & ~n4178;
  assign n4180 = n4134 & n4166;
  assign n4181 = Ng2950 & n4180;
  assign n4182 = Ng758 & n4175_1;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = ~n4179_1 & n4183;
  assign n4185 = n4174 & n4184;
  assign n4186 = ~n4136 & n4185;
  assign n4187 = n3828_1 & ~n4186;
  assign n4188_1 = n3828_1 & n4150;
  assign n4189 = Ng48 & n4188_1;
  assign n4190 = n4132 & n4189;
  assign n4191 = Ng4300 & n4190;
  assign n4192 = n4157 & n4168;
  assign n4193_1 = n3828_1 & n4192;
  assign n4194 = Ng4172 & n4193_1;
  assign n4195 = ~n4191 & ~n4194;
  assign n4196 = Ng16 & n3828_1;
  assign n4197 = Ng50 & n4196;
  assign n4198 = n4133 & n4197;
  assign n4199 = ~Ng4927 & n4198;
  assign n4200 = ~Pg53 & ~n4127;
  assign n4201 = Ng16 & n4200;
  assign n4202 = ~n4199 & ~n4201;
  assign n4203 = n3828_1 & n4137;
  assign n4204 = n4158 & n4203;
  assign n4205 = Ng1291 & n4204;
  assign n4206 = n4202 & ~n4205;
  assign n4207_1 = n4195 & n4206;
  assign n4208 = n4133 & n4188_1;
  assign n4209 = Ng947 & n4208;
  assign n4210 = n4158 & n4197;
  assign n4211 = ~Ng4737 & n4210;
  assign n4212 = ~n4209 & ~n4211;
  assign n4213 = n4207_1 & n4212;
  assign n2238_1 = n4187 | ~n4213;
  assign n4215 = Ng749 & n4175_1;
  assign n4216 = Ng608 & n4161_1;
  assign n4217 = ~Ng550 & n4159;
  assign n4218 = ~n4216 & ~n4217;
  assign n4219 = Ng2960 & n4180;
  assign n4220 = n4218 & ~n4219;
  assign n4221 = \[4433]  & n4141;
  assign n4222 = Ng790 & n4135;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = Ng2873 & n4164;
  assign n4225 = Ng572 & n4152;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = n4223 & n4226;
  assign n4228 = n4220 & n4227;
  assign n4229 = Ng2965 & n4148_1;
  assign n4230 = Ng2878 & n4169;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232_1 = ~n4179_1 & n4231;
  assign n4233 = n4228 & n4232_1;
  assign n4234 = ~n4215 & n4233;
  assign n4235 = n3828_1 & ~n4234;
  assign n4236 = Ng4253 & n4190;
  assign n4237 = ~Ng1296 & n4204;
  assign n4238 = n4157 & n4189;
  assign n4239 = Ng2130 & n4238;
  assign n4240_1 = ~n4237 & ~n4239;
  assign n4241 = Ng50 & n4200;
  assign n4242 = ~Ng952 & n4208;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = Ng4176 & n4193_1;
  assign n4245 = Ng52 & n4156;
  assign n4246 = n4189 & n4245;
  assign n4247 = Ng2689 & n4246;
  assign n4248 = ~n4244 & ~n4247;
  assign n4249 = n4243 & n4248;
  assign n4250_1 = n4240_1 & n4249;
  assign n4251 = ~n4236 & n4250_1;
  assign n4940_1 = n4235 | ~n4251;
  assign n4253 = n2238_1 & ~n4940_1;
  assign n4254 = ~n2238_1 & n4940_1;
  assign n4255_1 = ~n4253 & ~n4254;
  assign n4256 = Ng807 & n4135;
  assign n4257 = Ng2898 & n4169;
  assign n4258 = Ng763 & n4175_1;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260_1 = ~n4256 & n4259;
  assign n4261 = Ng542 & n4159;
  assign n4262 = Ng617 & n4161_1;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264_1 = Ng577 & n4152;
  assign n4265 = ~n4167 & ~n4264_1;
  assign n4266 = n4263 & n4265;
  assign n4267 = n4260_1 & n4266;
  assign n4268 = Ng2894 & n4192;
  assign n4269 = Ng2936 & n4180;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = Ng2941 & n4148_1;
  assign n4272 = Ng2988 & n4164;
  assign n4273_1 = ~n4271 & ~n4272;
  assign n4274 = n4270 & n4273_1;
  assign n4275 = n4267 & n4274;
  assign n4276 = ~n4179_1 & n4275;
  assign n4277 = n3828_1 & ~n4276;
  assign n4278_1 = Ng48 & n4200;
  assign n4279 = Ng4912 & n4198;
  assign n4280 = Ng5160 & n4238;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = ~n4278_1 & n4281;
  assign n4283 = Ng1135 & ~Ng947;
  assign n4284 = n4208 & n4283;
  assign n4285 = Ng4722 & n4210;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = Ng1478 & ~Ng1291;
  assign n4288 = n4204 & n4287;
  assign n4289 = Ng6545 & n4246;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n4286 & n4290;
  assign n4292 = n4282 & n4291;
  assign n1350_1 = n4277 | ~n4292;
  assign n4294 = Ng1129 & ~Ng947;
  assign n4295 = n4208 & n4294;
  assign n4296 = Ng4922 & n4198;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = Ng3502 & n4246;
  assign n4299 = Ng46 & n4200;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = n4297 & n4300;
  assign n4302 = Ng2999 & n4164;
  assign n4303 = Ng2852 & n4192;
  assign n4304 = Ng2917 & n4148_1;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = Ng590 & n4152;
  assign n4307 = n4305 & ~n4306;
  assign n4308 = Ng626 & n4161_1;
  assign n4309 = Ng2856 & n4169;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = n4307 & n4310;
  assign n4312 = ~Pg35 & ~n4177;
  assign n4313 = Ng772 & n4175_1;
  assign n4314 = Ng2912 & n4180;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = ~n4312 & n4315;
  assign n4317 = n4311 & n4316;
  assign n4318 = ~n4302 & n4317;
  assign n4319 = n3828_1 & ~n4318;
  assign n4320 = Ng5853 & n4238;
  assign n4321 = Ng4732 & n4210;
  assign n4322 = Ng1472 & ~Ng1291;
  assign n4323 = n4204 & n4322;
  assign n4324 = ~n4321 & ~n4323;
  assign n4325 = ~n4320 & n4324;
  assign n4326 = ~n4319 & n4325;
  assign n2739_1 = ~n4301 | ~n4326;
  assign n4328 = ~n1350_1 & ~n2739_1;
  assign n4329 = n1350_1 & n2739_1;
  assign n4330 = ~n4328 & ~n4329;
  assign n4331 = n4255_1 & n4330;
  assign n4332 = ~n4255_1 & ~n4330;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = Ng55 & ~n4125_1;
  assign n4335 = Ng604 & n4161_1;
  assign n4336 = \[4426]  & n4159;
  assign n4337 = ~n4335 & ~n4336;
  assign n4338 = Pg127 & n4164;
  assign n4339 = Pg92 & n4141;
  assign n4340 = Ng2970 & n4180;
  assign n4341 = Ng2886 & n4169;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~n4339 & n4342;
  assign n4344 = ~n4338 & n4343;
  assign n4345 = Ng2975 & n4148_1;
  assign n4346 = Ng744 & n4175_1;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = n4137 & n4147;
  assign n4349 = Ng2980 & n4348;
  assign n4350 = n4347 & ~n4349;
  assign n4351 = n4344 & n4350;
  assign n4352 = Ng785 & n4135;
  assign n4353 = Ng568 & n4152;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4179_1 & n4354;
  assign n4356 = n4351 & n4355;
  assign n4357 = n4337 & n4356;
  assign n4358 = n3828_1 & ~n4357;
  assign n4359 = Ng1283 & n4204;
  assign n4360 = Ng2697 & n4246;
  assign n4361 = Ng51 & n4200;
  assign n4362 = Ng939 & n4208;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = ~n4360 & n4363;
  assign n4365 = Ng2138 & n4238;
  assign n4366 = Ng4146 & n4193_1;
  assign n4367 = Ng4249 & n4190;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = ~n4365 & n4368;
  assign n4370_1 = n4364 & n4369;
  assign n4371 = ~n4359 & n4370_1;
  assign n2512 = n4358 | ~n4371;
  assign n4373 = n4334 & ~n2512;
  assign n4374 = ~n4334 & n2512;
  assign n4375_1 = ~n4373 & ~n4374;
  assign n4376 = Ng2890 & n4164;
  assign n4377 = Ng562 & n4152;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = Ng599 & n4161_1;
  assign n4380 = Ng2984 & n4348;
  assign n4381 = ~n4167 & ~n4380;
  assign n4382 = ~n4379 & n4381;
  assign n4383 = n4378 & n4382;
  assign n4384 = Pg100 & n4141;
  assign n4385 = Ng739 & n4175_1;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = Ng199 & n4159;
  assign n4388 = Ng781 & n4135;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390_1 = n4386 & n4389;
  assign n4391 = n4383 & n4390_1;
  assign n4392 = ~n4179_1 & n4391;
  assign n4393 = n3828_1 & ~n4392;
  assign n4394 = Ng2704 & n4246;
  assign n4395 = Ng2145 & n4238;
  assign n4396 = ~n4394 & ~n4395;
  assign n4397 = ~n4393 & n4396;
  assign n4398 = Ng52 & n4200;
  assign n4399 = Ng4245 & n4190;
  assign n4400 = Ng1287 & n4204;
  assign n4401 = Ng943 & n4208;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = ~n4399 & n4402;
  assign n4404 = ~n4398 & n4403;
  assign n4405 = Ng4157 & n4193_1;
  assign n4406 = n4404 & ~n4405;
  assign n1587_1 = ~n4397 | ~n4406;
  assign n4408_1 = ~Ng2994 & n4164;
  assign n4409 = Ng2922 & n4180;
  assign n4410 = ~n4408_1 & ~n4409;
  assign n4411 = Ng582 & n4152;
  assign n4412 = n4410 & ~n4411;
  assign n4413_1 = Ng2864 & n4169;
  assign n4414 = Ng767 & n4175_1;
  assign n4415 = Ng2860 & n4192;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n4413_1 & n4416;
  assign n4418 = n4412 & n4417;
  assign n4419 = Ng622 & n4161_1;
  assign n4420 = Ng546 & n4159;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = Ng554 & n4135;
  assign n4423_1 = Ng2927 & n4148_1;
  assign n4424 = ~n4422 & ~n4423_1;
  assign n4425 = n4421 & n4424;
  assign n4426 = n4418 & n4425;
  assign n4427 = ~n4179_1 & n4426;
  assign n4428 = n3828_1 & ~n4427;
  assign n4429 = Ng4907 & n4198;
  assign n4430 = Ng8 & n4200;
  assign n4431 = Ng1105 & ~Ng947;
  assign n4432 = n4208 & n4431;
  assign n4433 = ~n4430 & ~n4432;
  assign n4434 = ~n4429 & n4433;
  assign n4435 = Ng5507 & n4238;
  assign n4436 = Ng3151 & n4246;
  assign n4437 = Ng4717 & n4210;
  assign n4438_1 = ~n4436 & ~n4437;
  assign n4439 = Ng1448 & ~Ng1291;
  assign n4440 = n4204 & n4439;
  assign n4441 = n4438_1 & ~n4440;
  assign n4442 = ~n4435 & n4441;
  assign n4443 = n4434 & n4442;
  assign n3892 = n4428 | ~n4443;
  assign n4445 = Ng538 & n4159;
  assign n4446 = Ng632 & n4161_1;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448_1 = Ng2907 & n4180;
  assign n4449 = n4447 & ~n4448_1;
  assign n4450 = Ng595 & n4152;
  assign n4451 = Ng776 & n4175_1;
  assign n4452 = Ng2902 & n4148_1;
  assign n4453_1 = ~n4451 & ~n4452;
  assign n4454 = Ng2848 & n4169;
  assign n4455 = n4453_1 & ~n4454;
  assign n4456 = ~n4450 & n4455;
  assign n4457_1 = Ng2844 & n4192;
  assign n4458 = ~n4312 & ~n4457_1;
  assign n4459 = n4456 & n4458;
  assign n4460 = n4449 & n4459;
  assign n4461_1 = n3828_1 & ~n4460;
  assign n4462 = Ng6199 & n4238;
  assign n4463 = ~Ng1291 & Ng1300;
  assign n4464 = n4204 & n4463;
  assign n4465 = Ng4727 & n4210;
  assign n4466_1 = ~n4464 & ~n4465;
  assign n4467 = Ng4917 & n4198;
  assign n4468 = Ng956 & ~Ng947;
  assign n4469 = n4208 & n4468;
  assign n4470 = Ng45 & n4200;
  assign n4471_1 = ~n4469 & ~n4470;
  assign n4472 = ~n4467 & n4471_1;
  assign n4473 = Ng3853 & n4246;
  assign n4474 = n4472 & ~n4473;
  assign n4475 = n4466_1 & n4474;
  assign n4476_1 = ~n4462 & n4475;
  assign n2891_1 = n4461_1 | ~n4476_1;
  assign n4478 = n3892 & ~n2891_1;
  assign n4479 = ~n3892 & n2891_1;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481_1 = ~n1587_1 & n4480;
  assign n4482 = n1587_1 & ~n4480;
  assign n4483 = ~n4481_1 & ~n4482;
  assign n4484 = n4375_1 & ~n4483;
  assign n4485 = ~n4375_1 & n4483;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = ~n4333 & ~n4486;
  assign n4488 = n4333 & n4486;
  assign n3297 = ~n4487 & ~n4488;
  assign Pg34972 = ~Ng22 | n3297;
  assign n4491 = ~Pg72 & ~Ng4322;
  assign n4492 = Pg72 & Ng4322;
  assign n4493_1 = ~n4491 & ~n4492;
  assign n4494 = ~Pg73 & Ng4332;
  assign n4495 = Pg73 & ~Ng4332;
  assign n4496_1 = ~n4494 & ~n4495;
  assign n4497 = ~n4493_1 & n4496_1;
  assign n4498 = ~Ng4311 & n4497;
  assign n4499 = ~Ng4366 & n4498;
  assign Pg34956 = Ng4369 & ~n4499;
  assign Pg34927 = ~Ng22 | n2512;
  assign Pg34925 = ~Ng22 | n4940_1;
  assign Pg34923 = ~Ng22 | n2238_1;
  assign Pg34921 = ~Ng22 | n1350_1;
  assign Pg34919 = ~Ng22 | n3892;
  assign Pg34917 = ~Ng22 | n2739_1;
  assign Pg34915 = ~Ng22 | n1587_1;
  assign Pg34913 = ~Ng22 | n2891_1;
  assign n4509 = ~Pg72 & ~Ng482;
  assign n4510 = Pg72 & Ng482;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~Pg73 & Ng490;
  assign n4513 = Pg73 & ~Ng490;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4511 & n4514;
  assign n4516 = Ng479 & ~Ng528;
  assign n4517 = n4515 & n4516;
  assign Pg34788 = Ng890 & ~n4517;
  assign Pg34437 = ~Pg113 | ~Ng2868;
  assign Pg34436 = ~Pg113 | ~Ng2873;
  assign n4521 = ~Ng4082 & ~Ng4141;
  assign n4522 = ~Ng4098 & ~Ng4093;
  assign n4523 = ~Ng4087 & n4522;
  assign n4524 = Ng4076 & Ng4112;
  assign n4525_1 = n4523 & n4524;
  assign n4526 = n4521 & ~n4525_1;
  assign n4527 = ~Ng4064 & ~Ng4057;
  assign n4528 = ~n4526 & n4527;
  assign Pg34435 = ~Ng4125 & n4528;
  assign n4530 = Ng4311 & n4497;
  assign n4531 = Ng4349 & ~Ng4358;
  assign n4532 = Ng3288 & Ng3352;
  assign n4533 = n4531 & n4532;
  assign n4534 = Ng4349 & Ng4358;
  assign n4535 = Ng4054 & Ng3990;
  assign n4536 = n4534 & n4535;
  assign n4537 = ~Ng4349 & ~Ng4358;
  assign n4538 = Ng6682 & Ng6741;
  assign n4539 = n4537 & n4538;
  assign n4540 = ~Ng4349 & Ng4358;
  assign n4541 = Ng3639 & Ng3703;
  assign n4542 = n4540 & n4541;
  assign n4543 = ~n4539 & ~n4542;
  assign n4544 = ~n4536 & n4543;
  assign n4545_1 = ~n4533 & n4544;
  assign n4546 = n4530 & ~n4545_1;
  assign n4547 = Ng6336 & Ng6395;
  assign n4548 = n4534 & n4547;
  assign n4549 = Ng5703 & Ng5644;
  assign n4550 = n4531 & n4549;
  assign n4551 = Ng5990 & Ng6049;
  assign n4552 = n4540 & n4551;
  assign Pg31860 = Ng5297 & Ng5357;
  assign n4554 = n4537 & Pg31860;
  assign n4555_1 = ~n4552 & ~n4554;
  assign n4556 = ~n4550 & n4555_1;
  assign n4557 = ~n4548 & n4556;
  assign n4558 = n4498 & ~n4557;
  assign n3803_1 = n4546 | n4558;
  assign n4560_1 = Pg99 & Ng37;
  assign n4561 = ~Pg134 & ~n4560_1;
  assign n4562 = Pg113 & ~n4561;
  assign n4563 = n4497 & n4562;
  assign Pg34425 = n3803_1 | ~n4563;
  assign n4565_1 = Ng518 & n4515;
  assign n4566 = Ng528 & n4565_1;
  assign n4567 = ~Ng504 & n4566;
  assign n4568 = ~Ng2599 & Ng2629;
  assign n4569 = n4567 & n4568;
  assign n4570 = Ng504 & n4566;
  assign n4571 = ~Ng2465 & Ng2495;
  assign n4572 = n4570 & n4571;
  assign n4573 = ~Ng518 & n4515;
  assign n4574 = ~Ng528 & ~Ng504;
  assign n4575_1 = n4573 & n4574;
  assign Pg31862 = Ng1668 & ~Ng1636;
  assign n4577 = n4575_1 & Pg31862;
  assign n4578 = ~Ng528 & Ng504;
  assign n4579_1 = n4565_1 & n4578;
  assign n4580 = Ng1936 & ~Ng1906;
  assign n4581 = n4579_1 & n4580;
  assign n4582 = ~n4577 & ~n4581;
  assign n4583_1 = ~n4572 & n4582;
  assign n4584 = ~n4569 & n4583_1;
  assign n4585 = Ng528 & n4573;
  assign n4586 = Ng504 & n4585;
  assign n4587 = ~Ng2331 & Ng2361;
  assign n4588 = n4586 & n4587;
  assign n4589 = ~Ng504 & n4585;
  assign n4590 = Ng2227 & ~Ng2197;
  assign n4591 = n4589 & n4590;
  assign n4592 = n4573 & n4578;
  assign n4593 = Ng1802 & ~Ng1772;
  assign n4594 = n4592 & n4593;
  assign n4595 = n4565_1 & n4574;
  assign n4596 = ~Ng2040 & Ng2070;
  assign n4597 = n4595 & n4596;
  assign n4598_1 = ~n4594 & ~n4597;
  assign n4599 = ~n4591 & n4598_1;
  assign n4600 = ~n4588 & n4599;
  assign n5649_1 = ~n4584 | ~n4600;
  assign n4602 = n4515 & ~n5649_1;
  assign Pg34383 = ~n4562 | ~n4602;
  assign n4604 = Ng4878 & Ng4843;
  assign n4605 = Ng4849 & Ng4859;
  assign n4606 = n4604 & n4605;
  assign n4607 = Ng4899 & Ng4975;
  assign n4608_1 = Ng4983 & Ng4966;
  assign n4609 = ~Ng4991 & n4608_1;
  assign n4610 = n4607 & n4609;
  assign n4611 = n4606 & n4610;
  assign n4612 = n4530 & n4611;
  assign n4613_1 = Ng4709 & Ng4785;
  assign n4614 = Ng4776 & ~Ng4801;
  assign n4615 = Ng4793 & n4614;
  assign n4616 = n4613_1 & n4615;
  assign n4617 = Ng4653 & Ng4688;
  assign n4618_1 = Ng4659 & n4617;
  assign n4619 = Ng4669 & n4618_1;
  assign n4620 = n4498 & n4619;
  assign n4621 = n4616 & n4620;
  assign n4036_1 = n4612 | n4621;
  assign Pg34221 = ~n4563 | n4036_1;
  assign n4624 = ~Pg72 & ~Ng2759;
  assign n4625 = Pg72 & Ng2759;
  assign n4626 = ~n4624 & ~n4625;
  assign n4627 = ~Pg73 & Ng2763;
  assign n4628_1 = Pg73 & ~Ng2763;
  assign n4629 = ~n4627 & ~n4628_1;
  assign n4630 = ~n4626 & n4629;
  assign n4631 = Ng2756 & Ng2748;
  assign n4632 = Ng2741 & n4631;
  assign n4633 = n4630 & n4632;
  assign n4634 = Ng2610 & ~Ng2619;
  assign n4635 = n4633 & n4634;
  assign n4636 = Ng2748 & n4630;
  assign n4637 = Ng2741 & n4636;
  assign n4638 = ~Ng2756 & n4637;
  assign n4639 = Ng2051 & ~Ng2060;
  assign n4640 = n4638 & n4639;
  assign n4641 = ~n4635 & ~n4640;
  assign n4642 = Ng2756 & n4630;
  assign n4643 = ~Ng2748 & n4642;
  assign n4644 = ~Ng2741 & n4643;
  assign n4645_1 = Ng2208 & ~Ng2217;
  assign n4646 = n4644 & n4645_1;
  assign n4647 = ~Ng2741 & n4636;
  assign n4648 = Ng2756 & n4647;
  assign n4649_1 = ~Ng2485 & Ng2476;
  assign n4650 = n4648 & n4649_1;
  assign n4651 = ~n4646 & ~n4650;
  assign n4652 = n4641 & n4651;
  assign n4653 = ~Ng2756 & n4647;
  assign n4654 = ~Ng1926 & Ng1917;
  assign n4655 = n4653 & n4654;
  assign n4656 = ~Ng2756 & ~Ng2748;
  assign n4657 = Ng2741 & n4656;
  assign n4658_1 = n4630 & n4657;
  assign n4659 = Ng1783 & ~Ng1792;
  assign n4660 = n4658_1 & n4659;
  assign n4661 = ~n4655 & ~n4660;
  assign n4662 = ~Ng2741 & n4656;
  assign n4663 = n4630 & n4662;
  assign Pg31863 = ~Ng1657 & Ng1648;
  assign n4665 = n4663 & Pg31863;
  assign n4666 = Ng2741 & n4643;
  assign n4667 = Ng2342 & ~Ng2351;
  assign n4668_1 = n4666 & n4667;
  assign n4669 = ~n4665 & ~n4668_1;
  assign n4670 = n4661 & n4669;
  assign n2342_1 = ~n4652 | ~n4670;
  assign n4672 = n4562 & ~n2342_1;
  assign Pg34201 = ~n4630 | ~n4672;
  assign n4674 = ~Ng4793 & n4614;
  assign n4675 = Ng4669 & Ng4659;
  assign n4676 = Ng4653 & n4675;
  assign n4677 = n4674 & n4676;
  assign n4678_1 = ~Ng4709 & ~Ng4785;
  assign n4679 = Ng4698 & n4678_1;
  assign n4680 = n4677 & n4679;
  assign Pg33959 = Ng4646 & ~n4680;
  assign n4682 = Ng4955 & n4607;
  assign n4683_1 = ~Ng4899 & ~Ng4975;
  assign n4684 = Ng4888 & n4683_1;
  assign n4685 = ~n4682 & ~n4684;
  assign n4686 = Ng4899 & ~Ng4975;
  assign n4687 = Ng4944 & n4686;
  assign n4688_1 = ~Ng4899 & Ng4975;
  assign n4689 = Ng4933 & n4688_1;
  assign n4690 = ~n4687 & ~n4689;
  assign n6676 = ~n4685 | ~n4690;
  assign n4692 = \[4658]  & ~n4561;
  assign n4693_1 = \[4651]  & n4692;
  assign Pg33935 = n6676 | ~n4693_1;
  assign n4695 = Ng4507 & ~n4561;
  assign Pg33874 = \[4507]  | ~n4695;
  assign n4697 = ~Pg72 & ~Ng4108;
  assign n4698_1 = Pg72 & Ng4108;
  assign n4699 = ~n4697 & ~n4698_1;
  assign n4700 = ~Pg73 & Ng4104;
  assign n4701 = Pg73 & ~Ng4104;
  assign n4702 = ~n4700 & ~n4701;
  assign n4703 = ~n4699 & n4702;
  assign n4704 = Ng4098 & Ng4093;
  assign n4705 = Ng3530 & Ng3522;
  assign n4706 = Ng3518 & n4705;
  assign n4707 = n4704 & n4706;
  assign n4708_1 = Ng5180 & Ng5188;
  assign Pg32975 = Ng5176 & n4708_1;
  assign n4710 = n4522 & Pg32975;
  assign n4711 = ~n4707 & ~n4710;
  assign n4712 = Ng4098 & ~Ng4093;
  assign n4713 = Ng6573 & Ng6565;
  assign n4714 = Ng6561 & n4713;
  assign n4715 = n4712 & n4714;
  assign n4716 = ~Ng4098 & Ng4093;
  assign n4717 = Ng5873 & Ng5881;
  assign n4718_1 = Ng5869 & n4717;
  assign n4719 = n4716 & n4718_1;
  assign n4720 = ~n4715 & ~n4719;
  assign n4721 = n4711 & n4720;
  assign n4722 = ~Ng4087 & n4721;
  assign n4723 = Ng6219 & Ng6227;
  assign n4724 = Ng6215 & n4723;
  assign n4725 = n4716 & n4724;
  assign n4726 = Ng5535 & Ng5527;
  assign n4727 = Ng5523 & n4726;
  assign n4728_1 = n4522 & n4727;
  assign n4729 = ~n4725 & ~n4728_1;
  assign n4730 = Ng3179 & Ng3171;
  assign n4731 = Ng3167 & n4730;
  assign n4732_1 = n4712 & n4731;
  assign n4733 = Ng3873 & Ng3881;
  assign n4734 = Ng3869 & n4733;
  assign n4735 = n4704 & n4734;
  assign n4736 = ~n4732_1 & ~n4735;
  assign n4737 = Ng4087 & n4736;
  assign n4738 = n4729 & n4737;
  assign n4739 = n4703 & ~n4738;
  assign n2028 = ~n4722 & n4739;
  assign n4741 = n4562 & ~n2028;
  assign Pg33659 = ~n4703 | ~n4741;
  assign n4743 = Ng4765 & n4613_1;
  assign n4744 = Ng4709 & ~Ng4785;
  assign n4745 = Ng4754 & n4744;
  assign n4746 = ~n4743 & ~n4745;
  assign n4747 = ~Ng4709 & Ng4785;
  assign n4748 = Ng4743 & n4747;
  assign n4749 = ~n4679 & ~n4748;
  assign n2499 = ~n4746 | ~n4749;
  assign Pg33636 = ~n4693_1 | n2499;
  assign n4752 = ~Ng1205 & ~Ng1221;
  assign n4753 = ~Ng1211 & n4752;
  assign n4754 = ~Ng1216 & Ng1061;
  assign n4755 = Ng979 & n4754;
  assign n4756 = n4753 & n4755;
  assign n4757 = ~Ng1183 & n4756;
  assign n4758 = Ng1171 & n4757;
  assign Pg33533 = Pg17291 & ~n4758;
  assign n4760 = Ng2724 & Ng2787;
  assign n4761 = Ng2783 & ~Ng2724;
  assign n4762_1 = Ng2729 & ~n4761;
  assign n4763 = ~n4760 & n4762_1;
  assign n4764 = ~Ng2724 & ~Ng2729;
  assign n4765 = ~Ng2771 & n4764;
  assign n4766 = Ng2724 & ~Ng2729;
  assign n4767 = ~Ng2775 & n4766;
  assign n4768 = ~n4765 & ~n4767;
  assign Pg33435 = n4763 | ~n4768;
  assign n4770 = ~Ng2815 & ~Ng2724;
  assign n4771 = ~Ng2819 & Ng2724;
  assign n4772 = Ng2729 & ~n4771;
  assign n4773 = ~n4770 & n4772;
  assign n4774 = Ng2803 & n4764;
  assign n4775 = Ng2807 & n4766;
  assign n4776 = ~n4774 & ~n4775;
  assign Pg33079 = ~n4773 & n4776;
  assign n4778 = Ng2917 & Ng2912;
  assign n4779 = Ng2960 & Ng2965;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = Ng2955 & Ng2950;
  assign n4782 = n4780 & ~n4781;
  assign n4783 = Ng2975 & Ng2970;
  assign n4784 = Ng2941 & Ng2936;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = Ng2927 & Ng2922;
  assign n4787 = Ng2907 & Ng2902;
  assign n4788_1 = ~n4786 & ~n4787;
  assign n4789 = n4785 & n4788_1;
  assign Pg32185 = n4782 & n4789;
  assign n4791 = ~Ng5124 & ~Ng6163;
  assign n4792 = ~Ng5817 & n4791;
  assign n4793 = Pg35 & Ng5471;
  assign n4794 = ~n4792 & n4793;
  assign n4795 = ~Ng4427 & ~Ng4420;
  assign n4796 = Pg35 & Ng3466;
  assign n4797 = n4795 & ~n4796;
  assign n4798_1 = Pg35 & Ng6509;
  assign n4799 = n4797 & ~n4798_1;
  assign n4800 = Ng5124 & Ng6163;
  assign n4801 = ~Ng5817 & ~n4800;
  assign n4802 = Pg35 & ~n4791;
  assign n4803_1 = ~n4801 & n4802;
  assign n4804 = n4799 & ~n4803_1;
  assign n4805 = ~n4794 & n4804;
  assign n4806 = ~Ng5471 & n4792;
  assign n4807 = ~Ng3115 & n4806;
  assign n4808 = ~Ng3817 & n4807;
  assign n4809 = Pg35 & ~n4808;
  assign n4810 = ~n4795 & n4796;
  assign n4811 = ~n4797 & n4798_1;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = ~n4809 & n4812;
  assign n4814 = ~n4805 & ~n4813;
  assign n4815 = Ng3115 & ~n4806;
  assign n4816 = ~Ng3817 & ~n4815;
  assign n4817 = Pg35 & ~n4807;
  assign n4818 = ~n4816 & n4817;
  assign Pg31793 = ~n4814 & ~n4818;
  assign n4820 = Pg35 & ~Ng1306;
  assign Pg28042 = Ng962 | ~n4820;
  assign n4822 = ~Ng1312 & ~Ng1351;
  assign n4823 = Ng1536 & ~n4822;
  assign n4824 = ~Ng969 & ~Ng1008;
  assign n4825 = Ng1193 & ~n4824;
  assign n4826 = Pg35 & ~n4825;
  assign Pg28041 = n4823 | ~n4826;
  assign n4828_1 = ~Ng5831 & ~Ng5845;
  assign n4829 = ~Ng5499 & ~Ng5485;
  assign n4830 = ~Ng6537 & ~Ng6523;
  assign n4831 = ~Ng6177 & ~Ng6191;
  assign n4832 = n4830 & n4831;
  assign n4833 = n4829 & n4832;
  assign n4834 = n4828_1 & n4833;
  assign n4835 = ~Ng3831 & ~Ng3845;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~Ng3143 & ~Ng3129;
  assign n4838 = ~Ng5138 & ~Ng5152;
  assign n4839 = ~Ng3494 & ~Ng3480;
  assign n4840 = n4838 & n4839;
  assign n4841 = Pg35 & ~n4840;
  assign n4842 = n4837 & ~n4841;
  assign n4843_1 = ~n4830 & ~n4831;
  assign n4844 = n4828_1 & ~n4843_1;
  assign n4845 = ~n4833 & ~n4844;
  assign n4846 = ~n4829 & ~n4832;
  assign n4847_1 = ~n4845 & ~n4846;
  assign n4848 = n4842 & n4847_1;
  assign n4849 = ~n4836 & n4848;
  assign n4850 = n4834 & n4835;
  assign n4851 = ~n4838 & ~n4839;
  assign n4852 = n4837 & ~n4851;
  assign n4853 = ~n4840 & ~n4852;
  assign n4854 = n4850 & ~n4853;
  assign n4855 = Pg35 & ~n4854;
  assign Pg28030 = n4849 | ~n4855;
  assign n4857 = ~Ng1664 & ~Ng2047;
  assign n4858 = ~Ng1798 & ~Ng2066;
  assign n4859 = n4857 & n4858;
  assign n4860 = ~Ng1932 & ~Ng1644;
  assign n4861 = ~Ng1779 & n4860;
  assign n4862 = n4859 & n4861;
  assign n4863 = ~Ng1913 & n4862;
  assign n4864 = ~Ng2223 & ~Ng2625;
  assign n4865_1 = ~Ng2606 & ~Ng2357;
  assign n4866 = ~Ng2472 & n4865_1;
  assign n4867 = n4864 & n4866;
  assign n4868 = ~Ng2338 & ~Ng2491;
  assign n4869_1 = ~Ng2204 & n4868;
  assign n4870 = n4867 & n4869_1;
  assign n4871 = Pg35 & ~n4870;
  assign Pg26877 = n4863 | ~n4871;
  assign n4873 = ~Ng1858 & ~Ng1710;
  assign n4874_1 = ~Ng1844 & ~Ng1978;
  assign n4875 = ~Ng1992 & ~Ng2126;
  assign n4876 = n4874_1 & n4875;
  assign n4877 = ~Ng2112 & ~Ng1724;
  assign n4878 = n4876 & n4877;
  assign n4879 = n4873 & n4878;
  assign n4880 = ~Ng2671 & ~Ng2685;
  assign n4881 = ~Ng2269 & ~Ng2283;
  assign n4882 = n4880 & n4881;
  assign n4883 = ~Ng2417 & ~Ng2551;
  assign n4884 = ~Ng2403 & ~Ng2537;
  assign n4885 = n4883 & n4884;
  assign n4886 = n4882 & n4885;
  assign n4887 = Pg35 & ~n4886;
  assign Pg26876 = n4879 | ~n4887;
  assign n4889 = ~Ng1830 & ~Ng1964;
  assign n4890 = ~Ng1696 & ~Ng2098;
  assign n4891_1 = n4889 & n4890;
  assign n4892 = ~Ng2255 & ~Ng2523;
  assign n4893 = ~Ng2657 & n4892;
  assign n4894 = ~Ng2389 & n4893;
  assign n4895 = Pg35 & ~n4894;
  assign Pg26875 = n4891_1 | ~n4895;
  assign Pg23190 = ~Ng22 & ~Ng25;
  assign Pg21727 = ~Pg35 & Ng3003;
  assign n4899 = ~Pg35 & Ng5052;
  assign n4900 = Ng5029 & Ng5062;
  assign n4901 = Ng5016 & n4900;
  assign n4902 = Ng5033 & n4901;
  assign n4903 = Ng5037 & n4902;
  assign n4904 = Ng5041 & n4903;
  assign n4905_1 = Ng5046 & n4904;
  assign n4906 = Ng5052 & ~n4905_1;
  assign n4907 = Ng5022 & ~Ng5016;
  assign n4908 = ~Ng5029 & n4907;
  assign n4909 = ~Ng5033 & n4908;
  assign n4910 = ~Ng5037 & n4909;
  assign n4911 = ~Ng5041 & n4910;
  assign n4912 = ~Ng5046 & n4911;
  assign n4913 = ~Ng5052 & ~n4912;
  assign n4914 = ~n4906 & ~n4913;
  assign n4915 = ~Pg84 & ~Ng5052;
  assign n4916 = Pg84 & ~Ng5041;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = Ng5057 & ~Ng5046;
  assign n4919 = Ng5022 & n4918;
  assign n4920_1 = ~n4917 & n4919;
  assign n4921 = Pg35 & ~n4920_1;
  assign n4922 = Ng5057 & n4921;
  assign n4923 = ~n4914 & n4922;
  assign n4924 = ~n4899 & ~n4923;
  assign n4925_1 = ~Ng5057 & n4914;
  assign n4926 = Pg35 & n4925_1;
  assign n688 = ~n4924 | n4926;
  assign n4928 = ~Pg113 & ~n4561;
  assign n4929 = Ng2767 & ~n4928;
  assign n4930 = Ng2735 & n4632;
  assign n4931 = n4764 & n4930;
  assign n4932 = Ng85 & n4928;
  assign n4933 = n4931 & ~n4932;
  assign n4934 = ~n4929 & n4933;
  assign n4935 = Ng2771 & ~n4931;
  assign n4936 = Pg35 & ~n4935;
  assign n4937 = ~n4934 & n4936;
  assign n4938 = ~Pg35 & ~Ng2775;
  assign n693 = ~n4937 & ~n4938;
  assign n4940 = Ng1183 & n4756;
  assign n4941 = Ng1171 & n4940;
  assign n4942 = Pg17400 & ~n4941;
  assign n4943 = ~Ng209 & Ng691;
  assign n4944 = n4825 & n4943;
  assign n4945 = ~Pg134 & ~n4944;
  assign n4946 = ~n4294 & ~n4945;
  assign n4947 = Ng2130 & Ng2138;
  assign n4948 = ~Ng2145 & n4947;
  assign n4949 = n4946 & ~n4948;
  assign n4950 = ~n4942 & n4949;
  assign n4951 = Ng1862 & ~n4950;
  assign n4952 = Ng1936 & n4951;
  assign n4953 = Pg35 & ~n4952;
  assign n4954 = Ng1882 & n4953;
  assign n4955 = ~Pg35 & Ng1886;
  assign n4956 = \[4421]  & ~n4948;
  assign n4957 = Ng4180 & n4946;
  assign n4958 = ~n4949 & ~n4957;
  assign n4959 = ~n4956 & ~n4958;
  assign n4960 = Pg35 & ~n4959;
  assign n4961 = ~n4955 & ~n4960;
  assign n4962 = ~n4953 & ~n4961;
  assign n698_1 = n4954 | n4962;
  assign n4964 = ~Ng1564 & ~Ng1554;
  assign n4965 = ~Ng1559 & n4964;
  assign n4966 = Ng1404 & Ng1322;
  assign n4967 = ~Ng1548 & n4966;
  assign n4968 = n4965 & n4967;
  assign n4969 = ~Ng1514 & n4968;
  assign n4970 = Ng1526 & n4969;
  assign n4971 = Pg17404 & ~n4970;
  assign n4972 = n4823 & n4943;
  assign n4973 = ~Pg134 & ~n4972;
  assign n4974_1 = ~n4439 & ~n4973;
  assign n4975 = Ng2689 & ~Ng2697;
  assign n4976 = Ng2704 & n4975;
  assign n4977 = n4974_1 & ~n4976;
  assign n4978 = ~n4971 & n4977;
  assign n4979_1 = ~Ng2287 & ~Ng2361;
  assign n4980 = ~n4978 & n4979_1;
  assign n4981 = Pg35 & ~n4980;
  assign n4982 = ~Ng1585 & ~n4976;
  assign n4983 = Ng4180 & n4974_1;
  assign n4984 = ~n4977 & ~n4983;
  assign n4985 = ~n4982 & ~n4984;
  assign n4986 = Pg35 & ~n4985;
  assign n4987 = ~Pg35 & Ng2380;
  assign n4988_1 = ~n4986 & ~n4987;
  assign n4989 = ~n4981 & n4988_1;
  assign n4990 = ~Ng2299 & n4981;
  assign n703_1 = ~n4989 & ~n4990;
  assign n4992 = ~Pg35 & Ng4031;
  assign n4993_1 = Pg13966 & Pg11418;
  assign n4994 = Pg16659 & n4993_1;
  assign n4995 = Pg16775 & n4994;
  assign n4996 = ~Ng4040 & ~n4995;
  assign n4997 = Ng4040 & n4995;
  assign n4998 = Pg35 & ~n4997;
  assign n4999 = ~n4996 & n4998;
  assign n708_1 = n4992 | n4999;
  assign n5001 = Ng2719 & ~Ng2715;
  assign n5002 = ~Ng2735 & n4764;
  assign n5003_1 = ~n4662 & n4764;
  assign n5004 = ~n5002 & ~n5003_1;
  assign n5005 = n5001 & n5004;
  assign n5006 = Ng2815 & n4764;
  assign n5007 = n5005 & ~n5006;
  assign n5008_1 = Ng2485 & n5007;
  assign n5009 = Ng2453 & n5008_1;
  assign n5010 = Pg35 & ~n5009;
  assign n5011 = Ng2547 & n5010;
  assign n5012 = Ng2541 & ~n5010;
  assign n713_1 = n5011 | n5012;
  assign n5014 = ~Pg35 & ~Ng3227;
  assign n5015 = ~Ng3155 & Ng3161;
  assign n5016 = n4730 & n5015;
  assign n5017_1 = ~Ng4284 & Ng4180;
  assign n5018 = Pg35 & n5017_1;
  assign n5019 = n5016 & n5018;
  assign n5020 = Pg35 & ~Ng3243;
  assign n5021 = ~n5016 & n5020;
  assign n5022_1 = ~n5019 & ~n5021;
  assign n722_1 = ~n5014 & n5022_1;
  assign n5024 = Ng358 & Ng376;
  assign n5025 = Ng385 & n5024;
  assign n5026 = ~Ng370 & n5025;
  assign n5027_1 = Pg35 & ~n5026;
  assign n5028 = Ng452 & n5027_1;
  assign n5029 = Ng460 & ~n5027_1;
  assign n727_1 = n5028 | n5029;
  assign n5031 = ~Pg35 & ~Ng3546;
  assign n5032_1 = ~Ng3530 & Ng3522;
  assign n5033 = ~Ng3512 & ~Ng3518;
  assign n5034 = ~Ng3506 & n5033;
  assign n5035 = n5032_1 & n5034;
  assign n5036 = ~n5018 & n5035;
  assign n5037_1 = Pg35 & ~Ng3542;
  assign n5038 = ~n5035 & ~n5037_1;
  assign n5039 = ~n5036 & ~n5038;
  assign n732_1 = ~n5031 & ~n5039;
  assign n5041 = ~Ng5180 & Ng5188;
  assign n5042_1 = Ng5164 & ~Ng5170;
  assign n5043 = n5041 & n5042_1;
  assign n5044 = Pg35 & ~n5043;
  assign n5045 = ~Pg35 & ~Ng5208;
  assign n5046 = ~n5018 & ~n5045;
  assign n5047 = ~n5044 & ~n5046;
  assign n5048 = ~Ng5232 & n5044;
  assign n737_1 = ~n5047 & ~n5048;
  assign n5050 = Pg35 & ~n4718_1;
  assign n5051 = Ng5813 & n5050;
  assign n5052 = Ng5849 & ~n5050;
  assign n742_1 = n5051 | n5052;
  assign n5054 = Pg35 & Ng2907;
  assign n5055 = ~Pg35 & Ng2984;
  assign n747_1 = n5054 | n5055;
  assign n5057 = ~Ng1171 & n4940;
  assign n5058 = Pg17316 & ~n5057;
  assign n5059 = ~n4431 & ~n4945;
  assign n5060 = Ng2130 & ~Ng2138;
  assign n5061_1 = Ng2145 & n5060;
  assign n5062 = n5059 & ~n5061_1;
  assign n5063 = ~n5058 & n5062;
  assign n5064 = Ng1772 & ~n5063;
  assign n5065_1 = ~Ng1802 & n5064;
  assign n5066 = ~\[4421]  & ~n5061_1;
  assign n5067 = Ng4180 & n5059;
  assign n5068 = ~n5062 & ~n5067;
  assign n5069 = ~n5066 & ~n5068;
  assign n5070 = Pg35 & ~n5069;
  assign n5071 = n5065_1 & n5070;
  assign n5072 = ~Pg35 & Ng1736;
  assign n5073 = Pg35 & Ng1744;
  assign n5074 = ~n5065_1 & n5073;
  assign n5075 = ~n5072 & ~n5074;
  assign n752_1 = n5071 | ~n5075;
  assign n5077 = ~Ng5869 & ~Ng5857;
  assign n5078 = ~Ng5863 & n5077;
  assign n5079 = n4717 & n5078;
  assign n5080_1 = Pg35 & ~n5079;
  assign n5081 = Ng5909 & n5080_1;
  assign n5082 = ~Pg35 & Ng5913;
  assign n5083 = Pg35 & ~n5017_1;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = ~n5080_1 & ~n5084;
  assign n757_1 = n5081 | n5085;
  assign n5087 = Pg35 & n5063;
  assign n5088 = Ng1802 & n5087;
  assign n5089 = Ng112 & n4928;
  assign n5090 = n4592 & n5089;
  assign n5091 = Pg35 & n5090;
  assign n5092 = Ng1772 & ~n5091;
  assign n5093 = ~n5087 & n5092;
  assign n762_1 = n5088 | n5093;
  assign n5095 = Ng3518 & Ng3522;
  assign n5096 = ~Ng3530 & n5095;
  assign n5097 = n5018 & n5096;
  assign n5098 = ~Pg35 & ~Ng3602;
  assign n5099_1 = ~n5097 & ~n5098;
  assign n5100 = Pg35 & ~n5096;
  assign n5101 = ~Ng3554 & n5100;
  assign n767_1 = n5099_1 & ~n5101;
  assign n5103 = Ng43 & n4928;
  assign n5104_1 = n4703 & n5103;
  assign n5105 = Ng4087 & n5104_1;
  assign n5106 = n4716 & n5105;
  assign n5107 = ~Ng6219 & ~n5106;
  assign n5108_1 = Pg35 & ~n5107;
  assign n5109 = Ng6215 & ~n5108_1;
  assign n5110 = Pg35 & ~n5106;
  assign n5111 = ~Ng6215 & n5110;
  assign n5112_1 = Ng6219 & n5111;
  assign n772_1 = n5109 | n5112_1;
  assign n5114 = ~Pg35 & Ng794;
  assign n5115 = ~Ng736 & Pg11678;
  assign n5116 = ~Ng518 & ~Ng499;
  assign n5117_1 = ~Ng528 & ~Ng482;
  assign n5118 = n5116 & n5117_1;
  assign n5119 = ~Ng490 & n5118;
  assign n5120 = n5026 & n5119;
  assign n5121 = Ng807 & Ng554;
  assign n5122 = Ng718 & Ng655;
  assign n5123 = Ng753 & ~n5122;
  assign n5124 = ~Ng718 & ~Ng655;
  assign n5125 = ~Ng753 & ~n5124;
  assign n5126 = ~n5123 & ~n5125;
  assign n5127_1 = ~n5121 & ~n5126;
  assign n5128 = n5120 & n5127_1;
  assign n5129 = Pg12184 & ~Pg11678;
  assign n5130 = n5128 & ~n5129;
  assign n5131 = Ng739 & n5130;
  assign n5132 = ~n5115 & n5131;
  assign n5133 = Ng744 & n5132;
  assign n5134 = Ng749 & n5133;
  assign n5135 = Ng758 & n5134;
  assign n5136 = Ng763 & n5135;
  assign n5137 = Ng767 & n5136;
  assign n5138 = Ng772 & n5137;
  assign n5139 = Ng776 & n5138;
  assign n5140 = Ng781 & n5139;
  assign n5141 = Ng785 & n5140;
  assign n5142 = Ng790 & n5141;
  assign n5143 = Ng794 & n5142;
  assign n5144 = Ng807 & n5143;
  assign n5145 = Pg35 & ~n5115;
  assign n5146 = Ng807 & n5145;
  assign n5147 = ~n5143 & ~n5146;
  assign n5148 = ~n5144 & ~n5147;
  assign n777_1 = n5114 | n5148;
  assign n5150 = Ng370 & n5025;
  assign n5151 = Pg35 & ~n5150;
  assign n5152 = Ng847 & n5151;
  assign n5153 = Ng854 & ~n5151;
  assign n786_1 = n5152 | n5153;
  assign n5155 = Pg35 & ~Pg12919;
  assign n5156 = ~Ng1061 & n5155;
  assign n5157_1 = Pg35 & Ng1052;
  assign n5158 = ~Ng1061 & ~n5157_1;
  assign n5159 = ~n5155 & ~n5158;
  assign n5160 = Pg35 & ~Pg19334;
  assign n5161_1 = ~n5159 & ~n5160;
  assign n791_1 = n5156 | ~n5161_1;
  assign n5163 = ~Ng4172 & ~Ng4153;
  assign n796_1 = Pg35 & ~n5163;
  assign n5165 = ~Pg35 & ~Ng4366;
  assign n5166_1 = ~n4531 & ~n4540;
  assign n5167 = Ng4340 & n5166_1;
  assign n5168 = Ng4593 & ~Ng4601;
  assign n5169 = Ng4584 & ~Ng4608;
  assign n5170 = n5168 & n5169;
  assign n5171_1 = ~Ng4584 & Ng4608;
  assign n5172 = ~Ng4593 & n5171_1;
  assign n5173 = ~Ng4593 & Ng4601;
  assign n5174 = ~n5168 & ~n5173;
  assign n5175 = ~Ng4616 & n5174;
  assign n5176 = ~n5169 & n5175;
  assign n5177 = ~n5171_1 & n5176;
  assign n5178 = ~n5172 & ~n5177;
  assign n5179 = ~n5170 & n5178;
  assign n5180 = ~Pg135 & ~n5179;
  assign n5181 = ~n4537 & ~n5180;
  assign n5182 = ~Pg73 & ~Pg72;
  assign n5183 = Ng4322 & ~Ng4515;
  assign n5184 = n5182 & ~n5183;
  assign n5185 = ~Ng4332 & n5184;
  assign n5186 = ~Ng4322 & Ng4311;
  assign n5187 = Ng4332 & ~n5186;
  assign n5188 = ~n5185 & ~n5187;
  assign n5189 = ~Ng4332 & ~Ng4322;
  assign n5190 = ~Ng2994 & n5189;
  assign n5191_1 = Pg90 & n5190;
  assign n5192 = n4537 & ~n5191_1;
  assign n5193 = ~n5188 & n5192;
  assign n5194 = ~Ng4340 & ~n5193;
  assign n5195 = ~n5181 & n5194;
  assign n5196 = Pg35 & ~n5195;
  assign n5197 = ~n5167 & n5196;
  assign n801_1 = ~n5165 & ~n5197;
  assign n5199 = ~Pg35 & Ng3506;
  assign n5200 = ~Ng3512 & Ng3506;
  assign n5201 = Ng3512 & ~Ng3506;
  assign n5202 = ~n5200 & ~n5201;
  assign n5203 = ~Ng4087 & n5104_1;
  assign n5204 = n4704 & n5203;
  assign n5205 = Pg35 & ~n5204;
  assign n5206 = ~n5202 & n5205;
  assign n806_1 = n5199 | n5206;
  assign n5208 = ~Pg35 & Ng744;
  assign n5209 = Ng749 & n5145;
  assign n5210 = ~n5133 & ~n5209;
  assign n5211 = ~n5134 & ~n5210;
  assign n811_1 = n5208 | n5211;
  assign n5213 = Pg35 & ~n4706;
  assign n5214 = Ng3490 & n5213;
  assign n5215 = Ng3484 & ~n5213;
  assign n816_1 = n5214 | n5215;
  assign n5217 = Pg12350 & Pg14738;
  assign n5218 = ~Pg14738 & ~Pg17739;
  assign n5219 = ~n5217 & ~n5218;
  assign n5220 = Pg35 & ~Pg17646;
  assign n5221 = ~Pg17607 & ~Pg13068;
  assign n5222 = n5220 & n5221;
  assign n821_1 = ~n5219 & n5222;
  assign n5224 = ~n4283 & ~n4945;
  assign n5225 = ~Ng2145 & n5060;
  assign n5226 = n5224 & ~n5225;
  assign n5227 = ~Pg33533 & n5226;
  assign n5228 = ~Ng1636 & ~n5227;
  assign n5229 = Ng1592 & n5228;
  assign n5230 = Pg35 & ~n5229;
  assign n5231 = Ng1600 & n5230;
  assign n5232 = ~Pg35 & Ng1604;
  assign n5233 = \[4421]  & ~n5225;
  assign n5234 = Ng4180 & n5224;
  assign n5235 = ~n5226 & ~n5234;
  assign n5236 = ~n5233 & ~n5235;
  assign n5237 = Pg35 & ~n5236;
  assign n5238 = ~n5232 & ~n5237;
  assign n5239 = ~n5230 & ~n5238;
  assign n829_1 = n5231 | n5239;
  assign n5241 = ~Pg35 & Ng1710;
  assign n5242 = Pg35 & ~Ng1714;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = Pg35 & n5227;
  assign n5245 = ~Ng1668 & ~Ng1592;
  assign n5246 = Pg35 & ~n5245;
  assign n5247 = ~n5244 & ~n5246;
  assign n5248 = n5243 & n5247;
  assign n5249 = ~Ng1714 & ~n5247;
  assign n834_1 = ~n5248 & ~n5249;
  assign n5251 = n4712 & n5105;
  assign n5252 = Pg35 & ~n5251;
  assign n5253 = ~Ng3167 & n5252;
  assign n842_1 = ~Ng3155 & n5253;
  assign n5255 = ~Pg35 & Ng2217;
  assign n5256 = ~Ng2719 & ~Ng2715;
  assign n5257 = n5004 & n5256;
  assign n5258 = ~n4774 & n5257;
  assign n5259 = Pg35 & ~n5258;
  assign n5260 = Ng2236 & n5259;
  assign n5261 = Pg35 & n5258;
  assign n5262 = Ng2208 & ~Ng2185;
  assign n5263 = Ng2161 & n5262;
  assign n5264 = Ng2181 & n4645_1;
  assign n5265 = ~Ng2208 & Ng2185;
  assign n5266 = Ng2177 & n5265;
  assign n5267 = ~n5264 & ~n5266;
  assign n5268 = ~Ng2208 & Ng2217;
  assign n5269 = Ng2169 & n5268;
  assign n5270_1 = Ng2173 & ~Ng2217;
  assign n5271 = ~Ng2185 & n5270_1;
  assign n5272 = ~n5269 & ~n5271;
  assign n5273 = n5267 & n5272;
  assign n5274 = ~n5263 & n5273;
  assign n5275 = n5261 & ~n5274;
  assign n5276 = ~n5260 & ~n5275;
  assign n5277 = Ng2185 & Ng2217;
  assign n5278 = n5258 & n5277;
  assign n5279_1 = Ng2165 & n5278;
  assign n5280 = n5276 & ~n5279_1;
  assign n847_1 = n5255 | ~n5280;
  assign n5282 = Pg13926 & Pg11388;
  assign n5283 = Pg16627 & n5282;
  assign n5284 = Pg16744 & n5283;
  assign n5285 = Ng3689 & n5284;
  assign n5286 = Pg35 & n5285;
  assign n857_1 = Ng3694 & ~n5286;
  assign n5288 = ~Ng1772 & ~n5063;
  assign n5289_1 = Ng1728 & n5288;
  assign n5290 = Pg35 & ~n5289_1;
  assign n5291 = Ng1736 & n5290;
  assign n5292 = ~Pg35 & Ng1740;
  assign n5293 = ~n5070 & ~n5292;
  assign n5294_1 = ~n5290 & ~n5293;
  assign n862_1 = n5291 | n5294_1;
  assign n5296 = Ng2783 & n4764;
  assign n5297 = n5005 & ~n5296;
  assign n5298 = Ng1926 & n5297;
  assign n5299 = Ng1894 & n5298;
  assign n5300 = Pg35 & ~n5299;
  assign n5301 = ~Ng1968 & n5300;
  assign n5302 = Pg35 & ~Ng1968;
  assign n5303 = ~Pg35 & Ng1964;
  assign n5304 = ~n5302 & ~n5303;
  assign n5305 = ~n5300 & n5304;
  assign n867_1 = ~n5301 & ~n5305;
  assign n5307 = ~Ng4621 & ~Ng4639;
  assign n5308 = ~n4928 & n5182;
  assign n5309 = Ng65 & ~n5308;
  assign n5310 = ~Ng4643 & ~n5309;
  assign n5311 = Pg35 & n5310;
  assign n5312 = Ng4621 & Ng4639;
  assign n5313 = n5311 & ~n5312;
  assign n5314_1 = ~Pg35 & Ng4639;
  assign n5315 = ~n5313 & ~n5314_1;
  assign n872_1 = ~n5307 & ~n5315;
  assign n5317 = ~Ng5535 & Ng5527;
  assign n5318 = Ng5511 & Ng5517;
  assign n5319 = n5317 & n5318;
  assign n5320 = n5083 & n5319;
  assign n5321 = ~Pg35 & Ng5591;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = Pg35 & Ng5607;
  assign n5324 = ~n5319 & n5323;
  assign n877_1 = ~n5322 | n5324;
  assign n5326 = Ng2819 & n4764;
  assign n5327 = Ng2719 & Ng2715;
  assign n5328 = n5004 & n5327;
  assign n5329 = ~n5326 & n5328;
  assign n5330 = Pg35 & ~n5329;
  assign n5331 = Ng2610 & ~Ng2587;
  assign n5332 = Pg35 & ~n5331;
  assign n5333 = ~n5330 & ~n5332;
  assign n5334 = Ng2657 & ~n5333;
  assign n5335 = Pg35 & Ng2648;
  assign n5336 = ~Ng2652 & n5335;
  assign n5337 = Ng2652 & ~n5335;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = n5333 & ~n5338;
  assign n882_1 = n5334 | n5339;
  assign n5341 = Pg12300 & Pg14694;
  assign n5342 = ~Pg17711 & ~Pg14694;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = Pg35 & ~Pg17580;
  assign n5345 = ~Pg13049 & n5344;
  assign n5346 = ~Pg17604 & n5345;
  assign n887_1 = ~n5343 & n5346;
  assign n5348 = Ng667 & ~Ng686;
  assign n5349 = Pg35 & n5348;
  assign n5350 = Ng358 & Ng385;
  assign n5351 = ~Ng376 & n5350;
  assign n5352 = ~Ng513 & Ng518;
  assign n5353 = n5351 & n5352;
  assign n5354 = Ng490 & Ng482;
  assign n5355 = ~Ng528 & ~n5354;
  assign n5356 = n5353 & ~n5355;
  assign n5357 = Ng482 & n5356;
  assign n5358 = Pg35 & ~n5357;
  assign n5359 = Ng490 & n5358;
  assign n5360 = ~Ng490 & n5356;
  assign n5361 = Pg35 & ~n5360;
  assign n5362 = Ng482 & ~n5361;
  assign n5363 = ~n5359 & ~n5362;
  assign n891_1 = n5349 | ~n5363;
  assign n5365 = Pg6744 & Pg35;
  assign n5366 = ~Pg35 & Ng305;
  assign n896_1 = n5365 | n5366;
  assign n5368 = ~Pg35 & Ng767;
  assign n5369 = Ng772 & n5145;
  assign n5370 = ~n5137 & ~n5369;
  assign n5371 = ~n5138 & ~n5370;
  assign n901_1 = n5368 | n5371;
  assign n5373 = ~Ng5511 & Ng5517;
  assign n5374 = ~Ng5535 & ~Ng5527;
  assign n5375 = n5373 & n5374;
  assign n5376 = Pg35 & ~n5375;
  assign n5377 = ~Pg35 & ~Ng5571;
  assign n5378 = ~n5018 & ~n5377;
  assign n5379 = ~n5376 & ~n5378;
  assign n5380 = ~Ng5587 & n5376;
  assign n906_1 = ~n5379 & ~n5380;
  assign n5382 = Pg17685 & n4547;
  assign n5383 = Ng6381 & n5382;
  assign n5384 = n4677 & n4743;
  assign n5385 = Ng4688 & ~n5384;
  assign n5386 = n5383 & n5385;
  assign n5387 = Pg35 & ~n5386;
  assign n5388 = Pg35 & ~Ng6167;
  assign n5389 = Ng6173 & n5388;
  assign n5390 = ~Ng6173 & ~n5388;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~n5387 & ~n5391;
  assign n5393 = ~Ng6177 & n5387;
  assign n911_1 = ~n5392 & ~n5393;
  assign n5395 = ~Pg35 & Ng3161;
  assign n5396 = Ng3155 & Ng3161;
  assign n5397 = n5253 & n5396;
  assign n920_1 = n5395 | n5397;
  assign n5399 = n4726 & n5318;
  assign n5400 = Pg35 & ~n5399;
  assign n5401 = Ng5615 & n5400;
  assign n5402 = ~Pg35 & Ng5599;
  assign n5403 = ~n5083 & ~n5402;
  assign n5404 = ~n5400 & ~n5403;
  assign n925_1 = n5401 | n5404;
  assign n5406 = Pg35 & Ng4581;
  assign n5407 = Pg73 & ~Pg72;
  assign n5408 = n5406 & ~n5407;
  assign n5409 = Ng4575 & n5406;
  assign n5410 = Ng4543 & ~n5406;
  assign n5411 = ~n5409 & ~n5410;
  assign n930 = n5408 | ~n5411;
  assign n5413 = ~Ng3639 & Ng3703;
  assign n5414 = Ng3594 & n5413;
  assign n5415 = Pg16744 & n5414;
  assign n5416 = Ng3689 & ~Pg11388;
  assign n5417 = ~Ng3689 & Pg11388;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = Ng3639 & ~Ng3703;
  assign n5420 = Pg16627 & Ng3610;
  assign n5421 = n5419 & n5420;
  assign n5422 = ~Ng3639 & ~Ng3703;
  assign n5423 = Pg13926 & Ng3578;
  assign n5424 = n5422 & n5423;
  assign n5425 = ~n5421 & ~n5424;
  assign n5426 = ~n5418 & n5425;
  assign n5427 = ~n5415 & n5426;
  assign n5428 = Pg16744 & n4541;
  assign n5429 = Ng3586 & n5428;
  assign n5430 = Ng3570 & Pg13926;
  assign n5431 = n5419 & n5430;
  assign n5432_1 = Pg16627 & Ng3602;
  assign n5433 = n5422 & n5432_1;
  assign n5434 = ~n5431 & ~n5433;
  assign n5435 = n5418 & n5434;
  assign n5436 = ~n5429 & n5435;
  assign n5437 = ~n5427 & ~n5436;
  assign n5438 = Pg14451 & Ng3550;
  assign n5439 = Ng3680 & Ng3562;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = n5419 & ~n5440;
  assign n5442 = Ng3606 & Pg16722;
  assign n5443 = Ng3554 & Pg16656;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = n5413 & ~n5444;
  assign n5446 = ~n5441 & ~n5445;
  assign n5447_1 = Ng3574 & Pg16924;
  assign n5448 = Ng3558 & Pg11388;
  assign n5449 = ~n5447_1 & ~n5448;
  assign n5450 = n4541 & ~n5449;
  assign n5451 = ~Ng3689 & ~n5450;
  assign n5452 = Ng3590 & n5422;
  assign n5453 = Pg13881 & n5452;
  assign n5454 = n5451 & ~n5453;
  assign n5455 = n5446 & n5454;
  assign n5456 = Ng3566 & Pg16924;
  assign n5457_1 = Ng3542 & Pg11388;
  assign n5458 = ~n5456 & ~n5457_1;
  assign n5459 = n5413 & ~n5458;
  assign n5460 = Pg13881 & Ng3582;
  assign n5461 = n5419 & n5460;
  assign n5462 = Ng3689 & ~n5461;
  assign n5463 = Ng3598 & n4541;
  assign n5464 = Pg16722 & n5463;
  assign n5465 = Pg14451 & Ng3538;
  assign n5466 = Ng3680 & Ng3546;
  assign n5467 = ~n5465 & ~n5466;
  assign n5468 = n5422 & ~n5467;
  assign n5469 = ~n5464 & ~n5468;
  assign n5470 = n5462 & n5469;
  assign n5471 = ~n5459 & n5470;
  assign n5472 = ~n5455 & ~n5471;
  assign n5473 = ~n5437 & ~n5472;
  assign n5474 = Pg16656 & n4541;
  assign n5475 = Ng3689 & n5474;
  assign n5476 = Ng3614 & n5475;
  assign n5477 = n5473 & ~n5476;
  assign n5478 = ~Ng4983 & ~Ng4991;
  assign n5479 = Ng4966 & n5478;
  assign n5480 = Ng4843 & n4605;
  assign n5481 = n5479 & n5480;
  assign n5482 = n4687 & n5481;
  assign n5483 = Ng4871 & ~n5482;
  assign n5484 = Pg35 & n5483;
  assign n5485 = ~n5477 & n5484;
  assign n5486 = ~Ng3457 & n5485;
  assign n5487 = n5475 & n5483;
  assign n5488 = n5477 & n5487;
  assign n5489 = Pg35 & Ng3457;
  assign n5490 = ~n5473 & n5483;
  assign n5491 = ~n5475 & n5490;
  assign n5492 = n5489 & ~n5491;
  assign n5493 = ~n5488 & n5492;
  assign n5494 = ~Pg35 & Ng3462;
  assign n5495 = ~n5493 & ~n5494;
  assign n935_1 = n5486 | ~n5495;
  assign n5497 = Ng6209 & ~Ng6203;
  assign n5498 = ~Ng6219 & Ng6227;
  assign n5499 = n5497 & n5498;
  assign n5500 = Pg35 & ~n5499;
  assign n5501 = ~Pg35 & ~Ng6271;
  assign n5502 = ~n5018 & ~n5501;
  assign n5503 = ~n5500 & ~n5502;
  assign n5504 = ~Ng6287 & n5500;
  assign n940_1 = ~n5503 & ~n5504;
  assign n5506 = ~Ng1333 & ~Ng1322;
  assign n5507 = ~Ng1339 & ~Ng1322;
  assign n5508 = Ng1339 & Ng1322;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n5506 & n5509;
  assign n5511 = n4822 & n5510;
  assign n5512 = Ng1579 & Ng1322;
  assign n5513 = ~Ng1579 & ~Ng1322;
  assign n5514 = Pg35 & ~n5513;
  assign n5515 = ~n5512 & n5514;
  assign n5516 = n5511 & n5515;
  assign n5517 = ~Pg7946 & ~Pg19357;
  assign n5518 = ~Ng1333 & n5517;
  assign n5519 = ~Pg8475 & n5518;
  assign n5520 = ~Pg13272 & n5519;
  assign n5521 = n5516 & n5520;
  assign n5522 = Pg35 & n5520;
  assign n5523 = ~Pg35 & Ng1339;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n5516 & n5524;
  assign n945_1 = ~n5521 & ~n5525;
  assign n5527 = ~Ng1526 & n4969;
  assign n5528 = Ng1430 & ~n5527;
  assign n5529 = ~n4463 & ~n4973;
  assign n5530 = Ng2689 & Ng2697;
  assign n5531 = Ng2704 & n5530;
  assign n5532 = n5529 & ~n5531;
  assign n5533 = ~n5528 & n5532;
  assign n5534 = ~Ng2599 & ~n5533;
  assign n5535 = Ng2555 & n5534;
  assign n5536 = Pg35 & ~n5535;
  assign n5537 = Ng2563 & n5536;
  assign n5538 = ~Pg35 & Ng2567;
  assign n5539 = ~Ng1585 & ~n5531;
  assign n5540 = Ng4180 & n5529;
  assign n5541 = ~n5532 & ~n5540;
  assign n5542_1 = ~n5539 & ~n5541;
  assign n5543 = Pg35 & ~n5542_1;
  assign n5544 = ~n5538 & ~n5543;
  assign n5545 = ~n5536 & ~n5544;
  assign n949_1 = n5537 | n5545;
  assign n5547 = Ng63 & n4928;
  assign n5548 = n4498 & n5547;
  assign n5549 = Ng4793 & n4619;
  assign n5550 = Ng4776 & n5549;
  assign n5551 = ~n5548 & ~n5550;
  assign n5552 = Pg35 & n5551;
  assign n5553 = Ng4776 & n5552;
  assign n5554 = n5549 & n5551;
  assign n5555 = Pg35 & ~n5554;
  assign n5556 = Ng4801 & ~n5555;
  assign n954_1 = n5553 | n5556;
  assign n5558 = ~Pg35 & Ng4584;
  assign n5559 = Ng4621 & ~Ng4639;
  assign n5560 = Ng4340 & n5559;
  assign n5561 = Ng4628 & n5560;
  assign n5562 = Ng4349 & n5561;
  assign n5563 = Ng4358 & n5562;
  assign n5564 = Ng4332 & n5563;
  assign n5565 = Ng4322 & n5564;
  assign n5566 = Ng4584 & n5565;
  assign n5567 = Ng4616 & n5566;
  assign n5568 = ~n5309 & ~n5567;
  assign n5569 = Ng4593 & n5566;
  assign n5570 = Pg35 & Ng4593;
  assign n5571 = ~n5566 & ~n5570;
  assign n5572 = ~n5569 & ~n5571;
  assign n5573 = n5568 & n5572;
  assign n959_1 = n5558 | n5573;
  assign n964_1 = Pg35 & Ng6199;
  assign n5576 = ~Ng2331 & ~n4978;
  assign n5577 = Ng2287 & n5576;
  assign n5578 = Pg35 & ~n5577;
  assign n5579 = Ng2295 & n5578;
  assign n5580 = ~Pg35 & Ng2299;
  assign n5581 = ~n4986 & ~n5580;
  assign n5582 = ~n5578 & ~n5581;
  assign n969_1 = n5579 | n5582;
  assign n5584 = ~Pg35 & Ng1379;
  assign n5585 = ~Ng1384 & ~n5510;
  assign n5586 = ~Ng1384 & Ng1351;
  assign n5587 = n5510 & ~n5586;
  assign n5588 = Pg35 & ~n5587;
  assign n5589 = ~n5585 & n5588;
  assign n974_1 = n5584 | n5589;
  assign n5591 = Pg35 & Pg12923;
  assign n5592 = ~Pg35 & Ng1579;
  assign n979_1 = n5591 | n5592;
  assign n5594_1 = n4522 & n5203;
  assign n5595 = ~Ng5180 & ~n5594_1;
  assign n5596 = Pg35 & ~n5595;
  assign n5597 = Ng5176 & ~n5596;
  assign n5598 = Pg35 & ~n5594_1;
  assign n5599 = ~Ng5176 & n5598;
  assign n5600 = Ng5180 & n5599;
  assign n984_1 = n5597 | n5600;
  assign n5602 = Pg35 & Ng2844;
  assign n5603 = ~Pg35 & Ng2890;
  assign n989_1 = n5602 | n5603;
  assign n5605 = ~Pg35 & Ng1018;
  assign n5606 = ~Ng990 & ~Ng979;
  assign n5607 = ~Ng996 & ~Ng979;
  assign n5608 = Ng996 & Ng979;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = Ng1008 & ~Ng1046;
  assign n5611 = n5609 & ~n5610;
  assign n5612 = Ng1030 & Ng1018;
  assign n5613 = Ng1008 & n5612;
  assign n5614 = ~n5609 & n5613;
  assign n5615 = ~Ng969 & ~n5614;
  assign n5616 = ~n5611 & n5615;
  assign n5617 = ~Ng1002 & n5616;
  assign n5618 = ~n5606 & ~n5617;
  assign n5619 = ~Ng1018 & n5616;
  assign n5620 = n5618 & ~n5619;
  assign n5621 = ~Ng1024 & ~n5620;
  assign n5622 = ~Ng1024 & n5616;
  assign n5623 = n5620 & ~n5622;
  assign n5624_1 = Pg35 & ~n5623;
  assign n5625 = ~n5621 & n5624_1;
  assign n994_1 = n5605 | n5625;
  assign n5627 = n5317 & n5373;
  assign n5628 = n5018 & n5627;
  assign n5629_1 = ~Pg35 & ~Ng5575;
  assign n5630 = ~n5628 & ~n5629_1;
  assign n5631 = Pg35 & ~n5627;
  assign n5632 = ~Ng5591 & n5631;
  assign n999_1 = n5630 & ~n5632;
  assign n5634 = Ng3512 & Ng3506;
  assign n5635 = ~Ng3530 & ~Ng3522;
  assign n5636 = n5634 & n5635;
  assign n5637 = n5083 & n5636;
  assign n5638 = ~Pg35 & Ng3582;
  assign n5639_1 = ~n5637 & ~n5638;
  assign n5640 = Pg35 & Ng3598;
  assign n5641 = ~n5636 & n5640;
  assign n1004_1 = ~n5639_1 | n5641;
  assign n5643 = ~Ng4264 & ~Ng4258;
  assign n5687_1 = Pg35 & ~Ng4258;
  assign n5645 = Ng4264 & ~n5687_1;
  assign n5646 = ~Pg35 & Ng4258;
  assign n5647 = n5645 & ~n5646;
  assign n1009_1 = ~n5643 & ~n5647;
  assign n5649 = ~Pg35 & Ng763;
  assign n5650 = Ng767 & n5145;
  assign n5651 = ~n5136 & ~n5650;
  assign n5652 = ~n5137 & ~n5651;
  assign n1014_1 = n5649 | n5652;
  assign n1019_1 = Pg35 & Ng5853;
  assign n5655 = ~Ng1171 & n4757;
  assign n5656 = Ng1087 & ~n5655;
  assign n5657 = Ng2145 & n4947;
  assign n5658 = ~n4468 & ~n4945;
  assign n5659_1 = ~n5657 & n5658;
  assign n5660 = ~n5656 & n5659_1;
  assign n5661 = Pg35 & n5660;
  assign n5662 = ~Ng2070 & ~Ng1996;
  assign n5663 = Pg35 & ~n5662;
  assign n5664 = ~n5661 & ~n5663;
  assign n5665 = Ng2084 & n5664;
  assign n5666 = Ng2089 & ~n5664;
  assign n1027_1 = n5665 | n5666;
  assign n5668 = ~\[4661]  & ~n4561;
  assign n5669 = ~Ng4818 & n5668;
  assign n5670 = Ng71 & n5669;
  assign n5671 = n4609 & n4683_1;
  assign n5672_1 = ~n5670 & n5671;
  assign n5673 = Pg35 & ~n5672_1;
  assign n5674 = ~Ng4939 & ~n5673;
  assign n5675 = ~Ng4933 & ~n5671;
  assign n5676 = ~n5669 & ~n5675;
  assign n5677 = Pg35 & ~n5670;
  assign n5678 = ~n5676 & n5677;
  assign n1032_1 = ~n5674 & ~n5678;
  assign n5680 = ~Pg35 & ~Ng4512;
  assign n5681 = Ng4531 & n5406;
  assign n1037_1 = ~n5680 & ~n5681;
  assign n1042_1 = Pg35 & Ng5507;
  assign n5684 = n4723 & n5497;
  assign n5685 = n5018 & n5684;
  assign n5686 = Pg35 & ~Ng6291;
  assign n5687 = ~n5684 & n5686;
  assign n5688 = ~Pg35 & ~Ng6275;
  assign n5689 = ~n5687 & ~n5688;
  assign n1050_1 = ~n5685 & n5689;
  assign n5691_1 = ~Pg35 & Ng291;
  assign n5692 = ~Ng269 & ~Ng262;
  assign n5693 = ~Ng255 & n5692;
  assign n5694 = Ng246 & Ng239;
  assign n5695 = Ng225 & Ng232;
  assign n5696_1 = n5694 & n5695;
  assign n5697 = n5693 & n5696_1;
  assign n5698 = Ng278 & ~n5697;
  assign n5699 = Ng691 & ~n5128;
  assign n5700 = ~Ng225 & ~Ng232;
  assign n5701 = Ng269 & Ng262;
  assign n5702 = ~Ng246 & ~Ng239;
  assign n5703 = n5701 & n5702;
  assign n5704 = n5700 & n5703;
  assign n5705 = Ng255 & n5704;
  assign n5706 = ~Ng278 & ~n5705;
  assign n5707 = n5699 & ~n5706;
  assign n5708 = ~n5698 & n5707;
  assign n5709 = Ng287 & n5708;
  assign n5710 = Ng283 & n5709;
  assign n5711_1 = Ng291 & n5710;
  assign n5712 = Ng294 & n5711_1;
  assign n5713 = Pg35 & n5708;
  assign n5714 = Ng294 & n5713;
  assign n5715 = ~n5711_1 & ~n5714;
  assign n5716 = ~n5712 & ~n5715;
  assign n1055_1 = n5691_1 | n5716;
  assign n5718 = Ng5523 & Ng5527;
  assign n5719 = ~Ng5535 & n5718;
  assign n5720 = n5018 & n5719;
  assign n5721 = ~Pg35 & ~Ng5607;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = Pg35 & ~n5719;
  assign n5724 = ~Ng5559 & n5723;
  assign n1060 = n5722 & ~n5724;
  assign n1065_1 = Pg35 & Ng5881;
  assign n5727 = Pg35 & Ng6381;
  assign n5728 = ~Pg35 & Ng6098;
  assign n1069_1 = n5727 | n5728;
  assign n5730 = Pg35 & ~n4734;
  assign n5731 = Ng3813 & n5730;
  assign n5732 = Ng3849 & ~n5730;
  assign n1073_1 = n5731 | n5732;
  assign n5734 = ~Pg35 & Ng559;
  assign n5735 = Ng632 & Ng626;
  assign n5736 = ~Ng559 & Pg9048;
  assign n5737 = Pg35 & ~n5736;
  assign n5738 = ~Pg9048 & Pg12368;
  assign n5739_1 = \[4436]  & ~n5738;
  assign n5740 = Ng562 & n5739_1;
  assign n5741 = ~Ng562 & ~n5739_1;
  assign n5742 = ~n5740 & ~n5741;
  assign n5743 = n5737 & n5742;
  assign n5744 = ~n5735 & n5743;
  assign n1078_1 = n5734 | n5744;
  assign n5746 = ~Pg35 & Ng604;
  assign n5747 = ~n5736 & n5740;
  assign n5748 = Ng568 & n5747;
  assign n5749 = Ng572 & n5748;
  assign n5750 = Ng586 & n5749;
  assign n5751 = Ng577 & n5750;
  assign n5752 = Ng582 & n5751;
  assign n5753 = Ng590 & n5752;
  assign n5754 = Ng595 & n5753;
  assign n5755 = Ng599 & n5754;
  assign n5756 = Ng604 & n5755;
  assign n5757 = Ng608 & n5756;
  assign n5758 = Ng608 & n5737;
  assign n5759_1 = ~n5756 & ~n5758;
  assign n5760 = ~n5757 & ~n5759_1;
  assign n1083_1 = n5746 | n5760;
  assign n5762 = Pg35 & Ng1205;
  assign n5763 = ~Ng1087 & n5762;
  assign n5764_1 = Ng1087 & ~n5762;
  assign n1088_1 = n5763 | n5764_1;
  assign n5766 = ~Ng3869 & ~Ng3857;
  assign n5767 = ~Ng3863 & n5766;
  assign n5768 = n4733 & n5767;
  assign n5769_1 = Pg35 & ~n5768;
  assign n5770 = Ng3909 & n5769_1;
  assign n5771 = ~Pg35 & Ng3913;
  assign n5772 = ~n5083 & ~n5771;
  assign n5773_1 = ~n5769_1 & ~n5772;
  assign n1093_1 = n5770 | n5773_1;
  assign n5775 = Ng6215 & n5498;
  assign n5776 = n5083 & n5775;
  assign n5777 = ~Pg35 & Ng6303;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = Pg35 & Ng6259;
  assign n5780 = ~n5775 & n5779;
  assign n1098 = ~n5778 | n5780;
  assign n5782_1 = Ng5873 & Ng5869;
  assign n5783 = ~Ng5881 & n5782_1;
  assign n5784 = n5083 & n5783;
  assign n5785 = ~Pg35 & Ng5953;
  assign n5786 = ~n5784 & ~n5785;
  assign n5787_1 = Pg35 & Ng5905;
  assign n5788 = ~n5783 & n5787_1;
  assign n1103 = ~n5786 | n5788;
  assign n5790 = Pg35 & Ng921;
  assign n5791 = Ng904 & ~n5790;
  assign n5792_1 = ~Ng904 & n5790;
  assign n5793 = ~n5791 & ~n5792_1;
  assign n1108_1 = ~n5155 & ~n5793;
  assign n5795 = ~Pg35 & ~Ng2941;
  assign n5796 = Pg35 & n4850;
  assign n5797_1 = n4842 & n5796;
  assign n5798 = n4891_1 & ~n4895;
  assign n5799 = n4879 & ~n4887;
  assign n5800 = ~Ng2955 & n5799;
  assign n5801 = n5798 & n5800;
  assign n5802_1 = n4799 & ~n4809;
  assign n5803 = ~Ng2946 & n5802_1;
  assign n5804 = n5801 & n5803;
  assign n5805 = n5797_1 & n5804;
  assign n1113_1 = ~n5795 & ~n5805;
  assign n5807_1 = Pg8719 & Ng376;
  assign n5808 = Ng385 & n5807_1;
  assign n5809 = ~Pg35 & Ng385;
  assign n1118_1 = n5808 | n5809;
  assign n5811 = ~Ng1183 & Pg13259;
  assign n5812 = ~Ng1171 & n5811;
  assign n5813 = Pg35 & ~n5812;
  assign n5814 = Ng1099 & n5813;
  assign n5815 = Ng1152 & ~n5813;
  assign n1123 = n5814 | n5815;
  assign n5817 = n4530 & n5547;
  assign n5818 = Pg35 & n5817;
  assign n1128 = Ng4871 & ~n5818;
  assign n5820 = ~Ng5180 & ~Ng5188;
  assign n5821 = Ng5176 & n5820;
  assign n5822_1 = n5018 & n5821;
  assign n5823 = ~Pg35 & ~Ng5256;
  assign n5824 = ~n5822_1 & ~n5823;
  assign n5825 = Pg35 & ~n5821;
  assign n5826_1 = ~Ng5204 & n5825;
  assign n1133_1 = n5824 & ~n5826_1;
  assign n5828 = Ng3530 & ~Ng3522;
  assign n5829 = n5634 & n5828;
  assign n5830 = n5018 & n5829;
  assign n5831 = ~Pg35 & ~Ng3590;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = Pg35 & ~n5829;
  assign n5834_1 = ~Ng3606 & n5833;
  assign n1141_1 = n5832 & ~n5834_1;
  assign n5836 = Pg35 & n5297;
  assign n5837 = Ng1917 & n5836;
  assign n5838 = Pg35 & ~n5297;
  assign n5839_1 = Ng1926 & n5838;
  assign n5840 = ~n5837 & ~n5839_1;
  assign n5841 = n4653 & n5297;
  assign n5842 = Pg35 & n4928;
  assign n5843 = Ng110 & n5842;
  assign n5844 = n5841 & n5843;
  assign n5845 = ~Pg35 & Ng1932;
  assign n5846 = ~n5844 & ~n5845;
  assign n1146_1 = ~n5840 | ~n5846;
  assign n5848 = ~Pg35 & Ng6209;
  assign n5849 = Ng6209 & Ng6203;
  assign n5850 = n5111 & n5849;
  assign n1151_1 = n5848 | n5850;
  assign n5852 = ~Pg35 & ~Ng3570;
  assign n5853 = n5032_1 & n5201;
  assign n5854 = Pg35 & ~Ng3586;
  assign n5855 = ~n5853 & n5854;
  assign n5856_1 = n5018 & n5853;
  assign n5857 = ~n5855 & ~n5856_1;
  assign n1156_1 = ~n5852 & n5857;
  assign n5859 = ~Pg35 & Ng287;
  assign n5860 = Ng291 & n5713;
  assign n5861 = ~n5710 & ~n5860;
  assign n5862 = ~n5711_1 & ~n5861;
  assign n1161 = n5859 | n5862;
  assign n5864 = Pg35 & n5548;
  assign n1166_1 = Ng4646 & ~n5864;
  assign n5866 = n5032_1 & n5200;
  assign n5867 = n5018 & n5866;
  assign n5868 = ~Pg35 & ~Ng3542;
  assign n5869 = ~n5867 & ~n5868;
  assign n5870 = Pg35 & ~n5866;
  assign n5871 = ~Ng3570 & n5870;
  assign n1171 = n5869 & ~n5871;
  assign n5873 = Pg35 & n4950;
  assign n5874 = Ng1862 & n5873;
  assign n5875 = n4579_1 & n5089;
  assign n5876 = Pg35 & ~n5875;
  assign n5877 = ~Ng1936 & n5876;
  assign n5878 = ~n5874 & ~n5877;
  assign n5879 = ~Ng1906 & ~n4950;
  assign n5880 = ~Ng1862 & ~n5879;
  assign n1182_1 = ~n5878 & ~n5880;
  assign n5882 = Ng499 & n5354;
  assign n5883 = n4574 & n5882;
  assign n5884 = n5150 & n5883;
  assign n5885 = Ng671 & n5884;
  assign n5886 = ~n5122 & ~n5124;
  assign n5887 = Ng661 & Ng728;
  assign n5888 = ~Ng661 & ~Ng728;
  assign n5889_1 = ~n5887 & ~n5888;
  assign n5890 = Ng681 & ~Ng645;
  assign n5891 = ~Ng650 & Ng699;
  assign n5892 = n5890 & n5891;
  assign n5893 = ~n5889_1 & n5892;
  assign n5894 = ~n5886 & n5893;
  assign n5895 = n5884 & n5894;
  assign n5896 = Ng703 & ~n5895;
  assign n5897 = n5885 & n5896;
  assign n5898 = ~Ng676 & n5897;
  assign n5899_1 = Pg35 & n5896;
  assign n5900 = ~n5885 & n5899_1;
  assign n5901 = Ng676 & n5900;
  assign n5902 = ~Pg35 & Ng671;
  assign n5903 = ~n5901 & ~n5902;
  assign n1187_1 = n5898 | ~n5903;
  assign n5905 = Ng847 & n5150;
  assign n5906 = Ng843 & n5905;
  assign n5907 = ~Ng843 & ~n5905;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909_1 = Pg35 & ~n5908;
  assign n1192_1 = Ng837 & ~n5909_1;
  assign n5911 = ~n5309 & ~n5565;
  assign n5912 = Pg35 & n5911;
  assign n5913 = Ng4332 & n5912;
  assign n5914_1 = Ng4311 & n5563;
  assign n5915 = n5911 & n5914_1;
  assign n5916 = Pg35 & ~n5915;
  assign n5917 = Ng4322 & ~n5916;
  assign n1197_1 = n5913 | n5917;
  assign n5919 = ~Pg115 & Pg114;
  assign n5920 = Pg115 & ~Pg114;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = ~Ng4157 & n5921;
  assign n5923 = Pg126 & ~Pg120;
  assign n5924 = ~Pg126 & Pg120;
  assign n5925 = ~Ng4146 & ~n5924;
  assign n5926 = ~n5923 & n5925;
  assign n5927 = ~n5922 & ~n5926;
  assign n5928 = Pg35 & n5927;
  assign n5929_1 = ~Pg35 & ~Ng4122;
  assign n1202 = ~n5928 & ~n5929_1;
  assign n5931 = Pg35 & n5385;
  assign n5932 = Ng93 & n4928;
  assign n5933 = n4498 & n5932;
  assign n5934_1 = n4534 & n5933;
  assign n5935 = ~n4547 & ~n5934_1;
  assign n5936 = n5931 & ~n5935;
  assign n5937 = Pg35 & ~n5385;
  assign n5938 = Ng6395 & ~n5937;
  assign n5939 = Pg35 & Ng6336;
  assign n5940 = ~n5938 & ~n5939;
  assign n1210 = ~n5936 & ~n5940;
  assign n5942_1 = ~Pg35 & Ng617;
  assign n5943 = Ng613 & n5757;
  assign n5944 = Ng617 & n5943;
  assign n5945 = Ng622 & n5944;
  assign n5946 = Ng622 & n5737;
  assign n5947 = ~n5944 & ~n5946;
  assign n5948 = ~n5945 & ~n5947;
  assign n1215_1 = n5942_1 | n5948;
  assign n5950 = ~Ng3518 & n5205;
  assign n1220_1 = ~Ng3506 & n5950;
  assign n5952 = ~Pg35 & Ng4555;
  assign n5953 = Pg6748 & Pg35;
  assign n1225 = n5952 | n5953;
  assign n5955 = Pg35 & ~n4731;
  assign n5956 = Ng3111 & n5955;
  assign n5957 = Ng3147 & ~n5955;
  assign n1233_1 = n5956 | n5957;
  assign n5959 = n4662 & n5002;
  assign n5960 = Ng2819 & n5327;
  assign n5961 = ~Ng2719 & Ng2715;
  assign n5962 = Ng2807 & n5961;
  assign n5963 = ~n5960 & ~n5962;
  assign n5964 = Ng2803 & n5256;
  assign n5965 = Ng2815 & n5001;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967_1 = n5963 & n5966;
  assign n5968 = n5959 & ~n5967_1;
  assign n5969 = ~Ng2236 & n5256;
  assign n5970 = ~Ng2638 & n5327;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972_1 = ~Ng2370 & n5961;
  assign n5973 = ~Ng2504 & n5001;
  assign n5974 = ~n5972_1 & ~n5973;
  assign n5975 = n5971 & n5974;
  assign n5976_1 = ~n5959 & ~n5975;
  assign n5977 = Pg35 & ~n5976_1;
  assign n5978 = ~n5968 & n5977;
  assign n5979 = ~Pg35 & Ng2834;
  assign n1238_1 = n5978 | n5979;
  assign n1243_1 = Pg125 & Pg35;
  assign n5982 = ~Ng939 & ~Ng933;
  assign n5983 = Pg35 & n5982;
  assign n5984 = ~Pg35 & ~Ng952;
  assign n1248_1 = ~n5983 & ~n5984;
  assign n5986 = Pg35 & ~n5706;
  assign n1253_1 = ~n5697 & n5986;
  assign n5988 = ~Pg35 & Ng4489;
  assign n5989 = Pg6750 & Pg35;
  assign n1258_1 = n5988 | n5989;
  assign n1263_1 = Ng4836 & ~n5818;
  assign n5992 = ~Ng1030 & n5616;
  assign n5993 = Pg35 & n5992;
  assign n5994 = ~n5624_1 & ~n5993;
  assign n5995 = Ng1036 & ~n5994;
  assign n5996 = ~Ng1036 & n5616;
  assign n5997 = Pg35 & ~n5996;
  assign n5998 = Ng1030 & ~n5624_1;
  assign n5999 = ~n5997 & n5998;
  assign n1268_1 = n5995 | n5999;
  assign n6001 = ~Ng5297 & ~Ng5357;
  assign n6002 = Pg14662 & n6001;
  assign n6003 = Ng5236 & n6002;
  assign n6004 = \[4415]  & ~Pg12238;
  assign n6005 = ~\[4415]  & Pg12238;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = Ng5297 & ~Ng5357;
  assign n6008 = Ng5268 & Pg17519;
  assign n6009_1 = n6007 & n6008;
  assign n6010 = ~n6006 & ~n6009_1;
  assign n6011 = ~Ng5297 & Ng5357;
  assign n6012 = Ng5252 & n6011;
  assign n6013 = Pg17674 & n6012;
  assign n6014 = n6010 & ~n6013;
  assign n6015 = ~n6003 & n6014;
  assign n6016 = Pg14662 & Ng5228;
  assign n6017 = n6007 & n6016;
  assign n6018_1 = Ng5244 & Pg31860;
  assign n6019 = Pg17674 & n6018_1;
  assign n6020 = Pg17519 & Ng5260;
  assign n6021 = n6001 & n6020;
  assign n6022 = n6006 & ~n6021;
  assign n6023 = ~n6019 & n6022;
  assign n6024 = ~n6017 & n6023;
  assign n6025 = ~n6015 & ~n6024;
  assign n6026 = Pg17639 & Pg31860;
  assign n6027 = Ng5256 & n6026;
  assign n6028_1 = Pg13039 & Ng5196;
  assign n6029 = Ng5204 & Ng5339;
  assign n6030 = ~n6028_1 & ~n6029;
  assign n6031 = n6001 & ~n6030;
  assign n6032 = ~n6027 & ~n6031;
  assign n6033 = Pg17787 & Ng5224;
  assign n6034 = Pg12238 & Ng5200;
  assign n6035 = ~n6033 & ~n6034;
  assign n6036 = n6011 & ~n6035;
  assign n6037 = \[4415]  & ~n6036;
  assign n6038_1 = Ng5240 & n6007;
  assign n6039 = Pg14597 & n6038_1;
  assign n6040 = n6037 & ~n6039;
  assign n6041 = n6032 & n6040;
  assign n6042 = Ng5248 & n6001;
  assign n6043 = Pg14597 & n6042;
  assign n6044 = Ng5264 & Pg17639;
  assign n6045 = Pg17577 & Ng5212;
  assign n6046 = ~n6044 & ~n6045;
  assign n6047 = n6011 & ~n6046;
  assign n6048 = ~\[4415]  & ~n6047;
  assign n6049 = Ng5232 & Pg17787;
  assign n6050 = Pg12238 & Ng5216;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = Pg31860 & ~n6051;
  assign n6053_1 = Ng5208 & Pg13039;
  assign n6054 = Ng5339 & Ng5220;
  assign n6055 = ~n6053_1 & ~n6054;
  assign n6056 = n6007 & ~n6055;
  assign n6057 = ~n6052 & ~n6056;
  assign n6058 = n6048 & n6057;
  assign n6059 = ~n6043 & n6058;
  assign n6060 = ~n6041 & ~n6059;
  assign n6061 = ~n6025 & ~n6060;
  assign n6062 = ~Ng5272 & n6061;
  assign n6063 = \[4415]  & Pg31860;
  assign n6064 = Pg17577 & n6063;
  assign n6065 = n6061 & ~n6064;
  assign n6066 = Pg33959 & ~n6065;
  assign n6067_1 = Pg35 & n6066;
  assign n6068 = ~n6062 & n6067_1;
  assign n6069 = Pg35 & ~Pg33959;
  assign n6070 = \[4427]  & n6069;
  assign n6071 = ~Pg35 & Ng5272;
  assign n6072 = ~n6070 & ~n6071;
  assign n1273_1 = n6068 | ~n6072;
  assign n6074 = ~Pg35 & ~Ng1183;
  assign n6075 = ~Ng996 & Pg7916;
  assign n6076 = Pg35 & n6075;
  assign n6077 = Pg35 & ~Pg7916;
  assign n6078 = ~Ng1178 & n6077;
  assign n6079 = ~n6076 & ~n6078;
  assign n1278_1 = ~n6074 & n6079;
  assign n6081 = Ng3179 & ~Ng3171;
  assign n6082 = n5015 & n6081;
  assign n6083 = Pg35 & ~n6082;
  assign n6084 = ~Pg35 & ~Ng3223;
  assign n6085 = ~n5018 & ~n6084;
  assign n6086 = ~n6083 & ~n6085;
  assign n6087_1 = ~Ng3239 & n6083;
  assign n1283_1 = ~n6086 & ~n6087_1;
  assign n6089 = Ng417 & ~Ng424;
  assign n6090 = ~Ng411 & n6089;
  assign n6091 = ~Ng691 & ~n6090;
  assign n6092 = Ng691 & ~n5116;
  assign n6093 = n5026 & ~n6092;
  assign n6094 = ~n6091 & n6093;
  assign n6095 = Pg35 & ~n6094;
  assign n6096 = Ng718 & n6095;
  assign n6097 = Ng655 & ~n6095;
  assign n1288_1 = n6096 | n6097;
  assign n6099 = Ng6195 & ~n4724;
  assign n6100 = n5018 & n6099;
  assign n6101_1 = n5083 & ~n6099;
  assign n1293_1 = n6100 | n6101_1;
  assign n6103 = ~Pg35 & Ng1094;
  assign n6104 = Ng1099 & ~Ng1152;
  assign n6105 = Ng1171 & n5811;
  assign n6106 = Ng1094 & n6105;
  assign n6107 = n6104 & n6106;
  assign n6108 = Ng1135 & n6107;
  assign n6109 = Pg35 & Ng1135;
  assign n6110_1 = ~n6107 & ~n6109;
  assign n6111 = ~n6108 & ~n6110_1;
  assign n1298_1 = n6103 | n6111;
  assign n6113 = ~Pg35 & Ng6390;
  assign n6114 = n5931 & ~n5934_1;
  assign n6115 = ~Ng6395 & ~n6114;
  assign n6116 = ~n5938 & ~n6115;
  assign n1303_1 = n6113 | n6116;
  assign n6118 = ~Pg35 & Ng5339;
  assign n6119 = Pg12238 & Pg14662;
  assign n6120 = Pg17519 & n6119;
  assign n6121 = Pg17674 & n6120;
  assign n6122 = ~\[4415]  & ~n6121;
  assign n6123 = \[4415]  & n6121;
  assign n6124 = Pg35 & ~n6123;
  assign n6125 = ~n6122 & n6124;
  assign n1308_1 = n6118 | n6125;
  assign n6127 = Ng554 & n5145;
  assign n6128 = ~Pg35 & Ng807;
  assign n6129 = ~n5144 & ~n6128;
  assign n1313_1 = n6127 | ~n6129;
  assign n6131 = ~Ng269 & n5182;
  assign n6132 = Pg73 & ~Ng255;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = Pg73 & Pg72;
  assign n6135 = Pg72 & ~Ng262;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = Pg35 & n6136;
  assign n6138_1 = n6133 & n6137;
  assign n6139 = ~Pg35 & \[4432] ;
  assign n1318_1 = n6138_1 | n6139;
  assign n1323_1 = Pg35 & Ng3853;
  assign n6142 = Pg33959 & n6064;
  assign n6143_1 = Pg35 & ~n6142;
  assign n6144 = Ng5134 & n6143_1;
  assign n6145 = Ng5128 & ~n6143_1;
  assign n1328_1 = n6144 | n6145;
  assign n1336_1 = Pg35 & Ng3881;
  assign n6148_1 = ~Pg35 & Ng2491;
  assign n6149 = Pg35 & ~n5007;
  assign n6150 = Ng2485 & n6149;
  assign n6151 = ~n6148_1 & ~n6150;
  assign n6152 = n4648 & n5007;
  assign n6153_1 = n5843 & n6152;
  assign n6154 = Pg35 & n5007;
  assign n6155 = Ng2476 & n6154;
  assign n6156 = ~n6153_1 & ~n6155;
  assign n1340 = ~n6151 | ~n6156;
  assign n6158 = ~Pg35 & Ng918;
  assign n6159 = Ng921 & Ng904;
  assign n6160 = Pg12919 & n6159;
  assign n6161_1 = Ng936 & n6160;
  assign n6162 = Ng907 & n6161_1;
  assign n6163 = Ng911 & n6162;
  assign n6164 = Ng914 & n6163;
  assign n6165 = Ng918 & n6164;
  assign n6166_1 = Ng925 & n6165;
  assign n6167 = Pg35 & Pg12919;
  assign n6168 = Ng925 & n6167;
  assign n6169 = ~n6165 & ~n6168;
  assign n6170_1 = ~n6166_1 & ~n6169;
  assign n1345_1 = n6158 | n6170_1;
  assign n6172 = Ng5535 & ~Ng5527;
  assign n6173 = ~Ng5511 & ~Ng5517;
  assign n6174 = ~Ng5523 & n6173;
  assign n6175_1 = n6172 & n6174;
  assign n6176 = n5083 & n6175_1;
  assign n6177 = ~Pg35 & Ng5559;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = Pg35 & Ng5555;
  assign n6180_1 = ~n6175_1 & n6179;
  assign n1355_1 = ~n6178 | n6180_1;
  assign n6182 = ~Pg35 & Ng1783;
  assign n6183 = Ng2775 & n4764;
  assign n6184_1 = n5004 & n5961;
  assign n6185 = ~n6183 & n6184_1;
  assign n6186 = n4658_1 & n6185;
  assign n6187 = n4928 & n6186;
  assign n6188 = ~Ng1783 & Ng1792;
  assign n6189_1 = ~Ng110 & n6188;
  assign n6190 = Ng110 & ~n6188;
  assign n6191 = ~n6189_1 & ~n6190;
  assign n6192 = n6187 & n6191;
  assign n6193_1 = ~Ng1798 & ~n6187;
  assign n6194 = Pg35 & ~n6193_1;
  assign n6195 = ~n6192 & n6194;
  assign n1363_1 = n6182 | n6195;
  assign n6197_1 = Pg35 & ~Ng2841;
  assign n6198 = ~Pg35 & Ng4082;
  assign n6199 = ~n6197_1 & ~n6198;
  assign n6200 = Ng4064 & Ng4057;
  assign n6201 = Ng4141 & n6200;
  assign n6202_1 = Ng4082 & n6201;
  assign n6203 = Ng4076 & n6202_1;
  assign n6204 = Pg35 & Ng4076;
  assign n6205 = ~n6202_1 & ~n6204;
  assign n6206 = ~n6203 & ~n6205;
  assign n1368_1 = ~n6199 | n6206;
  assign n6208 = ~Pg35 & ~Ng2927;
  assign n6209 = Pg35 & ~Ng4072;
  assign n6210 = ~Ng4153 & ~Ng2941;
  assign n6211 = n6209 & n6210;
  assign n1373_1 = ~n6208 & ~n6211;
  assign n6213 = Ng3873 & Ng3869;
  assign n6214 = ~Ng3881 & n6213;
  assign n6215 = n5018 & n6214;
  assign n6216 = ~Pg35 & ~Ng3953;
  assign n6217_1 = ~n6215 & ~n6216;
  assign n6218 = Pg35 & ~n6214;
  assign n6219 = ~Ng3905 & n6218;
  assign n1378_1 = n6217_1 & ~n6219;
  assign n6221 = ~Pg35 & Ng758;
  assign n6222_1 = Ng763 & n5145;
  assign n6223 = ~n5135 & ~n6222_1;
  assign n6224 = ~n5136 & ~n6223;
  assign n1383_1 = n6221 | n6224;
  assign n6226 = ~Ng6215 & ~Ng6203;
  assign n6227_1 = ~Ng6209 & n6226;
  assign n6228 = n4723 & n6227_1;
  assign n6229 = n5018 & n6228;
  assign n6230 = ~Pg35 & ~Ng6259;
  assign n6231_1 = ~n6229 & ~n6230;
  assign n6232 = Pg35 & ~n6228;
  assign n6233 = ~Ng6255 & n6232;
  assign n1388_1 = n6231_1 & ~n6233;
  assign n4588_1 = Pg35 & Ng4423;
  assign n6236_1 = ~Pg35 & Ng4427;
  assign n1393_1 = n4588_1 | n6236_1;
  assign n1398_1 = Ng4864 & ~n5818;
  assign n6239 = Pg35 & Ng4722;
  assign n6240 = ~Pg35 & Ng4717;
  assign n1403_1 = n6239 | n6240;
  assign n6242 = ~Pg35 & Ng582;
  assign n6243 = Ng590 & n5737;
  assign n6244 = ~n5752 & ~n6243;
  assign n6245 = ~n5753 & ~n6244;
  assign n1408_1 = n6242 | n6245;
  assign n6247 = ~Pg35 & ~Ng1612;
  assign n6248 = Ng2771 & n4764;
  assign n6249 = n5257 & ~n6248;
  assign n6250 = ~Ng1657 & n6249;
  assign n6251 = Ng1648 & n6250;
  assign n6252 = Ng1632 & ~n6251;
  assign n6253 = ~Ng1592 & Ng1636;
  assign n6254 = n6251 & ~n6253;
  assign n6255 = Pg35 & ~n6254;
  assign n6256 = ~n6252 & n6255;
  assign n1416_1 = ~n6247 & ~n6256;
  assign n6258 = ~Pg14662 & ~Pg17674;
  assign n6259 = ~n6119 & ~n6258;
  assign n6260 = Pg35 & ~Pg13039;
  assign n6261 = ~Pg17577 & ~Pg17519;
  assign n6262 = n6260 & n6261;
  assign n1421_1 = ~n6259 & n6262;
  assign n6264 = Pg13272 & ~Ng1526;
  assign n6265 = ~Ng1514 & n6264;
  assign n6266_1 = Pg35 & ~n6265;
  assign n6267 = Ng1495 & n6266_1;
  assign n6268 = Ng1489 & ~n6266_1;
  assign n1429_1 = n6267 | n6268;
  assign n6270 = Ng1514 & n6264;
  assign n6271_1 = ~Ng1319 & n4823;
  assign n6272 = ~Ng1478 & n6271_1;
  assign n6273 = Ng1478 & ~n6271_1;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = n6270 & n6274;
  assign n6276_1 = ~Ng1442 & ~Ng1489;
  assign n6277 = n6270 & n6276_1;
  assign n6278 = ~Ng1437 & ~n6277;
  assign n6279 = Pg35 & ~n6278;
  assign n6280_1 = ~n6275 & n6279;
  assign n6281 = ~Pg35 & Ng1442;
  assign n1434 = n6280_1 | n6281;
  assign n6283 = ~Pg35 & Ng6159;
  assign n6284 = Ng6336 & ~Ng6395;
  assign n6285_1 = Ng6307 & Pg17649;
  assign n6286 = n6284 & n6285_1;
  assign n6287 = Pg12422 & ~Ng6381;
  assign n6288 = ~Pg12422 & Ng6381;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~Ng6336 & Ng6395;
  assign n6291 = Ng6291 & Pg17760;
  assign n6292 = n6290 & n6291;
  assign n6293 = ~n6289 & ~n6292;
  assign n6294_1 = ~Ng6336 & ~Ng6395;
  assign n6295 = Ng6275 & n6294_1;
  assign n6296 = Pg14779 & n6295;
  assign n6297 = n6293 & ~n6296;
  assign n6298_1 = ~n6286 & n6297;
  assign n6299 = Pg17649 & Ng6299;
  assign n6300 = n6294_1 & n6299;
  assign n6301 = Pg17760 & Ng6283;
  assign n6302 = n4547 & n6301;
  assign n6303_1 = n6289 & ~n6302;
  assign n6304 = Pg14779 & n6284;
  assign n6305 = Ng6267 & n6304;
  assign n6306 = n6303_1 & ~n6305;
  assign n6307_1 = ~n6300 & n6306;
  assign n6308 = ~n6298_1 & ~n6307_1;
  assign n6309 = Pg17743 & n4547;
  assign n6310 = Ng6295 & n6309;
  assign n6311_1 = Pg17845 & Ng6263;
  assign n6312 = Ng6239 & Pg12422;
  assign n6313 = ~n6311_1 & ~n6312;
  assign n6314 = n6290 & ~n6313;
  assign n6315 = ~n6310 & ~n6314;
  assign n6316_1 = Ng6235 & Pg13085;
  assign n6317 = Ng6377 & Ng6243;
  assign n6318 = ~n6316_1 & ~n6317;
  assign n6319 = n6294_1 & ~n6318;
  assign n6320 = Ng6381 & ~n6319;
  assign n6321_1 = Pg14705 & n6284;
  assign n6322 = Ng6279 & n6321_1;
  assign n6323 = n6320 & ~n6322;
  assign n6324 = n6315 & n6323;
  assign n6325 = Pg17743 & Ng6303;
  assign n6326_1 = Pg17685 & Ng6251;
  assign n6327 = ~n6325 & ~n6326_1;
  assign n6328 = n6290 & ~n6327;
  assign n6329 = Ng6247 & Pg13085;
  assign n6330 = Ng6377 & Ng6259;
  assign n6331_1 = ~n6329 & ~n6330;
  assign n6332 = n6284 & ~n6331_1;
  assign n6333 = ~Ng6381 & ~n6332;
  assign n6334 = Ng6271 & Pg17845;
  assign n6335 = Ng6255 & Pg12422;
  assign n6336_1 = ~n6334 & ~n6335;
  assign n6337 = n4547 & ~n6336_1;
  assign n6338 = Pg14705 & n6294_1;
  assign n6339 = Ng6287 & n6338;
  assign n6340 = ~n6337 & ~n6339;
  assign n6341 = n6333 & n6340;
  assign n6342 = ~n6328 & n6341;
  assign n6343 = ~n6324 & ~n6342;
  assign n6344 = ~n6308 & ~n6343;
  assign n6345_1 = Ng6311 & n5383;
  assign n6346 = n6344 & ~n6345_1;
  assign n6347 = n5386 & n6346;
  assign n6348 = Pg35 & Ng6154;
  assign n6349 = n5385 & ~n6344;
  assign n6350_1 = ~n5383 & n6349;
  assign n6351 = n6348 & ~n6350_1;
  assign n6352 = ~n6347 & n6351;
  assign n6353 = n5931 & ~n6346;
  assign n6354 = ~Ng6154 & n6353;
  assign n6355_1 = ~n6352 & ~n6354;
  assign n1439_1 = n6283 | ~n6355_1;
  assign n6357 = Ng5523 & n6172;
  assign n6358 = Pg35 & ~n6357;
  assign n6359 = Ng5567 & n6358;
  assign n6360_1 = ~Pg35 & Ng5611;
  assign n6361 = ~n5083 & ~n6360_1;
  assign n6362 = ~n6358 & ~n6361;
  assign n1448 = n6359 | n6362;
  assign n6364 = ~Ng1728 & Ng1772;
  assign n6365_1 = ~n5063 & n6364;
  assign n6366 = n5070 & n6365_1;
  assign n6367 = ~Pg35 & Ng1756;
  assign n6368 = Pg35 & Ng1752;
  assign n6369 = ~n6365_1 & n6368;
  assign n6370_1 = ~n6367 & ~n6369;
  assign n1453 = n6366 | ~n6370_1;
  assign n6372 = Ng1894 & ~n5838;
  assign n6373 = Ng1917 & n5838;
  assign n6374_1 = ~n5844 & ~n6373;
  assign n1458_1 = n6372 | ~n6374_1;
  assign n6376 = ~Pg35 & Ng739;
  assign n6377_1 = Ng744 & n5145;
  assign n6378 = ~n5132 & ~n6377_1;
  assign n6379 = ~n5133 & ~n6378;
  assign n1463 = n6376 | n6379;
  assign n6381_1 = Pg35 & Ng4737;
  assign n6382 = ~Pg35 & Ng4722;
  assign n1468_1 = n6381_1 | n6382;
  assign n1473 = Pg113 & Pg35;
  assign n6385 = Ng6219 & ~Ng6227;
  assign n6386 = ~Ng6209 & Ng6203;
  assign n6387 = n6385 & n6386;
  assign n6388 = n5083 & n6387;
  assign n6389 = ~Pg35 & Ng6239;
  assign n6390 = ~n6388 & ~n6389;
  assign n6391_1 = Pg35 & Ng6267;
  assign n6392 = ~n6387 & n6391_1;
  assign n1478_1 = ~n6390 | n6392;
  assign n6394 = Ng1442 & n6266_1;
  assign n6395 = Ng1495 & ~n6266_1;
  assign n1486 = n6394 | n6395;
  assign n6397 = Ng5965 & n5050;
  assign n6398 = ~Pg35 & Ng5961;
  assign n6399 = ~n5083 & ~n6398;
  assign n6400_1 = ~n5050 & ~n6399;
  assign n1491_1 = n6397 | n6400_1;
  assign n6402 = ~Pg35 & Ng1246;
  assign n6403 = ~Pg12919 & Pg17400;
  assign n6404_1 = ~Pg10500 & ~Pg17400;
  assign n6405 = Pg35 & ~n6404_1;
  assign n6406 = ~n6403 & n6405;
  assign n1501_1 = n6402 | n6406;
  assign n6408 = n5310 & n5559;
  assign n6409_1 = Pg35 & ~n6408;
  assign n1505_1 = Ng4633 & ~n6409_1;
  assign n6411 = ~Pg35 & ~Ng5248;
  assign n6412 = Ng5164 & Ng5170;
  assign n6413 = n5041 & n6412;
  assign n6414_1 = n5018 & n6413;
  assign n6415 = Pg35 & ~Ng5264;
  assign n6416 = ~n6413 & n6415;
  assign n6417 = ~n6414_1 & ~n6416;
  assign n1510_1 = ~n6411 & n6417;
  assign n6419 = Ng2587 & ~n5330;
  assign n6420 = Ng2610 & n5330;
  assign n6421 = n4633 & n5329;
  assign n6422 = n5843 & n6421;
  assign n6423_1 = ~n6420 & ~n6422;
  assign n1518_1 = n6419 | ~n6423_1;
  assign n1523_1 = Pg35 & Ng5160;
  assign n6426 = Ng5863 & ~Ng5857;
  assign n6427 = ~Ng5873 & ~Ng5881;
  assign n6428_1 = n6426 & n6427;
  assign n6429 = Pg35 & ~n6428_1;
  assign n6430 = Ng5933 & n6429;
  assign n6431 = ~Pg35 & Ng5917;
  assign n6432 = ~n5083 & ~n6431;
  assign n6433_1 = ~n6429 & ~n6432;
  assign n1528 = n6430 | n6433_1;
  assign n6435 = Ng1526 & ~Ng1514;
  assign n6436 = Pg13272 & n6435;
  assign n6437 = ~Ng1448 & n6271_1;
  assign n6438_1 = Ng1448 & ~n6271_1;
  assign n6439 = ~n6437 & ~n6438_1;
  assign n6440 = n6436 & n6439;
  assign n6441 = n6276_1 & n6436;
  assign n6442 = ~Ng1454 & ~n6441;
  assign n6443_1 = Pg35 & ~n6442;
  assign n6444 = ~n6440 & n6443_1;
  assign n6445 = ~Pg35 & Ng1478;
  assign n1533_1 = n6444 | n6445;
  assign n6447 = Pg35 & ~n5120;
  assign n6448_1 = Ng753 & n6447;
  assign n6449 = Ng732 & ~n6447;
  assign n1538 = n6448_1 | n6449;
  assign n6451 = ~Pg35 & ~Ng1291;
  assign n6452 = Pg35 & Ng1306;
  assign n6453_1 = ~Ng1296 & n6452;
  assign n1543_1 = ~n6451 & ~n6453_1;
  assign n1548_1 = Pg35 & Ng3151;
  assign n6456 = ~Ng2980 & ~Ng55;
  assign n6457 = Pg35 & n6456;
  assign n6458_1 = ~Pg35 & ~Ng2886;
  assign n1553 = ~n6457 & ~n6458_1;
  assign n6460 = ~Pg35 & Ng6723;
  assign n6461 = Pg14828 & Pg12470;
  assign n6462 = Pg17778 & n6461;
  assign n6463_1 = Pg17688 & n6462;
  assign n6464 = ~Ng6727 & ~n6463_1;
  assign n6465 = Ng6727 & n6463_1;
  assign n6466 = Pg35 & ~n6465;
  assign n6467 = ~n6464 & n6466;
  assign n1558_1 = n6460 | n6467;
  assign n6469 = ~Pg35 & Ng3522;
  assign n4157_1 = Pg35 & Ng3530;
  assign n6471 = ~n5095 & ~n4157_1;
  assign n6472 = ~n4706 & ~n6471;
  assign n6473_1 = ~n5204 & n6472;
  assign n1563_1 = n6469 | n6473_1;
  assign n6475 = Pg35 & Ng4104;
  assign n6476 = Ng4087 & n6203;
  assign n6477 = Ng4093 & n6476;
  assign n6478_1 = Ng4098 & n6477;
  assign n6479 = Pg35 & ~n6478_1;
  assign n6480 = Ng4108 & ~n6479;
  assign n6481 = n6475 & ~n6480;
  assign n6482 = ~n6475 & n6480;
  assign n6483_1 = ~n6481 & ~n6482;
  assign n1568 = n6197_1 | ~n6483_1;
  assign n6485 = ~Pg35 & Ng1306;
  assign n6486 = Pg7946 & ~Ng1521;
  assign n6487 = ~Pg7946 & ~Ng1532;
  assign n6488_1 = Pg35 & ~n6487;
  assign n6489 = ~n6486 & n6488_1;
  assign n1573 = n6485 | n6489;
  assign n1578_1 = Pg35 & ~Ng4308;
  assign n6492 = Ng1514 & n4968;
  assign n6493_1 = ~Ng1526 & n6492;
  assign n6494 = Pg17320 & ~n6493_1;
  assign n6495 = ~n4287 & ~n4973;
  assign n6496 = ~Ng2704 & n4975;
  assign n6497 = n6495 & ~n6496;
  assign n6498_1 = ~n6494 & n6497;
  assign n6499 = ~Ng2153 & Ng2197;
  assign n6500 = ~n6498_1 & n6499;
  assign n6501 = Ng1585 & ~n6496;
  assign n6502 = Ng4180 & n6495;
  assign n6503_1 = ~n6497 & ~n6502;
  assign n6504 = ~n6501 & ~n6503_1;
  assign n6505 = Pg35 & ~n6504;
  assign n6506 = n6500 & n6505;
  assign n6507 = ~Pg35 & Ng2181;
  assign n6508_1 = Ng2177 & ~n6500;
  assign n6509 = Pg35 & n6508_1;
  assign n6510 = ~n6507 & ~n6509;
  assign n1582_1 = n6506 | ~n6510;
  assign n6512 = n4615 & n4747;
  assign n6513_1 = Ng101 & n5669;
  assign n6514 = n6512 & ~n6513_1;
  assign n6515 = Pg35 & ~n6514;
  assign n6516 = ~Ng4760 & ~n6515;
  assign n6517 = ~Ng4754 & ~n6512;
  assign n6518_1 = ~n5669 & ~n6517;
  assign n6519 = Pg35 & ~n6513_1;
  assign n6520 = ~n6518_1 & n6519;
  assign n1592_1 = ~n6516 & ~n6520;
  assign n6522 = ~Pg35 & Ng962;
  assign n6523_1 = ~Ng1178 & Pg7916;
  assign n6524 = ~Ng1189 & ~Pg7916;
  assign n6525 = Pg35 & ~n6524;
  assign n6526 = ~n6523_1 & n6525;
  assign n1597_1 = n6522 | n6526;
  assign n6528 = Pg35 & n4978;
  assign n6529 = Ng2287 & n6528;
  assign n6530 = ~Ng2287 & ~n5576;
  assign n6531 = n4586 & n5089;
  assign n6532_1 = Pg35 & ~n6531;
  assign n6533 = ~Ng2361 & n6532_1;
  assign n6534 = ~n6530 & n6533;
  assign n1602_1 = n6529 | n6534;
  assign n6536 = Ng4269 & Ng4258;
  assign n6537_1 = Ng4264 & n6536;
  assign n6538 = Pg35 & Ng4273;
  assign n6539 = ~n6537_1 & n6538;
  assign n6540 = Ng4264 & ~Ng4273;
  assign n6541 = Pg35 & ~n6540;
  assign n6542_1 = Ng4269 & ~n5687_1;
  assign n6543 = ~n6541 & n6542_1;
  assign n1607_1 = n6539 | n6543;
  assign n6545 = ~Pg35 & Ng1384;
  assign n6546 = ~Ng1389 & ~n5587;
  assign n6547_1 = Pg35 & Ng1351;
  assign n6548 = ~Ng1389 & n6547_1;
  assign n6549 = ~n5588 & ~n6548;
  assign n6550 = ~n6546 & ~n6549;
  assign n1612_1 = n6545 | n6550;
  assign n6552_1 = Ng1700 & n5247;
  assign n6553 = Ng1706 & ~n5247;
  assign n1617_1 = n6552_1 | n6553;
  assign n6555 = n4677 & n4745;
  assign n6556_1 = Ng4681 & ~n6555;
  assign n6557 = Pg17646 & Ng6035;
  assign n6558 = n4551 & n6557;
  assign n6559 = n6556_1 & n6558;
  assign n6560 = Pg35 & ~n6559;
  assign n6561_1 = ~Ng5835 & n6560;
  assign n6562 = Pg35 & ~Ng5835;
  assign n6563 = ~Pg35 & Ng5831;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = ~n6560 & n6564;
  assign n1622_1 = ~n6561_1 & ~n6565;
  assign n6567 = Ng1178 & Ng996;
  assign n6568 = ~Ng1189 & n6567;
  assign n6569 = Ng1024 & Ng1002;
  assign n6570 = Ng1036 & n6569;
  assign n6571_1 = ~n5609 & n6570;
  assign n6572 = n4824 & ~n6571_1;
  assign n6573 = Pg7916 & ~n6572;
  assign n6574 = n6568 & n6573;
  assign n6575 = ~Ng1171 & Ng1183;
  assign n6576_1 = Ng1193 & ~n6575;
  assign n6577 = n6574 & ~n6576_1;
  assign n6578 = Pg35 & n6577;
  assign n6579 = Ng1171 & Pg7916;
  assign n6580 = ~Ng1171 & ~Pg7916;
  assign n6581_1 = Pg35 & ~n6580;
  assign n6582 = ~n6579 & n6581_1;
  assign n1627_1 = n6578 | n6582;
  assign n6584 = Pg35 & Ng4269;
  assign n6585 = ~n5645 & ~n6584;
  assign n6586_1 = n5645 & n6584;
  assign n1632_1 = ~n6585 & ~n6586_1;
  assign n6588 = Ng2399 & n4981;
  assign n6589 = Ng2393 & ~n4981;
  assign n1637 = n6588 | n6589;
  assign n6591_1 = ~Ng4983 & ~n4606;
  assign n6592 = Ng4983 & n4606;
  assign n6593 = n4606 & n4608_1;
  assign n6594 = ~n5817 & ~n6593;
  assign n6595 = Pg35 & n6594;
  assign n6596_1 = ~n6592 & n6595;
  assign n6597 = ~n6591_1 & n6596_1;
  assign n6598 = ~Pg35 & Ng4818;
  assign n1642_1 = n6597 | n6598;
  assign n6600 = n5318 & n6172;
  assign n6601_1 = n5083 & n6600;
  assign n6602 = ~Pg35 & Ng5595;
  assign n6603 = ~n6601_1 & ~n6602;
  assign n6604 = Pg35 & Ng5611;
  assign n6605 = ~n6600 & n6604;
  assign n1647_1 = ~n6603 | n6605;
  assign n6607 = Ng4983 & n6676;
  assign n6608 = Ng4927 & n4607;
  assign n6609 = ~n4683_1 & n5478;
  assign n6610 = ~n6608 & n6609;
  assign n6611_1 = ~n6607 & ~n6610;
  assign n6612 = ~Ng4966 & ~n6611_1;
  assign n6613 = Ng4907 & n4688_1;
  assign n6614 = Ng4922 & n4686;
  assign n6615 = Ng4917 & n4607;
  assign n6616_1 = ~n6614 & ~n6615;
  assign n6617 = Ng4912 & n4683_1;
  assign n6618 = n6616_1 & ~n6617;
  assign n6619 = ~n6613 & n6618;
  assign n6620 = ~n6676 & n6619;
  assign n6621_1 = n6676 & ~n6619;
  assign n6622 = ~n6620 & ~n6621_1;
  assign n6623 = n5479 & n6622;
  assign n6624 = ~Ng4864 & ~Ng4836;
  assign n6625_1 = ~Ng4871 & n6624;
  assign n6626 = ~Ng4878 & n6625_1;
  assign n6627 = ~n4609 & n6626;
  assign n6628 = ~n6623 & n6627;
  assign n6629 = ~n6612 & n6628;
  assign n6630_1 = Ng5011 & Ng4836;
  assign n6631 = Ng4864 & ~Ng3333;
  assign n6632 = ~n6630_1 & ~n6631;
  assign n6633 = Ng4871 & Ng3684;
  assign n6634 = Ng4878 & ~Ng4035;
  assign n6635_1 = ~n6633 & ~n6634;
  assign n6636 = ~n6626 & n6635_1;
  assign n6637 = n6632 & n6636;
  assign n6638 = Pg35 & ~n6637;
  assign n1655_1 = ~n6629 & n6638;
  assign n6640 = Pg35 & ~Ng3133;
  assign n6641 = Ng3139 & n6640;
  assign n6642 = ~Ng3139 & ~n6640;
  assign n6643_1 = ~n6641 & ~n6642;
  assign n6644 = ~n5955 & ~n6643_1;
  assign n6645 = ~Ng3143 & n5955;
  assign n1660_1 = ~n6644 & ~n6645;
  assign n6647_1 = ~Ng2898 & n5797_1;
  assign n6648 = ~Pg35 & ~Ng2864;
  assign n1665 = ~n6647_1 & ~n6648;
  assign n6650 = ~Pg35 & Ng3338;
  assign n6651 = Pg13895 & Pg11349;
  assign n6652_1 = Pg16718 & n6651;
  assign n6653 = Pg16603 & n6652_1;
  assign n6654 = Ng3338 & n6653;
  assign n6655 = Pg35 & ~n6654;
  assign n6656 = ~Ng3347 & n6655;
  assign n1670_1 = n6650 | n6656;
  assign n6658 = ~Ng3179 & Ng3171;
  assign n6659 = n5015 & n6658;
  assign n6660 = Pg35 & ~n6659;
  assign n6661 = ~Pg35 & ~Ng3219;
  assign n6662_1 = ~n5018 & ~n6661;
  assign n6663 = ~n6660 & ~n6662_1;
  assign n6664 = ~Ng3235 & n6660;
  assign n1675_1 = ~n6663 & ~n6664;
  assign n6666_1 = Ng4578 & n5406;
  assign n6667 = Ng4540 & ~n5406;
  assign n6668 = ~n5408 & ~n6667;
  assign n1680 = n6666_1 | ~n6668;
  assign n6670 = n5200 & n5635;
  assign n6671_1 = n5083 & n6670;
  assign n6672 = ~Pg35 & Ng3538;
  assign n6673 = ~n6671_1 & ~n6672;
  assign n6674 = Pg35 & Ng3566;
  assign n6675 = ~n6670 & n6674;
  assign n1685_1 = ~n6673 | n6675;
  assign n6677 = ~Ng2988 & n5182;
  assign n6678 = Pg35 & ~n6677;
  assign n6679 = Ng4558 & Ng4564;
  assign n6680 = Ng4561 & n6679;
  assign n6681_1 = Ng4555 & n6680;
  assign n6682 = ~n6678 & ~n6681_1;
  assign n6683 = ~Ng4552 & ~n5182;
  assign n6684 = ~Ng4581 & n6683;
  assign n6685 = ~n6682 & ~n6684;
  assign n6686 = ~Pg35 & Ng4564;
  assign n1690_1 = n6685 | n6686;
  assign n6688 = n4682 & n5481;
  assign n6689 = Ng4878 & ~n6688;
  assign n6690 = ~Ng4054 & ~Ng4045;
  assign n6691 = Ng4054 & ~Ng4049;
  assign n6692 = ~n6690 & ~n6691;
  assign n6693 = Ng3990 & n6692;
  assign n6694 = ~Ng3990 & ~n6692;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = n6689 & ~n6695;
  assign n6697 = ~Ng4961 & ~n6696;
  assign n6698 = Pg35 & ~n6689;
  assign n6699 = Ng4961 & n6698;
  assign n6700 = n4609 & n4686;
  assign n6701 = Pg35 & n6700;
  assign n6702 = ~n6699 & ~n6701;
  assign n1695_1 = ~n6697 & ~n6702;
  assign n6704 = Pg35 & Ng4927;
  assign n6705 = ~Pg35 & Ng4912;
  assign n1700_1 = n6704 | n6705;
  assign n6707 = Pg35 & ~n5278;
  assign n6708 = ~Ng2259 & n6707;
  assign n6709 = Pg35 & ~Ng2259;
  assign n6710 = ~Pg35 & Ng2255;
  assign n6711 = ~n6709 & ~n6710;
  assign n6712 = ~n6707 & n6711;
  assign n1705 = ~n6708 & ~n6712;
  assign n6714 = ~Pg35 & Ng2827;
  assign n6715 = Pg35 & ~Ng2827;
  assign n6716 = ~n5842 & ~n6715;
  assign n6717 = Ng2729 & n4930;
  assign n6718 = Ng2724 & n6717;
  assign n6719 = Ng111 & n4928;
  assign n6720 = n6718 & ~n6719;
  assign n6721 = ~n6716 & n6720;
  assign n6722 = Ng2819 & ~n6718;
  assign n6723 = Pg35 & n6722;
  assign n6724 = ~n6721 & ~n6723;
  assign n1710_1 = n6714 | ~n6724;
  assign n6726 = ~Pg7257 & ~Pg7243;
  assign n6727 = ~Ng4375 & ~Ng4405;
  assign n6728 = ~Ng4411 & n6727;
  assign n6729 = n6726 & n6728;
  assign n6730 = Pg35 & Ng4392;
  assign n6731 = n6729 & n6730;
  assign n6732 = Pg35 & ~Ng4382;
  assign n6733 = Ng4375 & ~n6732;
  assign n1715_1 = n6731 | n6733;
  assign n6735 = Pg35 & Ng2852;
  assign n6736 = ~Pg35 & Ng2844;
  assign n1723 = n6735 | n6736;
  assign n6738 = Ng417 & n5151;
  assign n6739 = Pg35 & Ng385;
  assign n6740 = n5024 & n6739;
  assign n6741 = Ng370 & n6740;
  assign n6742 = Ng446 & n6741;
  assign n1728 = n6738 | n6742;
  assign n6744 = Ng681 & n6095;
  assign n6745 = Ng645 & ~n6095;
  assign n1733_1 = n6744 | n6745;
  assign n6747 = Ng437 & n5151;
  assign n6748 = Ng441 & ~n5151;
  assign n1738 = n6747 | n6748;
  assign n6750 = Pg35 & Ng347;
  assign n6751 = Pg35 & Pg7540;
  assign n6752 = ~Ng347 & ~n6751;
  assign n1743_1 = ~n6750 & ~n6752;
  assign n6754 = ~Ng5873 & Ng5881;
  assign n6755 = n5078 & n6754;
  assign n6756 = n5083 & n6755;
  assign n6757 = ~Pg35 & Ng5905;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = Pg35 & Ng5901;
  assign n6760 = ~n6755 & n6759;
  assign n1748 = ~n6758 | n6760;
  assign n6762 = ~Ng2886 & ~Ng2946;
  assign n6763 = Pg35 & n6762;
  assign n6764 = ~Pg35 & ~Ng2878;
  assign n1753_1 = ~n6763 & ~n6764;
  assign n6766 = Ng3494 & n5213;
  assign n6767 = Pg35 & ~Ng3484;
  assign n6768 = Ng3490 & ~n6767;
  assign n6769 = ~Ng3490 & n6767;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = ~n5213 & ~n6770;
  assign n1758_1 = n6766 | n6771;
  assign n6773 = n4522 & n5105;
  assign n6774 = Pg35 & ~n6773;
  assign n6775 = ~Ng5523 & n6774;
  assign n1763_1 = ~Ng5511 & n6775;
  assign n6777 = ~Pg35 & Ng3512;
  assign n6778 = n5634 & n5950;
  assign n1768_1 = n6777 | n6778;
  assign n6780 = ~Pg35 & Ng1687;
  assign n6781 = ~n5237 & ~n6780;
  assign n6782 = n5247 & n6781;
  assign n6783 = ~Ng1604 & ~n5247;
  assign n1773_1 = ~n6782 & ~n6783;
  assign n6785 = Ng5092 & Ng5084;
  assign n6786 = Pg35 & ~n6785;
  assign n6787 = ~Ng5092 & ~Ng5084;
  assign n6788 = n6786 & ~n6787;
  assign n6789 = ~Pg35 & Ng5084;
  assign n1778 = n6788 | n6789;
  assign n6791 = Pg35 & n6556_1;
  assign n6792 = ~Ng5990 & Ng6049;
  assign n6793 = Pg17739 & n6792;
  assign n6794 = Ng5945 & n6793;
  assign n6795 = ~Ng5990 & ~Ng6049;
  assign n6796 = Ng5929 & n6795;
  assign n6797 = Pg14738 & n6796;
  assign n6798 = ~n6794 & ~n6797;
  assign n6799 = Pg12350 & ~Ng6035;
  assign n6800 = ~Pg12350 & Ng6035;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = Ng5990 & ~Ng6049;
  assign n6803 = Pg17607 & Ng5961;
  assign n6804 = n6802 & n6803;
  assign n6805 = ~n6801 & ~n6804;
  assign n6806 = n6798 & n6805;
  assign n6807 = Pg14738 & Ng5921;
  assign n6808 = n6802 & n6807;
  assign n6809 = Pg17607 & Ng5953;
  assign n6810 = n6795 & n6809;
  assign n6811 = Pg17739 & Ng5937;
  assign n6812 = n4551 & n6811;
  assign n6813 = ~n6810 & ~n6812;
  assign n6814 = n6801 & n6813;
  assign n6815 = ~n6808 & n6814;
  assign n6816 = ~n6806 & ~n6815;
  assign n6817 = Ng5941 & n6795;
  assign n6818 = Pg14673 & n6817;
  assign n6819 = Pg17715 & Ng5957;
  assign n6820 = Ng5905 & Pg17646;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = n6792 & ~n6821;
  assign n6823 = ~n6818 & ~n6822;
  assign n6824 = Pg17819 & Ng5925;
  assign n6825 = Ng5909 & Pg12350;
  assign n6826 = ~n6824 & ~n6825;
  assign n6827 = n4551 & ~n6826;
  assign n6828 = Ng5901 & Pg13068;
  assign n6829 = Ng6031 & Ng5913;
  assign n6830 = ~n6828 & ~n6829;
  assign n6831 = n6802 & ~n6830;
  assign n6832 = ~Ng6035 & ~n6831;
  assign n6833 = ~n6827 & n6832;
  assign n6834 = n6823 & n6833;
  assign n6835 = Pg17715 & Ng5949;
  assign n6836 = Ng5965 & Pg17646;
  assign n6837 = ~n6835 & ~n6836;
  assign n6838 = n4551 & ~n6837;
  assign n6839 = Ng5889 & Pg13068;
  assign n6840 = Ng6031 & Ng5897;
  assign n6841 = ~n6839 & ~n6840;
  assign n6842 = n6795 & ~n6841;
  assign n6843 = Ng5917 & Pg17819;
  assign n6844 = Pg12350 & Ng5893;
  assign n6845 = ~n6843 & ~n6844;
  assign n6846 = n6792 & ~n6845;
  assign n6847 = Ng5933 & Pg14673;
  assign n6848 = n6802 & n6847;
  assign n6849 = Ng6035 & ~n6848;
  assign n6850 = ~n6846 & n6849;
  assign n6851 = ~n6842 & n6850;
  assign n6852 = ~n6838 & n6851;
  assign n6853 = ~n6834 & ~n6852;
  assign n6854 = ~n6816 & ~n6853;
  assign n6855 = n6791 & ~n6854;
  assign n6856 = Pg35 & ~n6556_1;
  assign n6857 = Ng4831 & n6856;
  assign n6858 = ~Pg35 & Ng5965;
  assign n6859 = ~n6857 & ~n6858;
  assign n1783_1 = n6855 | ~n6859;
  assign n6861 = Pg35 & ~n6729;
  assign n6862 = ~Ng4375 & Ng4382;
  assign n6863 = n6861 & n6862;
  assign n6864 = Pg35 & ~Ng4392;
  assign n6865 = n6729 & n6864;
  assign n6866 = ~Ng4417 & n6865;
  assign n6867 = Ng4375 & n6732;
  assign n6868 = ~Pg35 & Ng4388;
  assign n6869 = ~n6867 & ~n6868;
  assign n6870 = ~n6866 & n6869;
  assign n1788_1 = n6863 | ~n6870;
  assign n6872 = ~Pg35 & Ng6381;
  assign n6873 = Pg14779 & Pg12422;
  assign n6874 = Pg17649 & n6873;
  assign n6875 = Pg17760 & n6874;
  assign n6876 = Ng6381 & n6875;
  assign n6877 = Pg35 & ~n6876;
  assign n6878 = ~Ng6390 & n6877;
  assign n1793_1 = n6872 | n6878;
  assign n6880 = Ng203 & n5352;
  assign n6881 = Ng174 & Ng168;
  assign n6882 = ~Ng182 & ~n6881;
  assign n6883 = n6880 & ~n6882;
  assign n6884 = ~Ng174 & ~Ng168;
  assign n6885 = Pg35 & ~n6884;
  assign n1798_1 = n6883 & n6885;
  assign n6887 = Ng3965 & n5730;
  assign n6888 = ~Pg35 & Ng3961;
  assign n6889 = ~n5083 & ~n6888;
  assign n6890 = ~n5730 & ~n6889;
  assign n1803 = n6887 | n6890;
  assign n6892 = n4677 & n4748;
  assign n6893 = Ng4674 & ~n6892;
  assign n6894 = Pg35 & ~n6893;
  assign n6895 = Ng4749 & n6894;
  assign n6896 = ~Ng5694 & ~Ng5703;
  assign n6897 = Ng5703 & ~Ng5698;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = ~Ng5644 & ~n6898;
  assign n6900 = Ng5644 & n6898;
  assign n6901 = ~Ng4749 & ~n6900;
  assign n6902 = ~n6899 & n6901;
  assign n6903 = n4615 & n4678_1;
  assign n6904 = Pg35 & n6893;
  assign n6905 = n6903 & n6904;
  assign n6906 = ~n6902 & n6905;
  assign n1808_1 = n6895 | n6906;
  assign n6908 = ~\[4421]  & ~n5657;
  assign n6909 = Ng4180 & n5658;
  assign n6910 = ~n5659_1 & ~n6909;
  assign n6911 = ~n6908 & ~n6910;
  assign n6912 = Pg35 & ~n6911;
  assign n6913 = ~Pg35 & Ng2089;
  assign n6914 = n5664 & ~n6913;
  assign n6915 = ~n6912 & n6914;
  assign n6916 = ~Ng2008 & ~n5664;
  assign n1813_1 = ~n6915 & ~n6916;
  assign n6918 = Ng3863 & ~Ng3857;
  assign n6919 = ~Ng3873 & ~Ng3881;
  assign n6920 = n6918 & n6919;
  assign n6921 = n5018 & n6920;
  assign n6922 = ~Pg35 & ~Ng3917;
  assign n6923 = ~n6921 & ~n6922;
  assign n6924 = Pg35 & ~n6920;
  assign n6925 = ~Ng3933 & n6924;
  assign n1822 = n6923 & ~n6925;
  assign n6927 = Ng298 & n5712;
  assign n6928 = Ng142 & n6927;
  assign n6929 = Pg35 & n6928;
  assign n6930 = ~Pg35 & Ng301;
  assign n1827_1 = n6929 | n6930;
  assign n6932 = ~Ng3100 & Pg8215;
  assign n6933 = ~Ng3050 & ~n6932;
  assign n6934 = Pg35 & ~Pg8277;
  assign n6935 = ~n6933 & n6934;
  assign n6936 = ~Pg35 & Ng3100;
  assign n1832_1 = n6935 | n6936;
  assign n6938 = ~Ng990 & ~Pg19334;
  assign n6939 = ~Pg7916 & n6938;
  assign n6940 = Pg12919 & ~n6939;
  assign n6941 = Ng1052 & n6940;
  assign n6942 = ~Ng979 & ~n6941;
  assign n6943 = ~Ng1052 & ~n6940;
  assign n6944 = Pg35 & ~n6943;
  assign n1837_1 = n6942 & n6944;
  assign n6946 = Ng2787 & n4764;
  assign n6947 = n5328 & ~n6946;
  assign n6948 = Ng2060 & n6947;
  assign n6949 = Ng2028 & n6948;
  assign n6950 = Pg35 & ~n6949;
  assign n6951 = Ng2122 & n6950;
  assign n6952 = Ng2116 & ~n6950;
  assign n1845_1 = n6951 | n6952;
  assign n6954 = Ng1526 & n6492;
  assign n6955 = Pg17423 & ~n6954;
  assign n6956 = ~Ng2704 & n5530;
  assign n6957 = ~n4322 & ~n4973;
  assign n6958 = ~n6956 & n6957;
  assign n6959 = ~n6955 & n6958;
  assign n6960 = Ng2421 & ~n6959;
  assign n6961 = n4570 & n5089;
  assign n6962 = Pg35 & ~n6961;
  assign n6963 = n6960 & n6962;
  assign n6964 = ~Pg35 & Ng2472;
  assign n6965 = Pg35 & n6959;
  assign n6966 = Ng2465 & n6965;
  assign n6967 = ~n6964 & ~n6966;
  assign n1850 = n6963 | ~n6967;
  assign n6969 = ~Pg35 & ~Ng5881;
  assign n6970 = n5078 & n6427;
  assign n6971 = Pg35 & ~Ng5889;
  assign n6972 = ~n6970 & n6971;
  assign n6973 = n5018 & n6970;
  assign n6974 = ~n6972 & ~n6973;
  assign n1855_1 = ~n6969 & n6974;
  assign n6976 = Ng4572 & n5406;
  assign n6977 = Ng4480 & ~n5406;
  assign n6978 = ~n5408 & ~n6977;
  assign n1860_1 = n6976 | ~n6978;
  assign n6980 = Pg35 & ~Ng358;
  assign n1865_1 = ~Pg8719 & n6980;
  assign n6982 = Pg35 & Ng4653;
  assign n6983 = ~Ng4688 & ~n6982;
  assign n6984 = Ng4688 & n6982;
  assign n6985 = ~n6983 & ~n6984;
  assign n1869_1 = ~n5864 & n6985;
  assign n6987 = ~Pg35 & Ng3171;
  assign n6988 = Ng3167 & Ng3171;
  assign n2084_1 = Pg35 & Ng3179;
  assign n6990 = ~n6988 & ~n2084_1;
  assign n6991 = ~n4731 & ~n5251;
  assign n6992 = ~n6990 & n6991;
  assign n1874 = n6987 | n6992;
  assign n6994 = Ng1728 & n5087;
  assign n6995 = ~Ng1728 & ~n5288;
  assign n6996 = Pg35 & ~n5090;
  assign n6997 = ~Ng1802 & n6996;
  assign n6998 = ~n6995 & n6997;
  assign n1879_1 = n6994 | n6998;
  assign n7000 = Ng1585 & ~n6956;
  assign n7001 = Ng4180 & n6957;
  assign n7002 = ~n6958 & ~n7001;
  assign n7003 = ~n7000 & ~n7002;
  assign n7004 = Pg35 & ~n7003;
  assign n7005 = ~Pg35 & Ng2514;
  assign n7006 = ~n7004 & ~n7005;
  assign n7007 = ~Ng2495 & ~Ng2421;
  assign n7008 = Pg35 & ~n7007;
  assign n7009 = ~n6965 & ~n7008;
  assign n7010 = n7006 & n7009;
  assign n7011 = ~Ng2433 & ~n7009;
  assign n1884_1 = ~n7010 & ~n7011;
  assign n7013 = ~Pg35 & Ng3831;
  assign n7014 = Ng4040 & n4535;
  assign n7015 = Pg16693 & n7014;
  assign n7016 = n6689 & n7015;
  assign n7017 = Pg35 & ~n7016;
  assign n7018 = Ng3835 & n7017;
  assign n7019 = Pg35 & ~Ng3835;
  assign n7020 = n7016 & n7019;
  assign n7021 = ~n7018 & ~n7020;
  assign n1889_1 = n7013 | ~n7021;
  assign n7023 = Pg35 & ~n4724;
  assign n7024 = Ng6187 & n7023;
  assign n7025 = Ng6181 & ~n7023;
  assign n1894 = n7024 | n7025;
  assign n1899 = Pg35 & Ng4917;
  assign n7028 = ~Pg35 & Ng1199;
  assign n7029 = Pg7916 & ~n6568;
  assign n7030 = n6575 & n7029;
  assign n7031 = Ng1199 & n7030;
  assign n7032 = Pg35 & Ng1070;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = Ng1070 & n7031;
  assign n7035 = ~n6577 & ~n7034;
  assign n7036 = ~n7033 & n7035;
  assign n1904 = n7028 | n7036;
  assign n7038 = Ng817 & n5150;
  assign n7039 = Ng832 & n7038;
  assign n7040 = ~Ng822 & ~n7039;
  assign n7041 = Ng822 & n7039;
  assign n7042 = Ng847 & Ng812;
  assign n7043 = Ng847 & ~Ng837;
  assign n7044 = ~n7042 & ~n7043;
  assign n7045 = Pg35 & n7044;
  assign n7046 = ~n7041 & n7045;
  assign n7047 = ~n7040 & n7046;
  assign n7048 = ~Pg35 & Ng832;
  assign n1909_1 = n7047 | n7048;
  assign n7050 = ~Pg35 & Ng911;
  assign n7051 = Ng914 & n6167;
  assign n7052 = ~n6163 & ~n7051;
  assign n7053 = ~n6164 & ~n7052;
  assign n1917 = n7050 | n7053;
  assign n7055 = Pg35 & Ng4157;
  assign n7056 = Pg116 & n7055;
  assign n7057 = Pg114 & ~Ng4157;
  assign n7058 = Pg35 & n7057;
  assign n7059 = ~Pg35 & Ng4153;
  assign n7060 = ~n7058 & ~n7059;
  assign n1926 = n7056 | ~n7060;
  assign n7062 = ~n5606 & n5609;
  assign n7063 = Pg35 & ~n7062;
  assign n7064 = Ng969 & n7063;
  assign n7065 = Ng1046 & n5609;
  assign n7066 = n5613 & ~n7065;
  assign n7067 = ~Ng1008 & n6571_1;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = Pg35 & ~n5606;
  assign n7070 = ~n7068 & n7069;
  assign n1931_1 = n7064 | n7070;
  assign n7072 = ~Pg35 & Ng2815;
  assign n7073 = Pg35 & ~Ng2811;
  assign n7074 = ~n5842 & ~n7073;
  assign n7075 = n4766 & n4930;
  assign n7076 = ~n6719 & n7075;
  assign n7077 = ~n7074 & n7076;
  assign n7078 = Ng2807 & ~n7075;
  assign n7079 = Pg35 & n7078;
  assign n7080 = ~n7077 & ~n7079;
  assign n1936_1 = n7072 | ~n7080;
  assign n7082 = Pg35 & ~Ng4054;
  assign n7083 = n4530 & n5932;
  assign n7084 = n4534 & n7083;
  assign n7085 = n6689 & ~n7084;
  assign n7086 = n7082 & ~n7085;
  assign n7087 = ~Pg35 & Ng4049;
  assign n7088 = ~n6698 & ~n7082;
  assign n7089 = ~n7087 & n7088;
  assign n1941_1 = ~n7086 & ~n7089;
  assign n7091 = Pg35 & ~Ng6181;
  assign n7092 = Ng6187 & n7091;
  assign n7093 = ~Ng6187 & ~n7091;
  assign n7094 = ~n7092 & ~n7093;
  assign n7095 = ~n7023 & ~n7094;
  assign n7096 = ~Ng6191 & n7023;
  assign n1946 = ~n7095 & ~n7096;
  assign n7098 = Pg35 & ~Ng5069;
  assign n1951 = Ng5073 & ~n7098;
  assign n7100 = ~Pg35 & Ng5517;
  assign n7101 = n5318 & n6775;
  assign n1956_1 = n7100 | n7101;
  assign n7103 = ~Ng6549 & Ng6555;
  assign n7104 = n4713 & n7103;
  assign n7105 = n5018 & n7104;
  assign n7106 = ~Pg35 & ~Ng6621;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = Pg35 & ~n7104;
  assign n7109 = ~Ng6637 & n7108;
  assign n1965_1 = n7107 & ~n7109;
  assign n7111 = Ng174 & n5027_1;
  assign n7112 = Ng182 & ~n5027_1;
  assign n1970_1 = n7111 | n7112;
  assign n7114 = ~Pg35 & Ng1668;
  assign n7115 = ~Ng1682 & n5227;
  assign n7116 = Ng1246 & ~n5225;
  assign n7117 = ~n5235 & ~n7116;
  assign n7118 = Ng1682 & ~n5245;
  assign n7119 = n7117 & n7118;
  assign n7120 = ~n7117 & ~n7118;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = ~n5227 & n7121;
  assign n7123 = Pg35 & ~n7122;
  assign n7124 = ~n7115 & n7123;
  assign n1975_1 = n7114 | n7124;
  assign n7126 = ~Pg35 & Ng351;
  assign n7127 = ~Ng355 & ~Ng333;
  assign n7128 = Pg35 & ~Ng351;
  assign n7129 = ~n7127 & n7128;
  assign n1980_1 = n7126 | n7129;
  assign n7131 = ~Pg35 & Ng1111;
  assign n7132 = Pg13259 & n6575;
  assign n7133 = Ng1111 & n7132;
  assign n7134 = n6104 & n7133;
  assign n7135 = ~Ng1105 & n7134;
  assign n7136 = Pg35 & Ng1105;
  assign n7137 = ~n7134 & n7136;
  assign n7138 = ~n7135 & ~n7137;
  assign n1989 = n7131 | ~n7138;
  assign n7140 = Ng2807 & n4764;
  assign n7141 = n6184_1 & ~n7140;
  assign n7142 = Pg35 & ~n7141;
  assign n7143 = Ng2319 & ~n7142;
  assign n7144 = Ng2342 & n7142;
  assign n7145 = n4666 & n7141;
  assign n7146 = n5843 & n7145;
  assign n7147 = ~n7144 & ~n7146;
  assign n1994_1 = n7143 | ~n7147;
  assign n7149 = n4723 & n5849;
  assign n7150 = Pg35 & ~n7149;
  assign n7151 = Ng6307 & n7150;
  assign n7152 = ~Pg35 & Ng6291;
  assign n7153 = ~n5083 & ~n7152;
  assign n7154 = ~n7150 & ~n7153;
  assign n1999_1 = n7151 | n7154;
  assign n7156 = Ng6159 & n7023;
  assign n7157 = Ng6195 & ~n7023;
  assign n2008_1 = n7156 | n7157;
  assign n7159 = Pg35 & ~n5262;
  assign n7160 = ~n5259 & ~n7159;
  assign n7161 = ~Ng2255 & ~n7160;
  assign n7162 = Pg35 & Ng2246;
  assign n7163 = Ng2250 & n7162;
  assign n7164 = ~Ng2250 & ~n7162;
  assign n7165 = ~n7163 & ~n7164;
  assign n7166 = n7160 & ~n7165;
  assign n2013_1 = ~n7161 & ~n7166;
  assign n7168 = ~Pg35 & Ng2819;
  assign n7169 = Pg35 & ~Ng2823;
  assign n7170 = ~n5842 & ~n7169;
  assign n7171 = ~Ng2724 & n6717;
  assign n7172 = ~n6719 & n7171;
  assign n7173 = ~n7170 & n7172;
  assign n7174 = Pg35 & Ng2815;
  assign n7175 = ~n7171 & n7174;
  assign n7176 = ~n7173 & ~n7175;
  assign n2018 = n7168 | ~n7176;
  assign n7178 = ~Pg35 & Ng907;
  assign n7179 = Ng911 & n6167;
  assign n7180 = ~n6162 & ~n7179;
  assign n7181 = ~n6163 & ~n7180;
  assign n2023_1 = n7178 | n7181;
  assign n7183 = Ng1728 & ~n5063;
  assign n7184 = Ng1802 & n7183;
  assign n7185 = Pg35 & ~n7184;
  assign n7186 = Ng1748 & n7185;
  assign n7187 = ~Pg35 & Ng1752;
  assign n7188 = ~n5070 & ~n7187;
  assign n7189 = ~n7185 & ~n7188;
  assign n2036_1 = n7186 | n7189;
  assign n7191 = Ng5523 & n5374;
  assign n7192 = Pg35 & ~n7191;
  assign n7193 = ~Pg35 & ~Ng5603;
  assign n7194 = ~n5018 & ~n7193;
  assign n7195 = ~n7192 & ~n7194;
  assign n7196 = ~Ng5551 & n7192;
  assign n2041 = ~n7195 & ~n7196;
  assign n7198 = n4705 & n5034;
  assign n7199 = n5018 & n7198;
  assign n7200 = ~Pg35 & ~Ng3562;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = Pg35 & ~n7198;
  assign n7203 = ~Ng3558 & n7202;
  assign n2046_1 = n7201 & ~n7203;
  assign n7205 = Pg35 & ~n4727;
  assign n7206 = Ng5499 & n7205;
  assign n7207 = Pg35 & ~Ng5489;
  assign n7208 = ~Ng5495 & n7207;
  assign n7209 = Ng5495 & ~n7207;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = ~n7205 & ~n7210;
  assign n2051_1 = n7206 | n7211;
  assign n7213 = Pg35 & Ng2960;
  assign n7214 = ~Pg35 & Ng2950;
  assign n2056 = n7213 | n7214;
  assign n7216 = ~Ng3873 & Ng3881;
  assign n7217 = n5767 & n7216;
  assign n7218 = n5018 & n7217;
  assign n7219 = ~Pg35 & ~Ng3905;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = Pg35 & ~n7217;
  assign n7222 = ~Ng3901 & n7221;
  assign n2061 = n7220 & ~n7222;
  assign n7224 = n4610 & ~n5670;
  assign n7225 = Pg35 & ~n7224;
  assign n7226 = ~Ng4894 & ~n7225;
  assign n7227 = ~Ng4888 & ~n4610;
  assign n7228 = ~n5669 & ~n7227;
  assign n7229 = n5677 & ~n7228;
  assign n2066 = ~n7226 & ~n7229;
  assign n7231 = Ng6219 & Ng6215;
  assign n7232 = ~Ng6227 & n7231;
  assign n7233 = Pg35 & ~n7232;
  assign n7234 = Ng6251 & n7233;
  assign n7235 = ~Pg35 & Ng6299;
  assign n7236 = ~n5083 & ~n7235;
  assign n7237 = ~n7233 & ~n7236;
  assign n2071 = n7234 | n7237;
  assign n7239 = ~Pg35 & Ng1367;
  assign n7240 = ~Ng1389 & Ng1351;
  assign n7241 = n5509 & ~n7240;
  assign n7242 = Ng1373 & Ng1361;
  assign n7243 = Ng1351 & n7242;
  assign n7244 = ~n5509 & n7243;
  assign n7245 = ~Ng1312 & ~n7244;
  assign n7246 = ~n7241 & n7245;
  assign n7247 = ~Ng1345 & n7246;
  assign n7248 = ~n5506 & ~n7247;
  assign n7249 = ~Ng1361 & n7246;
  assign n7250 = n7248 & ~n7249;
  assign n7251 = ~Ng1367 & n7246;
  assign n7252 = n7250 & ~n7251;
  assign n7253 = Pg35 & ~n7252;
  assign n7254 = ~Ng1373 & n7246;
  assign n7255 = Pg35 & n7254;
  assign n7256 = ~n7253 & ~n7255;
  assign n7257 = ~Ng1373 & ~n7252;
  assign n7258 = ~n7256 & ~n7257;
  assign n2079_1 = n7239 | n7258;
  assign n7260 = ~Pg35 & Ng153;
  assign n7261 = ~Ng182 & n6884;
  assign n7262 = n6880 & ~n7261;
  assign n7263 = n5699 & ~n7262;
  assign n7264 = Ng146 & n6880;
  assign n7265 = n7263 & n7264;
  assign n7266 = Ng164 & n7265;
  assign n7267 = Ng150 & n7266;
  assign n7268 = Ng153 & n7267;
  assign n7269 = Ng157 & n7268;
  assign n7270 = Pg35 & n7263;
  assign n7271 = Ng157 & n7270;
  assign n7272 = ~n7268 & ~n7271;
  assign n7273 = ~n7269 & ~n7272;
  assign n2088_1 = n7260 | n7273;
  assign n7275 = ~Pg35 & Ng2787;
  assign n7276 = Ng2783 & ~n7171;
  assign n7277 = Pg35 & n7276;
  assign n7278 = ~n7275 & ~n7277;
  assign n7279 = Pg35 & ~Ng2791;
  assign n7280 = ~n5842 & ~n7279;
  assign n7281 = ~n4932 & n7171;
  assign n7282 = ~n7280 & n7281;
  assign n2093_1 = ~n7278 | n7282;
  assign n7284 = n5200 & n5828;
  assign n7285 = Pg35 & ~n7284;
  assign n7286 = Ng3574 & n7285;
  assign n7287 = ~Pg35 & Ng3550;
  assign n7288 = ~n5083 & ~n7287;
  assign n7289 = ~n7285 & ~n7288;
  assign n2102 = n7286 | n7289;
  assign n7291 = ~Ng2112 & ~n5664;
  assign n7292 = Pg35 & ~Ng2102;
  assign n7293 = ~Ng2108 & n7292;
  assign n7294 = Ng2108 & ~n7292;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = n5664 & n7295;
  assign n2107_1 = ~n7291 & ~n7296;
  assign n7298 = ~Ng1283 & ~Ng1277;
  assign n7299 = Pg35 & n7298;
  assign n7300 = ~Pg35 & ~Ng1296;
  assign n2112 = ~n7299 & ~n7300;
  assign n7302 = ~Pg35 & Ng437;
  assign n7303 = Ng433 & n5151;
  assign n7304 = Ng269 & n6741;
  assign n7305 = ~n7303 & ~n7304;
  assign n2117_1 = n7302 | ~n7305;
  assign n7307 = ~Pg35 & Ng749;
  assign n7308 = Ng758 & n5145;
  assign n7309 = ~n5134 & ~n7308;
  assign n7310 = ~n5135 & ~n7309;
  assign n2132 = n7307 | n7310;
  assign n2137 = ~Ng4639 & n5311;
  assign n7313 = Pg35 & ~n4714;
  assign n7314 = Pg35 & ~Ng6527;
  assign n7315 = Ng6533 & n7314;
  assign n7316 = ~Ng6533 & ~n7314;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = ~n7313 & ~n7317;
  assign n7319 = ~Ng6537 & n7313;
  assign n2142_1 = ~n7318 & ~n7319;
  assign n7321 = n5374 & n6174;
  assign n7322 = n5083 & n7321;
  assign n7323 = ~Pg35 & Ng5535;
  assign n7324 = ~n7322 & ~n7323;
  assign n7325 = Pg35 & Ng5543;
  assign n7326 = ~n7321 & n7325;
  assign n2147_1 = ~n7324 | n7326;
  assign n7328 = Ng5863 & Ng5857;
  assign n7329 = n4717 & n7328;
  assign n7330 = n5083 & n7329;
  assign n7331 = ~Pg35 & Ng5945;
  assign n7332 = ~n7330 & ~n7331;
  assign n7333 = Pg35 & Ng5961;
  assign n7334 = ~n7329 & n7333;
  assign n2155 = ~n7332 | n7334;
  assign n7336 = ~Ng6219 & ~Ng6227;
  assign n7337 = Ng6215 & n7336;
  assign n7338 = Pg35 & ~n7337;
  assign n7339 = Ng6243 & n7338;
  assign n7340 = ~Pg35 & Ng6295;
  assign n7341 = ~n5083 & ~n7340;
  assign n7342 = ~n7338 & ~n7341;
  assign n2160_1 = n7339 | n7342;
  assign n7344 = ~Pg35 & Ng626;
  assign n7345 = Ng626 & n5945;
  assign n7346 = Ng632 & n7345;
  assign n7347 = Ng632 & n5737;
  assign n7348 = ~n7345 & ~n7347;
  assign n7349 = ~n7346 & ~n7348;
  assign n2165 = n7344 | n7349;
  assign n7351 = Pg35 & \[4432] ;
  assign n7352 = ~Pg35 & Ng1211;
  assign n2170_1 = n7351 | n7352;
  assign n7354 = n5767 & n6919;
  assign n7355 = Pg35 & ~n7354;
  assign n7356 = Ng3889 & n7355;
  assign n7357 = ~Pg35 & Ng3881;
  assign n7358 = ~n5083 & ~n7357;
  assign n7359 = ~n7355 & ~n7358;
  assign n2174 = n7356 | n7359;
  assign n7361 = Pg35 & ~n5487;
  assign n7362 = Ng3476 & n7361;
  assign n7363 = Ng3470 & ~n7361;
  assign n2179 = n7362 | n7363;
  assign n7365 = n4663 & n6249;
  assign n7366 = n4928 & n7365;
  assign n7367 = Ng1664 & ~n7366;
  assign n7368 = Pg35 & n7367;
  assign n7369 = Ng1657 & ~Ng1648;
  assign n7370 = Ng110 & n7369;
  assign n7371 = ~Ng110 & ~n7369;
  assign n7372 = ~n7370 & ~n7371;
  assign n7373 = n5842 & n7372;
  assign n7374 = n7365 & n7373;
  assign n7375 = ~Pg35 & Ng1648;
  assign n7376 = ~n7374 & ~n7375;
  assign n2184 = n7368 | ~n7376;
  assign n7378 = ~Pg35 & \[4421] ;
  assign n2189 = n6167 | n7378;
  assign n7380 = ~Ng6573 & Ng6565;
  assign n7381 = n7103 & n7380;
  assign n7382 = n5083 & n7381;
  assign n7383 = ~Pg35 & Ng6613;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = Pg35 & Ng6629;
  assign n7386 = ~n7381 & n7385;
  assign n2194_1 = ~n7384 | n7386;
  assign n7388 = ~Ng862 & ~Ng896;
  assign n7389 = Ng890 & n7388;
  assign n7390 = Pg35 & n7389;
  assign n7391 = Pg14167 & n7390;
  assign n7392 = ~Pg35 & Ng269;
  assign n7393 = Pg35 & ~n7389;
  assign n7394 = Ng246 & n7393;
  assign n7395 = ~n7392 & ~n7394;
  assign n2199 = n7391 | ~n7395;
  assign n7397 = Pg35 & n4997;
  assign n2204_1 = Ng4045 & ~n7397;
  assign n7399 = Ng4438 & ~n6732;
  assign n7400 = ~Ng4452 & ~Pg7245;
  assign n7401 = ~Pg7260 & ~Ng4438;
  assign n7402 = ~Ng4443 & n7401;
  assign n7403 = n7400 & n7402;
  assign n7404 = n6730 & n7403;
  assign n2209_1 = n7399 | n7404;
  assign n7406 = Pg35 & Pg9251;
  assign n7407 = Ng4308 & ~n7406;
  assign n7408 = Pg9251 & n1578_1;
  assign n2213 = n7407 | n7408;
  assign n7410 = Ng4727 & n4613_1;
  assign n7411 = Ng4717 & n4747;
  assign n7412 = Ng4722 & n4678_1;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = Ng4732 & n4744;
  assign n7415 = n7413 & ~n7414;
  assign n7416 = ~n7410 & n7415;
  assign n7417 = ~n2499 & n7416;
  assign n7418 = n2499 & ~n7416;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = n4674 & n7419;
  assign n7421 = ~Ng4674 & ~Ng4646;
  assign n7422 = ~Ng4681 & n7421;
  assign n7423 = ~Ng4688 & n7422;
  assign n7424 = Ng4793 & n2499;
  assign n7425 = Ng4737 & n4613_1;
  assign n7426 = ~Ng4801 & ~Ng4793;
  assign n7427 = ~n4678_1 & n7426;
  assign n7428 = ~n7425 & n7427;
  assign n7429 = ~n7424 & ~n7428;
  assign n7430 = ~Ng4776 & ~n7429;
  assign n7431 = n7423 & ~n7430;
  assign n7432 = ~n7420 & n7431;
  assign n7433 = ~n4615 & n7432;
  assign n7434 = Ng4831 & Ng4681;
  assign n7435 = \[4427]  & Ng4646;
  assign n7436 = ~n7434 & ~n7435;
  assign n7437 = ~Ng4826 & Ng4688;
  assign n7438 = Ng4674 & ~Ng4821;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~n7423 & n7439;
  assign n7441 = n7436 & n7440;
  assign n7442 = Pg35 & ~n7441;
  assign n6681 = ~n7433 & n7442;
  assign n7444 = ~Pg35 & \[4437] ;
  assign n2218_1 = n6681 | n7444;
  assign n7446 = ~Pg35 & Ng4093;
  assign n7447 = ~Ng4098 & ~n6477;
  assign n7448 = n6479 & ~n7447;
  assign n7449 = ~n6197_1 & ~n7448;
  assign n2223_1 = n7446 | ~n7449;
  assign n7451 = \[4437]  & n5406;
  assign n7452 = Ng4495 & ~n5406;
  assign n7453 = ~n5408 & ~n7452;
  assign n2228_1 = n7451 | ~n7453;
  assign n7455 = ~Pg35 & ~Ng518;
  assign n7456 = ~Ng528 & ~n5353;
  assign n7457 = ~n5356 & ~n7456;
  assign n7458 = Pg35 & ~n7457;
  assign n7459 = ~n5349 & ~n7458;
  assign n2233_1 = ~n7455 & n7459;
  assign n7461 = Ng3139 & n5955;
  assign n7462 = Ng3133 & ~n5955;
  assign n2243_1 = n7461 | n7462;
  assign n7464 = ~Ng232 & n5407;
  assign n7465 = ~Pg73 & Pg72;
  assign n7466 = ~Ng239 & n7465;
  assign n7467 = ~n7464 & ~n7466;
  assign n7468 = ~Ng225 & n6134;
  assign n7469 = ~Ng246 & n5182;
  assign n7470 = ~n7468 & ~n7469;
  assign n7471 = n7467 & n7470;
  assign n7472 = Pg35 & n7471;
  assign n7473 = ~Pg35 & Ng479;
  assign n2248_1 = n7472 | n7473;
  assign n7475 = ~Pg35 & Ng4332;
  assign n7476 = Pg35 & n5568;
  assign n7477 = ~Ng4584 & ~n5565;
  assign n7478 = ~n5566 & ~n7477;
  assign n7479 = n7476 & n7478;
  assign n2253_1 = n7475 | n7479;
  assign n7481 = ~Pg35 & Ng298;
  assign n7482 = Ng142 & n5713;
  assign n7483 = ~n6927 & ~n7482;
  assign n7484 = ~n6928 & ~n7483;
  assign n2258_1 = n7481 | n7484;
  assign n7486 = Ng5831 & n6560;
  assign n7487 = Pg35 & ~Ng5821;
  assign n7488 = Ng5827 & ~n7487;
  assign n7489 = ~Ng5827 & n7487;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = ~n6560 & ~n7490;
  assign n2266_1 = n7486 | n7491;
  assign n7493 = Pg14125 & n7390;
  assign n7494 = ~Pg35 & Ng262;
  assign n7495 = Ng239 & n7393;
  assign n7496 = ~n7494 & ~n7495;
  assign n2271_1 = n7493 | ~n7496;
  assign n7498 = ~Pg35 & Ng1221;
  assign n7499 = Ng1205 & Ng1087;
  assign n7500 = Ng1221 & n7499;
  assign n7501 = Ng1216 & n7500;
  assign n7502 = Ng1211 & n7500;
  assign n7503 = Pg35 & ~n7502;
  assign n7504 = ~Ng1216 & ~n7500;
  assign n7505 = n7503 & ~n7504;
  assign n7506 = ~n7501 & n7505;
  assign n2276_1 = n7498 | n7506;
  assign n7508 = Pg35 & ~Ng2848;
  assign n7509 = n5798 & n7508;
  assign n7510 = ~Pg35 & ~\[4433] ;
  assign n2281_1 = ~n7509 & ~n7510;
  assign n7512 = Pg9553 & ~Ng5112;
  assign n7513 = ~Ng5022 & ~n7512;
  assign n7514 = Pg35 & ~Pg9497;
  assign n7515 = ~n7513 & n7514;
  assign n7516 = ~Pg35 & Ng5112;
  assign n2286 = n7515 | n7516;
  assign n7518 = ~Pg35 & Ng1024;
  assign n7519 = ~Ng1030 & ~n5623;
  assign n7520 = ~n5994 & ~n7519;
  assign n2294_1 = n7518 | n7520;
  assign n7522 = ~Ng3179 & ~Ng3171;
  assign n7523 = n5015 & n7522;
  assign n7524 = Pg35 & ~n7523;
  assign n7525 = ~Pg35 & ~Ng3215;
  assign n7526 = ~n5018 & ~n7525;
  assign n7527 = ~n7524 & ~n7526;
  assign n7528 = ~Ng3231 & n7524;
  assign n2302_1 = ~n7527 & ~n7528;
  assign n7530 = Pg35 & Ng6727;
  assign n7531 = ~Pg35 & Ng6444;
  assign n2307 = n7530 | n7531;
  assign n7533 = ~Pg35 & Ng2227;
  assign n7534 = ~Ng2241 & n6498_1;
  assign n7535 = Ng1589 & ~n6496;
  assign n7536 = ~n6503_1 & ~n7535;
  assign n7537 = ~Ng2153 & ~Ng2227;
  assign n7538 = Ng2241 & ~n7537;
  assign n7539 = n7536 & n7538;
  assign n7540 = ~n7536 & ~n7538;
  assign n7541 = ~n7539 & ~n7540;
  assign n7542 = ~n6498_1 & n7541;
  assign n7543 = Pg35 & ~n7542;
  assign n7544 = ~n7534 & n7543;
  assign n2319_1 = n7533 | n7544;
  assign n7546 = ~Pg35 & Ng1548;
  assign n7547 = Ng1430 & Ng1548;
  assign n7548 = Ng1564 & n7547;
  assign n7549 = Pg35 & Ng1564;
  assign n7550 = ~n7547 & ~n7549;
  assign n7551 = ~n7548 & ~n7550;
  assign n2324 = n7546 | n7551;
  assign n7553 = Pg35 & Ng6035;
  assign n7554 = ~Pg35 & Ng5752;
  assign n2329_1 = n7553 | n7554;
  assign n7556 = Ng6549 & Ng6555;
  assign n7557 = Ng6573 & ~Ng6565;
  assign n7558 = n7556 & n7557;
  assign n7559 = Pg35 & ~n7558;
  assign n7560 = Ng6649 & n7559;
  assign n7561 = ~Pg35 & Ng6633;
  assign n7562 = ~n5083 & ~n7561;
  assign n7563 = ~n7559 & ~n7562;
  assign n2337 = n7560 | n7563;
  assign n7565 = Ng225 & n7393;
  assign n7566 = Pg14189 & n7390;
  assign n7567 = ~Pg35 & Ng872;
  assign n7568 = ~n7566 & ~n7567;
  assign n2350 = n7565 | ~n7568;
  assign n7570 = ~Pg35 & Ng4483;
  assign n2355_1 = n5953 | n7570;
  assign n7572 = n5406 & ~n7465;
  assign n7573 = Ng4501 & ~n5406;
  assign n7574 = ~n7451 & ~n7573;
  assign n2360 = n7572 | ~n7574;
  assign n7576 = n4716 & n5203;
  assign n7577 = ~Ng5873 & ~n7576;
  assign n7578 = Pg35 & ~n7577;
  assign n7579 = Ng5869 & ~n7578;
  assign n7580 = Pg35 & ~n7576;
  assign n7581 = ~Ng5869 & n7580;
  assign n7582 = Ng5873 & n7581;
  assign n2365 = n7579 | n7582;
  assign n7584 = ~n4902 & ~n4909;
  assign n7585 = Pg35 & ~Ng5037;
  assign n7586 = ~n7584 & n7585;
  assign n7587 = ~Ng5057 & Ng5046;
  assign n7588 = n4917 & n7587;
  assign n7589 = Ng5062 & n7588;
  assign n7590 = Pg35 & ~n7589;
  assign n7591 = ~n4920_1 & n7590;
  assign n7592 = Ng5037 & n7584;
  assign n7593 = n7591 & n7592;
  assign n7594 = ~Pg35 & Ng5033;
  assign n7595 = ~n7593 & ~n7594;
  assign n2370_1 = n7586 | ~n7595;
  assign n7597 = Ng2319 & n7142;
  assign n7598 = Ng2342 & ~Ng2319;
  assign n7599 = Pg35 & ~n7598;
  assign n7600 = n7141 & n7599;
  assign n7601 = ~Ng2351 & n7600;
  assign n7602 = ~n7597 & ~n7601;
  assign n7603 = ~Pg35 & Ng2327;
  assign n7604 = ~n7146 & ~n7603;
  assign n2375 = ~n7602 | ~n7604;
  assign n7606 = Ng5495 & n7205;
  assign n7607 = Ng5489 & ~n7205;
  assign n2380_1 = n7606 | n7607;
  assign n7609 = Ng4164 & Ng4253;
  assign n7610 = Ng4145 & ~Ng4253;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = Pg35 & n7611;
  assign n7613 = ~Pg35 & Ng4180;
  assign n2385_1 = n7612 | n7613;
  assign n7615 = ~Ng5164 & ~Ng5170;
  assign n7616 = ~Ng5176 & n7615;
  assign n7617 = n5041 & n7616;
  assign n7618 = Pg35 & ~n7617;
  assign n7619 = ~Pg35 & ~Ng5212;
  assign n7620 = ~n5018 & ~n7619;
  assign n7621 = ~n7618 & ~n7620;
  assign n7622 = ~Ng5208 & n7618;
  assign n2389 = ~n7621 & ~n7622;
  assign n7624 = Ng5511 & ~Ng5517;
  assign n7625 = n6172 & n7624;
  assign n7626 = Pg35 & ~n7625;
  assign n7627 = Ng5579 & n7626;
  assign n7628 = ~Pg35 & Ng5555;
  assign n7629 = ~n5083 & ~n7628;
  assign n7630 = ~n7626 & ~n7629;
  assign n2394_1 = n7627 | n7630;
  assign n7632 = ~Pg35 & Ng5863;
  assign n7633 = n7328 & n7581;
  assign n2399_1 = n7632 | n7633;
  assign n7635 = ~Pg35 & Ng1585;
  assign n2404_1 = n5591 | n7635;
  assign n7637 = Pg9617 & ~Ng5802;
  assign n7638 = ~Ng5752 & ~n7637;
  assign n7639 = Pg35 & ~Pg9680;
  assign n7640 = ~n7638 & n7639;
  assign n7641 = ~Pg35 & Ng5802;
  assign n2409_1 = n7640 | n7641;
  assign n7643 = n5497 & n7336;
  assign n7644 = Pg35 & ~n7643;
  assign n7645 = Ng6279 & n7644;
  assign n7646 = ~Pg35 & Ng6263;
  assign n7647 = ~n5083 & ~n7646;
  assign n7648 = ~n7644 & ~n7647;
  assign n2414_1 = n7645 | n7648;
  assign n7650 = ~Ng5863 & Ng5857;
  assign n7651 = n6427 & n7650;
  assign n7652 = n5083 & n7651;
  assign n7653 = ~Pg35 & Ng5889;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = Pg35 & Ng5917;
  assign n7656 = ~n7651 & n7655;
  assign n2419_1 = ~n7654 | n7656;
  assign n7658 = ~Pg35 & ~Ng2965;
  assign n7659 = Ng962 & n6452;
  assign n7660 = ~Ng2975 & n7659;
  assign n2424_1 = ~n7658 & ~n7660;
  assign n7662 = ~Ng6167 & n7023;
  assign n7663 = ~Pg35 & Ng6163;
  assign n7664 = ~n5388 & ~n7663;
  assign n7665 = ~n7023 & n7664;
  assign n2429 = ~n7662 & ~n7665;
  assign n7667 = ~Pg35 & Ng2606;
  assign n7668 = Pg35 & n5533;
  assign n7669 = Ng2599 & n7668;
  assign n7670 = Ng2555 & ~n5533;
  assign n7671 = n4567 & n5089;
  assign n7672 = Pg35 & ~n7671;
  assign n7673 = n7670 & n7672;
  assign n7674 = ~n7669 & ~n7673;
  assign n2437_1 = n7667 | ~n7674;
  assign n7676 = ~Pg35 & Ng1454;
  assign n7677 = ~Ng1495 & Ng1442;
  assign n7678 = Ng1454 & n6436;
  assign n7679 = n7677 & n7678;
  assign n7680 = ~Ng1448 & n7679;
  assign n7681 = ~n7676 & ~n7680;
  assign n7682 = Pg35 & Ng1448;
  assign n7683 = ~n7679 & n7682;
  assign n2442 = ~n7681 | n7683;
  assign n7685 = ~Pg35 & Ng2351;
  assign n7686 = Ng2319 & n7141;
  assign n7687 = Ng2351 & n7686;
  assign n7688 = Ng2299 & n7687;
  assign n7689 = ~n7685 & ~n7688;
  assign n7690 = Pg35 & n7141;
  assign n7691 = Ng2319 & Ng2311;
  assign n7692 = ~Ng2342 & n7691;
  assign n7693 = Ng2315 & n4667;
  assign n7694 = Ng2295 & n7598;
  assign n7695 = ~n7693 & ~n7694;
  assign n7696 = ~Ng2342 & Ng2351;
  assign n7697 = Ng2303 & n7696;
  assign n7698 = ~Ng2319 & Ng2307;
  assign n7699 = ~Ng2351 & n7698;
  assign n7700 = ~n7697 & ~n7699;
  assign n7701 = n7695 & n7700;
  assign n7702 = ~n7692 & n7701;
  assign n7703 = n7690 & ~n7702;
  assign n7704 = Ng2370 & n7142;
  assign n7705 = ~n7703 & ~n7704;
  assign n2450_1 = ~n7689 | ~n7705;
  assign n2455 = ~Ng5164 & n5599;
  assign n7708 = ~Pg35 & Ng150;
  assign n7709 = Ng153 & n7270;
  assign n7710 = ~n7267 & ~n7709;
  assign n7711 = ~n7268 & ~n7710;
  assign n2464_1 = n7708 | n7711;
  assign n7713 = n4712 & n5203;
  assign n7714 = Pg35 & ~n7713;
  assign n7715 = ~Ng6561 & n7714;
  assign n2469_1 = ~Ng6549 & n7715;
  assign n7717 = ~Pg35 & Ng4076;
  assign n7718 = Pg35 & Ng2841;
  assign n7719 = ~Ng4087 & ~n6203;
  assign n7720 = ~n6476 & ~n7719;
  assign n7721 = n7718 & n7720;
  assign n2474_1 = n7717 | n7721;
  assign n7723 = ~Ng4801 & n5554;
  assign n7724 = ~n5549 & n5552;
  assign n7725 = Ng4801 & n7724;
  assign n7726 = ~Pg35 & Ng4793;
  assign n7727 = ~n7725 & ~n7726;
  assign n2479_1 = n7723 | ~n7727;
  assign n7729 = ~Pg35 & ~Ng2980;
  assign n7730 = ~Pg54 & ~Pg53;
  assign n7731 = ~Pg56 & n7730;
  assign n7732 = n3297 & n7731;
  assign n7733 = Pg35 & ~Ng2984;
  assign n7734 = ~n7732 & n7733;
  assign n2484_1 = ~n7729 & ~n7734;
  assign n7736 = Ng3863 & Ng3857;
  assign n7737 = n4733 & n7736;
  assign n7738 = Pg35 & ~n7737;
  assign n7739 = ~Pg35 & ~Ng3945;
  assign n7740 = ~n5018 & ~n7739;
  assign n7741 = ~n7738 & ~n7740;
  assign n7742 = ~Ng3961 & n7738;
  assign n2489_1 = ~n7741 & ~n7742;
  assign n7744 = ~Pg35 & Ng1178;
  assign n7745 = Ng1171 & Ng1183;
  assign n7746 = n6075 & n7745;
  assign n7747 = Pg35 & Ng962;
  assign n7748 = Pg35 & Ng1183;
  assign n7749 = n6579 & n7748;
  assign n7750 = ~n7747 & ~n7749;
  assign n7751 = ~n7746 & ~n7750;
  assign n2494 = n7744 | n7751;
  assign n7753 = ~Ng6573 & ~Ng6565;
  assign n7754 = n7103 & n7753;
  assign n7755 = n5083 & n7754;
  assign n7756 = ~Pg35 & Ng6609;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = Pg35 & Ng6625;
  assign n7759 = ~n7754 & n7758;
  assign n2507_1 = ~n7757 | n7759;
  assign n7761 = ~Pg35 & Ng1002;
  assign n7762 = ~Ng1018 & ~n5618;
  assign n7763 = Pg35 & ~n5620;
  assign n7764 = ~n7762 & n7763;
  assign n2517_1 = n7761 | n7764;
  assign n7766 = Ng1554 & n7548;
  assign n7767 = ~n5511 & n7766;
  assign n7768 = Pg35 & ~Pg17320;
  assign n7769 = ~Pg17404 & ~Pg17423;
  assign n7770 = n7768 & n7769;
  assign n2522_1 = ~n7767 & n7770;
  assign n7772 = ~Pg35 & Ng4040;
  assign n7773 = ~Ng4049 & n4998;
  assign n2526_1 = n7772 | n7773;
  assign n7775 = Pg13272 & Ng1514;
  assign n7776 = Ng1526 & n7775;
  assign n7777 = ~Ng1472 & n6271_1;
  assign n7778 = Ng1472 & ~n6271_1;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = n7776 & n7779;
  assign n7781 = n6276_1 & n7776;
  assign n7782 = ~Ng1467 & ~n7781;
  assign n7783 = Pg35 & ~n7782;
  assign n7784 = ~n7780 & n7783;
  assign n7785 = ~Pg35 & Ng1448;
  assign n2531 = n7784 | n7785;
  assign n7787 = Pg35 & ~n4649_1;
  assign n7788 = ~n6149 & ~n7787;
  assign n7789 = Ng2461 & ~n7788;
  assign n7790 = Ng2465 & ~Ng2421;
  assign n7791 = Pg35 & ~n7790;
  assign n7792 = ~Pg35 & Ng2441;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = n7788 & ~n7793;
  assign n2536_1 = n7789 | n7794;
  assign n7796 = ~Pg35 & ~Ng2748;
  assign n7797 = Ng2724 & n5327;
  assign n7798 = Ng2729 & n7797;
  assign n7799 = n4930 & n7798;
  assign n7800 = Ng2735 & n7798;
  assign n7801 = Ng2741 & n7800;
  assign n7802 = ~Ng2756 & ~n7801;
  assign n7803 = ~n4656 & ~n7802;
  assign n7804 = ~n7799 & n7803;
  assign n7805 = n7718 & ~n7804;
  assign n2541_1 = ~n7796 & ~n7805;
  assign n7807 = Ng6049 & ~n6856;
  assign n7808 = Pg35 & Ng5990;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = n4540 & n5933;
  assign n7811 = ~n4551 & ~n7810;
  assign n7812 = n6791 & ~n7811;
  assign n2546_1 = ~n7809 & ~n7812;
  assign n7814 = ~Pg35 & Ng1252;
  assign n7815 = Ng1249 & Pg12923;
  assign n7816 = Ng1266 & n7815;
  assign n7817 = Ng1280 & n7816;
  assign n7818 = Ng1252 & n7817;
  assign n7819 = Ng1256 & n7818;
  assign n7820 = Ng1256 & n5591;
  assign n7821 = ~n7818 & ~n7820;
  assign n7822 = ~n7819 & ~n7821;
  assign n2551_1 = n7814 | n7822;
  assign n7824 = Ng5029 & ~n4920_1;
  assign n7825 = ~Ng5062 & ~n7824;
  assign n7826 = ~n4900 & ~n7825;
  assign n7827 = Pg35 & ~n7826;
  assign n7828 = Ng5016 & ~n7827;
  assign n7829 = ~Ng5016 & n7591;
  assign n7830 = ~Ng5022 & Ng5029;
  assign n7831 = n7829 & n7830;
  assign n7832 = Pg35 & n4908;
  assign n7833 = ~n7831 & ~n7832;
  assign n2556 = n7828 | ~n7833;
  assign n7835 = n4684 & n5481;
  assign n7836 = Ng4836 & ~n7835;
  assign n7837 = Ng6727 & n4538;
  assign n7838 = Pg17722 & n7837;
  assign n7839 = n7836 & n7838;
  assign n7840 = Pg35 & ~n7839;
  assign n7841 = Ng6519 & n7840;
  assign n7842 = Ng6513 & ~n7840;
  assign n2561_1 = n7841 | n7842;
  assign n7844 = ~Pg35 & Ng1802;
  assign n7845 = ~Ng1816 & n5063;
  assign n7846 = ~Ng1246 & ~n5061_1;
  assign n7847 = ~n5068 & ~n7846;
  assign n7848 = ~Ng1802 & ~Ng1728;
  assign n7849 = Ng1816 & ~n7848;
  assign n7850 = n7847 & n7849;
  assign n7851 = ~n7847 & ~n7849;
  assign n7852 = ~n7850 & ~n7851;
  assign n7853 = ~n5063 & n7852;
  assign n7854 = Pg35 & ~n7853;
  assign n7855 = ~n7845 & n7854;
  assign n2566 = n7844 | n7855;
  assign n7857 = ~Pg35 & ~Ng4459;
  assign n7858 = Pg35 & ~Ng4473;
  assign n2571_1 = ~n7857 & ~n7858;
  assign n7860 = ~Pg35 & Ng4572;
  assign n2576_1 = n1655_1 | n7860;
  assign n7862 = ~Ng4507 & ~n4561;
  assign n7863 = n5182 & ~n7862;
  assign n7864 = Ng26960 & ~n7863;
  assign n7865 = ~Ng4477 & n7864;
  assign n7866 = Ng10384 & Ng4462;
  assign n7867 = ~n7865 & n7866;
  assign n2581 = Pg35 & ~n7867;
  assign n7869 = Ng3831 & n7017;
  assign n7870 = Pg35 & ~Ng3821;
  assign n7871 = Ng3827 & ~n7870;
  assign n7872 = ~Ng3827 & n7870;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = ~n7017 & ~n7873;
  assign n2586_1 = n7869 | n7874;
  assign n7876 = Ng2509 & n7009;
  assign n7877 = Ng2514 & ~n7009;
  assign n2591_1 = n7876 | n7877;
  assign n7879 = n4689 & n5481;
  assign n7880 = Ng4864 & ~n7879;
  assign n7881 = n4531 & n7880;
  assign n7882 = n7083 & n7881;
  assign n7883 = Ng3288 & ~n7880;
  assign n7884 = ~n4532 & n7880;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n7882 & ~n7885;
  assign n7887 = Pg35 & ~n7886;
  assign n7888 = Pg35 & Ng3288;
  assign n7889 = ~Ng3352 & ~n7888;
  assign n2596 = ~n7887 & ~n7889;
  assign n7891 = Pg35 & ~Ng2393;
  assign n7892 = Ng2399 & ~n7891;
  assign n7893 = ~Ng2399 & n7891;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n4981 & n7894;
  assign n7896 = ~Ng2403 & n4981;
  assign n2601_1 = ~n7895 & ~n7896;
  assign n7898 = Pg35 & Ng2145;
  assign n7899 = ~Pg35 & Ng2138;
  assign n2606_1 = n7898 | n7899;
  assign n7901 = Ng1657 & n6249;
  assign n7902 = Ng1624 & n7901;
  assign n7903 = Pg35 & ~n7902;
  assign n7904 = ~Ng1700 & n7903;
  assign n7905 = Pg35 & ~Ng1700;
  assign n7906 = ~Pg35 & Ng1696;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = ~n7903 & n7907;
  assign n2611_1 = ~n7904 & ~n7908;
  assign n7910 = Pg35 & ~n5351;
  assign n7911 = Ng513 & n7910;
  assign n7912 = ~n5349 & ~n7910;
  assign n7913 = Ng504 & n7912;
  assign n2616_1 = n7911 | n7913;
  assign n7915 = ~Pg35 & Ng5357;
  assign n7916 = n4537 & n5933;
  assign n7917 = ~Pg31860 & ~n7916;
  assign n7918 = Pg33959 & ~n7917;
  assign n7919 = Pg35 & Ng5297;
  assign n7920 = Pg33959 & n6011;
  assign n7921 = ~n7919 & ~n7920;
  assign n7922 = ~n7918 & ~n7921;
  assign n2625_1 = n7915 | n7922;
  assign n7924 = Pg35 & Ng2763;
  assign n7925 = Pg35 & ~n7799;
  assign n7926 = Ng2759 & ~n7925;
  assign n7927 = n7924 & ~n7926;
  assign n7928 = ~n7924 & n7926;
  assign n7929 = ~n7927 & ~n7928;
  assign n2630_1 = n6197_1 | ~n7929;
  assign n7931 = ~Ng4793 & ~n4619;
  assign n7932 = n7724 & ~n7931;
  assign n2635_1 = n6598 | n7932;
  assign n7934 = ~Pg35 & ~Ng947;
  assign n7935 = ~Ng952 & n7747;
  assign n2640_1 = ~n7934 & ~n7935;
  assign n7937 = ~Pg35 & Ng1259;
  assign n7938 = Ng1259 & n7819;
  assign n7939 = Ng1263 & n7938;
  assign n7940 = Ng1263 & n5591;
  assign n7941 = ~n7938 & ~n7940;
  assign n7942 = ~n7939 & ~n7941;
  assign n2645_1 = n7937 | n7942;
  assign n7944 = ~Pg35 & Ng1936;
  assign n7945 = ~Ng1950 & n4950;
  assign n7946 = Ng1246 & ~n4948;
  assign n7947 = ~n4958 & ~n7946;
  assign n7948 = ~Ng1862 & ~Ng1936;
  assign n7949 = Ng1950 & ~n7948;
  assign n7950 = n7947 & n7949;
  assign n7951 = ~n7947 & ~n7949;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~n4950 & n7952;
  assign n7954 = Pg35 & ~n7953;
  assign n7955 = ~n7945 & n7954;
  assign n2650_1 = n7944 | n7955;
  assign n7957 = Ng5138 & n6143_1;
  assign n7958 = Pg35 & ~Ng5128;
  assign n7959 = n6142 & n7958;
  assign n7960 = ~Ng5134 & n7959;
  assign n7961 = ~n7957 & ~n7960;
  assign n7962 = Ng5134 & ~n7958;
  assign n7963 = ~n6143_1 & n7962;
  assign n2655_1 = ~n7961 | n7963;
  assign n7965 = Ng2287 & ~n4978;
  assign n7966 = Ng2361 & n7965;
  assign n7967 = Pg35 & ~n7966;
  assign n7968 = Ng2307 & n7967;
  assign n7969 = ~Pg35 & Ng2311;
  assign n7970 = ~n4986 & ~n7969;
  assign n7971 = ~n7967 & ~n7970;
  assign n2660_1 = n7968 | n7971;
  assign n7973 = Pg35 & Ng4040;
  assign n7974 = ~Pg35 & Ng3752;
  assign n2669_1 = n7973 | n7974;
  assign n7976 = ~Pg35 & Ng4659;
  assign n7977 = ~n4619 & ~n5548;
  assign n7978 = Pg35 & n7977;
  assign n7979 = Ng4664 & n4618_1;
  assign n7980 = ~Ng4664 & ~n4618_1;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = n7978 & n7981;
  assign n2673_1 = n7976 | n7982;
  assign n7984 = n4644 & n5258;
  assign n7985 = n4928 & n7984;
  assign n7986 = Ng2223 & ~n7985;
  assign n7987 = Pg35 & n7986;
  assign n7988 = Ng110 & n5268;
  assign n7989 = ~Ng110 & ~n5268;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = n5842 & n7990;
  assign n7992 = n7984 & n7991;
  assign n7993 = ~Pg35 & Ng2208;
  assign n7994 = ~n7992 & ~n7993;
  assign n2678_1 = n7987 | ~n7994;
  assign n7996 = ~Pg35 & Ng5813;
  assign n7997 = n6559 & n6854;
  assign n7998 = Pg35 & Ng5808;
  assign n7999 = n6556_1 & ~n6558;
  assign n8000 = ~n6854 & n7999;
  assign n8001 = n7998 & ~n8000;
  assign n8002 = ~n7997 & n8001;
  assign n8003 = ~Ng5808 & n6855;
  assign n8004 = ~n8002 & ~n8003;
  assign n2683_1 = n7996 | ~n8004;
  assign n8006 = ~Pg35 & ~Ng6629;
  assign n8007 = n7380 & n7556;
  assign n8008 = n5018 & n8007;
  assign n8009 = Pg35 & ~Ng6645;
  assign n8010 = ~n8007 & n8009;
  assign n8011 = ~n8008 & ~n8010;
  assign n2688_1 = ~n8006 & n8011;
  assign n8013 = Ng1996 & ~n5660;
  assign n8014 = Ng2070 & n8013;
  assign n8015 = Pg35 & ~n8014;
  assign n8016 = Ng2016 & n8015;
  assign n8017 = ~Pg35 & Ng2020;
  assign n8018 = ~n6912 & ~n8017;
  assign n8019 = ~n8015 & ~n8018;
  assign n2693_1 = n8016 | n8019;
  assign n8021 = n4704 & n5105;
  assign n8022 = ~Ng3873 & ~n8021;
  assign n8023 = Pg35 & ~n8022;
  assign n8024 = Ng3869 & ~n8023;
  assign n8025 = Pg35 & ~n8021;
  assign n8026 = ~Ng3869 & n8025;
  assign n8027 = Ng3873 & n8026;
  assign n2698_1 = n8024 | n8027;
  assign n8029 = n4587 & ~n4978;
  assign n8030 = Pg35 & ~n8029;
  assign n8031 = ~Ng2315 & n8030;
  assign n8032 = ~Pg35 & Ng2303;
  assign n8033 = ~n4986 & ~n8030;
  assign n8034 = ~n8032 & n8033;
  assign n2706_1 = ~n8031 & ~n8034;
  assign n8036 = Pg35 & ~n4657;
  assign n8037 = Ng2811 & n8036;
  assign n8038 = Pg35 & ~n4930;
  assign n8039 = ~n4656 & n8038;
  assign n8040 = ~Ng2327 & n8039;
  assign n8041 = ~Pg35 & Ng2799;
  assign n8042 = ~n8040 & ~n8041;
  assign n2711_1 = n8037 | ~n8042;
  assign n8044 = n6754 & n7328;
  assign n8045 = n5018 & n8044;
  assign n8046 = ~Pg35 & ~Ng5941;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = Pg35 & ~n8044;
  assign n8049 = ~Ng5957 & n8048;
  assign n2716_1 = n8047 & ~n8049;
  assign n8051 = ~Pg35 & Ng1996;
  assign n8052 = ~Ng112 & ~n4596;
  assign n8053 = Ng112 & n4596;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = n4595 & n5656;
  assign n8056 = n8054 & n8055;
  assign n8057 = n5842 & n8056;
  assign n8058 = ~n8051 & ~n8057;
  assign n8059 = n4928 & n8055;
  assign n8060 = Ng2047 & ~n8059;
  assign n8061 = Pg35 & n8060;
  assign n2721_1 = ~n8058 | n8061;
  assign n8063 = ~Pg35 & Ng3863;
  assign n8064 = n7736 & n8026;
  assign n2726_1 = n8063 | n8064;
  assign n8066 = n5317 & n7624;
  assign n8067 = Pg35 & ~n8066;
  assign n8068 = Ng5575 & n8067;
  assign n8069 = ~Pg35 & Ng5547;
  assign n8070 = ~n5083 & ~n8069;
  assign n8071 = ~n8067 & ~n8070;
  assign n2734_1 = n8068 | n8071;
  assign n8073 = Pg8344 & ~Ng3802;
  assign n8074 = ~Ng3752 & ~n8073;
  assign n8075 = Pg35 & ~Pg8398;
  assign n8076 = ~n8074 & n8075;
  assign n8077 = ~Pg35 & Ng3802;
  assign n2744_1 = n8076 | n8077;
  assign n8079 = ~Ng3863 & Ng3857;
  assign n8080 = n6919 & n8079;
  assign n8081 = n5083 & n8080;
  assign n8082 = ~Pg35 & Ng3889;
  assign n8083 = ~n8081 & ~n8082;
  assign n8084 = Pg35 & Ng3917;
  assign n8085 = ~n8080 & n8084;
  assign n2749 = ~n8083 | n8085;
  assign n8087 = Pg35 & Ng4411;
  assign n8088 = Ng4401 & ~n6864;
  assign n8089 = ~n6861 & n8088;
  assign n2761_1 = n8087 | n8089;
  assign n8091 = n4723 & n6386;
  assign n8092 = Pg35 & ~n8091;
  assign n8093 = ~Pg35 & ~Ng6255;
  assign n8094 = ~n5018 & ~n8093;
  assign n8095 = ~n8092 & ~n8094;
  assign n8096 = ~Ng6275 & n8092;
  assign n2766_1 = ~n8095 & ~n8096;
  assign n8098 = Ng6311 & n7023;
  assign n8099 = ~Pg35 & Ng6307;
  assign n8100 = ~n5083 & ~n8099;
  assign n8101 = ~n7023 & ~n8100;
  assign n2771_1 = n8098 | n8101;
  assign n8103 = ~Ng1041 & Ng1008;
  assign n8104 = n7062 & ~n8103;
  assign n8105 = Pg35 & n8104;
  assign n8106 = ~Pg35 & ~Ng1036;
  assign n8107 = ~Ng1041 & n7063;
  assign n8108 = ~n8106 & ~n8107;
  assign n2779_1 = ~n8105 & n8108;
  assign n8110 = ~Pg35 & ~Ng2575;
  assign n8111 = ~Ng2619 & n5329;
  assign n8112 = Ng2610 & n8111;
  assign n8113 = Ng2599 & ~Ng2555;
  assign n8114 = n8112 & ~n8113;
  assign n8115 = Ng2595 & ~n8112;
  assign n8116 = Pg35 & ~n8115;
  assign n8117 = ~n8114 & n8116;
  assign n2784_1 = ~n8110 & ~n8117;
  assign n8119 = ~Ng2537 & ~n7009;
  assign n8120 = Pg35 & ~Ng2527;
  assign n8121 = Ng2533 & n8120;
  assign n8122 = ~Ng2533 & ~n8120;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = n7009 & ~n8123;
  assign n2789_1 = ~n8119 & ~n8124;
  assign n8126 = Pg35 & \[4426] ;
  assign n8127 = ~Pg35 & Ng550;
  assign n2794_1 = n8126 | n8127;
  assign n8129 = Pg35 & Ng4443;
  assign n8130 = Pg35 & ~n7403;
  assign n8131 = Ng4434 & ~n6864;
  assign n8132 = ~n8130 & n8131;
  assign n2799_1 = n8129 | n8132;
  assign n8134 = ~Pg35 & Ng4561;
  assign n2804_1 = n5989 | n8134;
  assign n8136 = Ng4826 & n5937;
  assign n8137 = ~Pg35 & Ng6311;
  assign n8138 = ~n8136 & ~n8137;
  assign n2809_1 = n6353 | ~n8138;
  assign n8140 = n6227_1 & n6385;
  assign n8141 = n5083 & n8140;
  assign n8142 = ~Pg35 & Ng6243;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = Pg35 & Ng6239;
  assign n8145 = ~n8140 & n8144;
  assign n2814_1 = ~n8143 | n8145;
  assign n8147 = Ng232 & n7393;
  assign n8148 = ~Pg35 & Ng255;
  assign n8149 = Pg14217 & n7390;
  assign n8150 = ~n8148 & ~n8149;
  assign n2819 = n8147 | ~n8150;
  assign n8152 = n4708_1 & n6412;
  assign n8153 = n5083 & n8152;
  assign n8154 = ~Pg35 & Ng5252;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = Pg35 & Ng5268;
  assign n8157 = ~n8152 & n8156;
  assign n2824_1 = ~n8155 | n8157;
  assign n2829_1 = Pg35 & Ng6545;
  assign n8160 = Pg35 & ~n7687;
  assign n8161 = Pg35 & ~Ng2407;
  assign n8162 = Ng2413 & n8161;
  assign n8163 = ~Ng2413 & ~n8161;
  assign n8164 = ~n8162 & ~n8163;
  assign n8165 = ~n8160 & ~n8164;
  assign n8166 = ~Ng2417 & n8160;
  assign n2834_1 = ~n8165 & ~n8166;
  assign n8168 = n6996 & n7183;
  assign n8169 = ~Pg35 & Ng1779;
  assign n8170 = Ng1772 & n5087;
  assign n8171 = ~n8169 & ~n8170;
  assign n2839_1 = n8168 | ~n8171;
  assign n8173 = ~Pg35 & Ng5046;
  assign n8174 = Pg35 & n4912;
  assign n8175 = ~n4905_1 & ~n8174;
  assign n8176 = ~Ng5052 & ~n8175;
  assign n8177 = n4906 & n7591;
  assign n8178 = ~n4912 & n8177;
  assign n8179 = ~n8176 & ~n8178;
  assign n2844_1 = n8173 | ~n8179;
  assign n8181 = Pg35 & Ng5689;
  assign n8182 = ~Pg35 & Ng5406;
  assign n2849_1 = n8181 | n8182;
  assign n8184 = ~Pg35 & Ng1878;
  assign n8185 = n4580 & ~n4950;
  assign n8186 = Pg35 & ~n8185;
  assign n8187 = ~n4960 & ~n8186;
  assign n8188 = ~n8184 & n8187;
  assign n8189 = ~Ng1890 & n8186;
  assign n2853_1 = ~n8188 & ~n8189;
  assign n8191 = Pg35 & n7671;
  assign n8192 = Ng2599 & ~n7668;
  assign n8193 = ~n8191 & n8192;
  assign n8194 = Ng2629 & n7668;
  assign n2858_1 = n8193 | n8194;
  assign n8196 = ~Pg35 & Ng568;
  assign n8197 = Ng572 & n5737;
  assign n8198 = ~n5748 & ~n8197;
  assign n8199 = ~n5749 & ~n8198;
  assign n2863_1 = n8196 | n8199;
  assign n2868_1 = Pg35 & Ng2130;
  assign n8202 = ~Ng4108 & ~n6478_1;
  assign n8203 = ~n6480 & ~n8202;
  assign n8204 = ~Pg35 & Ng4098;
  assign n8205 = ~n6197_1 & ~n8204;
  assign n2873_1 = n8203 | ~n8205;
  assign n8207 = ~Pg35 & Ng424;
  assign n8208 = Ng475 & n5151;
  assign n8209 = Ng246 & n6741;
  assign n8210 = ~n8208 & ~n8209;
  assign n2882_1 = n8207 | ~n8210;
  assign n3848 = Pg64 & Pg35;
  assign n8213 = ~Pg35 & Ng753;
  assign n2896 = n3848 | n8213;
  assign n8215 = ~Pg35 & Ng4054;
  assign n8216 = ~n4535 & ~n7084;
  assign n8217 = n6689 & ~n8216;
  assign n8218 = Ng4054 & ~Ng3990;
  assign n8219 = n6689 & n8218;
  assign n8220 = Pg35 & Ng3990;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = ~n8217 & ~n8221;
  assign n2900_1 = n8215 | n8222;
  assign n8224 = ~Pg35 & Ng5873;
  assign n8225 = n1065_1 & ~n5782_1;
  assign n8226 = ~n5783 & ~n8225;
  assign n8227 = ~n7576 & ~n8226;
  assign n2905_1 = n8224 | n8227;
  assign n8229 = Ng1992 & n5300;
  assign n8230 = Pg35 & ~Ng1982;
  assign n8231 = n5299 & n8230;
  assign n8232 = ~Ng1988 & n8231;
  assign n8233 = ~n8229 & ~n8232;
  assign n8234 = Ng1988 & ~n8230;
  assign n8235 = ~n5300 & n8234;
  assign n2910_1 = ~n8233 | n8235;
  assign n8237 = ~Ng3171 & ~n5251;
  assign n8238 = Pg35 & ~n8237;
  assign n8239 = Ng3167 & ~n8238;
  assign n8240 = Ng3171 & n5253;
  assign n2915_1 = n8239 | n8240;
  assign n8242 = ~Pg35 & Ng843;
  assign n8243 = Ng812 & n5906;
  assign n8244 = Pg35 & Ng812;
  assign n8245 = ~n5906 & ~n8244;
  assign n8246 = Ng837 & ~n8245;
  assign n8247 = ~n8243 & n8246;
  assign n2920_1 = n8242 | n8247;
  assign n8249 = ~n7038 & n7045;
  assign n8250 = Ng832 & n8249;
  assign n8251 = ~Ng832 & n7044;
  assign n8252 = n5150 & n8251;
  assign n8253 = Pg35 & ~n8252;
  assign n8254 = Ng817 & ~n8253;
  assign n2925_1 = n8250 | n8254;
  assign n8256 = Ng5869 & n6427;
  assign n8257 = Pg35 & ~n8256;
  assign n8258 = Ng5897 & n8257;
  assign n8259 = ~Pg35 & Ng5949;
  assign n8260 = ~n5083 & ~n8259;
  assign n8261 = ~n8257 & ~n8260;
  assign n2930_1 = n8258 | n8261;
  assign n8263 = ~Pg35 & ~Ng2970;
  assign n8264 = Pg35 & ~Ng301;
  assign n8265 = n4943 & n8264;
  assign n8266 = ~Ng2902 & n8265;
  assign n2947_1 = ~n8263 & ~n8266;
  assign n8268 = Pg35 & ~Ng305;
  assign n8269 = ~Ng311 & n8268;
  assign n8270 = ~Ng26885 & n8269;
  assign n8271 = ~Ng329 & ~n8270;
  assign n8272 = Pg35 & Ng329;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = Ng305 & Ng324;
  assign n8275 = Ng311 & ~Ng324;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = Pg35 & ~n8276;
  assign n8278 = Ng336 & Ng305;
  assign n8279 = Ng311 & ~Ng336;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = ~Ng26885 & n8280;
  assign n8282 = n8277 & ~n8281;
  assign n2952_1 = n8273 | n8282;
  assign n8284 = Ng168 & n5027_1;
  assign n8285 = Ng174 & ~n5027_1;
  assign n2957_1 = n8284 | n8285;
  assign n8287 = ~Ng2461 & n8039;
  assign n8288 = ~Pg35 & Ng2811;
  assign n8289 = ~n8036 & ~n8288;
  assign n8290 = ~n7169 & ~n8289;
  assign n2962_1 = n8287 | n8290;
  assign n8292 = Pg35 & ~n5483;
  assign n8293 = Ng3684 & n8292;
  assign n8294 = ~Pg35 & Ng3614;
  assign n8295 = ~n8293 & ~n8294;
  assign n2967_1 = n5485 | ~n8295;
  assign n8297 = ~Pg35 & Ng3703;
  assign n8298 = n5413 & n5483;
  assign n8299 = Pg35 & Ng3639;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = n4540 & n7083;
  assign n8302 = ~n4541 & ~n8301;
  assign n8303 = n5483 & ~n8302;
  assign n8304 = ~n8300 & ~n8303;
  assign n2972_1 = n8297 | n8304;
  assign n8306 = ~Pg35 & Ng3329;
  assign n8307 = ~Ng3338 & ~n6653;
  assign n8308 = n6655 & ~n8307;
  assign n2980_1 = n8306 | n8308;
  assign n8310 = Pg9555 & ~Ng5456;
  assign n8311 = ~Ng5406 & ~n8310;
  assign n8312 = Pg35 & ~Pg9615;
  assign n8313 = ~n8311 & n8312;
  assign n8314 = ~Pg35 & Ng5456;
  assign n2985 = n8313 | n8314;
  assign n8316 = Ng269 & n7393;
  assign n8317 = Pg14147 & n7390;
  assign n8318 = ~Pg35 & Ng239;
  assign n8319 = ~n8317 & ~n8318;
  assign n2990_1 = n8316 | ~n8319;
  assign n8321 = Ng401 & n5151;
  assign n8322 = Ng429 & ~n5151;
  assign n2995_1 = n8321 | n8322;
  assign n8324 = ~Pg35 & Ng6035;
  assign n8325 = Pg17607 & n5217;
  assign n8326 = Pg17739 & n8325;
  assign n8327 = Ng6035 & n8326;
  assign n8328 = Pg35 & ~n8327;
  assign n8329 = ~Ng6044 & n8328;
  assign n3000_1 = n8324 | n8329;
  assign n8331 = Ng441 & n5151;
  assign n8332 = Ng475 & ~n5151;
  assign n3005_1 = n8331 | n8332;
  assign n8334 = Pg35 & \[4415] ;
  assign n8335 = ~Pg35 & Ng5062;
  assign n3010_1 = n8334 | n8335;
  assign n8337 = ~Pg35 & Ng3813;
  assign n8338 = ~Ng4054 & ~Ng3990;
  assign n8339 = Pg16659 & n8338;
  assign n8340 = Ng3953 & n8339;
  assign n8341 = ~Ng4054 & Ng3990;
  assign n8342 = Ng3921 & n8341;
  assign n8343 = Pg13966 & n8342;
  assign n8344 = ~n8340 & ~n8343;
  assign n8345 = Ng4040 & ~Pg11418;
  assign n8346 = ~Ng4040 & Pg11418;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = Pg16775 & Ng3937;
  assign n8349 = n4535 & n8348;
  assign n8350 = n8347 & ~n8349;
  assign n8351 = n8344 & n8350;
  assign n8352 = Pg16775 & Ng3945;
  assign n8353 = n8218 & n8352;
  assign n8354 = Pg13966 & Ng3929;
  assign n8355 = n8338 & n8354;
  assign n8356 = ~n8353 & ~n8355;
  assign n8357 = Ng3961 & n8341;
  assign n8358 = Pg16659 & n8357;
  assign n8359 = n8356 & ~n8358;
  assign n8360 = ~n8347 & n8359;
  assign n8361 = ~n8351 & ~n8360;
  assign n8362 = Pg16955 & Ng3925;
  assign n8363 = Ng3909 & Pg11418;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n4535 & ~n8364;
  assign n8366 = Ng3941 & n8338;
  assign n8367 = Pg13906 & n8366;
  assign n8368 = ~n8365 & ~n8367;
  assign n8369 = Ng3901 & Pg14518;
  assign n8370 = Ng4031 & Ng3913;
  assign n8371 = ~n8369 & ~n8370;
  assign n8372 = n8341 & ~n8371;
  assign n8373 = Ng3957 & Pg16748;
  assign n8374 = Ng3905 & Pg16693;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = n8218 & ~n8375;
  assign n8377 = ~Ng4040 & ~n8376;
  assign n8378 = ~n8372 & n8377;
  assign n8379 = n8368 & n8378;
  assign n8380 = Ng3889 & Pg14518;
  assign n8381 = Ng3897 & Ng4031;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = n8338 & ~n8382;
  assign n8384 = Pg16955 & Ng3917;
  assign n8385 = Pg11418 & Ng3893;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n8218 & ~n8386;
  assign n8388 = Ng4040 & ~n8387;
  assign n8389 = Ng3949 & n4535;
  assign n8390 = Pg16748 & n8389;
  assign n8391 = Pg13906 & n8341;
  assign n8392 = Ng3933 & n8391;
  assign n8393 = ~n8390 & ~n8392;
  assign n8394 = n8388 & n8393;
  assign n8395 = ~n8383 & n8394;
  assign n8396 = ~n8379 & ~n8395;
  assign n8397 = ~n8361 & ~n8396;
  assign n8398 = ~Ng3965 & n8397;
  assign n8399 = n7015 & ~n8398;
  assign n8400 = n6689 & ~n8397;
  assign n8401 = ~n7016 & ~n8400;
  assign n8402 = ~n8399 & ~n8401;
  assign n8403 = Pg35 & ~n8402;
  assign n8404 = Ng3808 & n8403;
  assign n8405 = Pg35 & ~n8401;
  assign n8406 = ~n8398 & n8405;
  assign n8407 = ~Ng3808 & n8406;
  assign n8408 = ~n8404 & ~n8407;
  assign n3014_1 = n8337 | ~n8408;
  assign n8410 = Pg35 & ~n7865;
  assign n8411 = Ng10384 & Ng4473;
  assign n8412 = ~Ng4462 & ~n8411;
  assign n3019_1 = ~n8410 | ~n8412;
  assign n8414 = n7216 & n7736;
  assign n8415 = n5018 & n8414;
  assign n8416 = ~Pg35 & ~Ng3941;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = Pg35 & ~n8414;
  assign n8419 = ~Ng3957 & n8418;
  assign n3024_1 = n8417 & ~n8419;
  assign n8421 = ~Pg35 & Ng4087;
  assign n8422 = Pg35 & Ng4093;
  assign n8423 = ~n6476 & ~n8422;
  assign n8424 = Ng2841 & ~n6477;
  assign n8425 = ~n8423 & n8424;
  assign n3029_1 = n8421 | n8425;
  assign n8427 = ~Pg35 & Ng1768;
  assign n8428 = ~Ng1760 & Ng1783;
  assign n8429 = Pg35 & ~n8428;
  assign n8430 = n6185 & n8429;
  assign n8431 = ~Ng1792 & n8430;
  assign n8432 = ~n8427 & ~n8431;
  assign n8433 = n5843 & n6186;
  assign n8434 = Pg35 & ~n6185;
  assign n8435 = Ng1760 & n8434;
  assign n8436 = ~n8433 & ~n8435;
  assign n3034_1 = ~n8432 | ~n8436;
  assign n8438 = ~Pg14779 & ~Pg17760;
  assign n8439 = ~n6873 & ~n8438;
  assign n8440 = Pg35 & ~Pg17649;
  assign n8441 = ~Pg13085 & n8440;
  assign n8442 = ~Pg17685 & n8441;
  assign n3039_1 = ~n8439 & n8442;
  assign n8444 = ~Pg35 & Ng157;
  assign n8445 = ~Ng160 & n7269;
  assign n8446 = ~n8444 & ~n8445;
  assign n8447 = ~n7269 & n7270;
  assign n8448 = Ng160 & n8447;
  assign n3043_1 = ~n8446 | n8448;
  assign n8450 = Ng2279 & n6707;
  assign n8451 = Ng2273 & ~n6707;
  assign n3048_1 = n8450 | n8451;
  assign n8453 = Ng3498 & ~n4706;
  assign n8454 = n5018 & n8453;
  assign n8455 = n5083 & ~n8453;
  assign n3053_1 = n8454 | n8455;
  assign n8457 = ~Pg35 & Ng572;
  assign n8458 = Ng586 & n5737;
  assign n8459 = ~n5749 & ~n8458;
  assign n8460 = ~n5750 & ~n8459;
  assign n3058 = n8457 | n8460;
  assign n8462 = ~Pg35 & Ng2625;
  assign n8463 = Pg35 & n5329;
  assign n8464 = Ng2610 & n8463;
  assign n8465 = ~n8462 & ~n8464;
  assign n8466 = Ng2619 & n5330;
  assign n8467 = ~n6422 & ~n8466;
  assign n3066 = ~n8465 | ~n8467;
  assign n8469 = Ng1171 & ~n6077;
  assign n8470 = ~n7748 & ~n8469;
  assign n8471 = ~n7749 & ~n8470;
  assign n3071_1 = n6578 | n8471;
  assign n8473 = ~Pg35 & Ng1600;
  assign n8474 = ~Ng1668 & Ng1636;
  assign n8475 = ~n5227 & n8474;
  assign n8476 = Pg35 & ~n8475;
  assign n8477 = ~n5237 & ~n8476;
  assign n8478 = ~n8473 & n8477;
  assign n8479 = ~Ng1608 & n8476;
  assign n3076 = ~n8478 & ~n8479;
  assign n8481 = ~Pg35 & Ng1728;
  assign n8482 = ~Ng112 & ~n4593;
  assign n8483 = Ng112 & n4593;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 = n4592 & n5058;
  assign n8486 = n8484 & n8485;
  assign n8487 = n5842 & n8486;
  assign n8488 = ~n8481 & ~n8487;
  assign n8489 = n4928 & n8485;
  assign n8490 = Ng1779 & ~n8489;
  assign n8491 = Pg35 & n8490;
  assign n3087 = ~n8488 | n8491;
  assign n8493 = Ng2638 & ~n5330;
  assign n8494 = Ng2652 & ~n5333;
  assign n8495 = ~n8493 & n8494;
  assign n8496 = n8493 & ~n8494;
  assign n3092_1 = n8495 | n8496;
  assign n8498 = ~Pg35 & ~Ng2173;
  assign n8499 = ~Ng2217 & n5258;
  assign n8500 = Ng2208 & n8499;
  assign n8501 = Ng2193 & ~n8500;
  assign n8502 = ~n6499 & n8500;
  assign n8503 = Pg35 & ~n8502;
  assign n8504 = ~n8501 & n8503;
  assign n3097 = ~n8498 & ~n8504;
  assign n8506 = ~Ng2393 & n8160;
  assign n8507 = ~Pg35 & Ng2389;
  assign n8508 = ~n7891 & ~n8507;
  assign n8509 = ~n8160 & n8508;
  assign n3102 = ~n8506 & ~n8509;
  assign n8511 = ~Ng718 & ~n6095;
  assign n8512 = ~Ng661 & n6095;
  assign n3107_1 = ~n8511 & ~n8512;
  assign n8514 = Ng4950 & n8292;
  assign n8515 = ~Ng3694 & ~Ng3703;
  assign n8516 = ~Ng3698 & Ng3703;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = Ng3639 & n8517;
  assign n8519 = ~Ng3639 & ~n8517;
  assign n8520 = ~n8518 & ~n8519;
  assign n8521 = n5483 & ~n8520;
  assign n8522 = ~Ng4950 & ~n8521;
  assign n8523 = n4609 & n4688_1;
  assign n8524 = Pg35 & n8523;
  assign n8525 = ~n8522 & n8524;
  assign n3112 = n8514 | n8525;
  assign n8527 = ~Pg35 & Ng5527;
  assign n3337_1 = Pg35 & Ng5535;
  assign n8529 = ~n5718 & n3337_1;
  assign n8530 = ~n5719 & ~n8529;
  assign n8531 = ~n6773 & ~n8530;
  assign n3117 = n8527 | n8531;
  assign n8533 = ~Pg35 & Ng2803;
  assign n3122_1 = n5978 | n8533;
  assign n8535 = ~Pg35 & Ng1345;
  assign n8536 = ~Ng1361 & ~n7248;
  assign n8537 = Pg35 & ~n7250;
  assign n8538 = ~n8536 & n8537;
  assign n3127 = n8535 | n8538;
  assign n8540 = n6227_1 & n7336;
  assign n8541 = n5083 & n8540;
  assign n8542 = ~Pg35 & Ng6227;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = Pg35 & Ng6235;
  assign n8545 = ~n8540 & n8544;
  assign n3132_1 = ~n8543 | n8545;
  assign n8547 = Pg35 & n5812;
  assign n8548 = ~Ng1099 & n8547;
  assign n8549 = Ng1152 & n5812;
  assign n8550 = Pg35 & Ng1146;
  assign n8551 = ~n8549 & n8550;
  assign n3137_1 = n8548 | n8551;
  assign n8553 = n4928 & n6421;
  assign n8554 = Ng2625 & ~n8553;
  assign n8555 = Pg35 & n8554;
  assign n8556 = ~Ng2610 & Ng2619;
  assign n8557 = Ng110 & n8556;
  assign n8558 = ~Ng110 & ~n8556;
  assign n8559 = ~n8557 & ~n8558;
  assign n8560 = n5842 & n8559;
  assign n8561 = n6421 & n8560;
  assign n8562 = ~Pg35 & Ng2610;
  assign n8563 = ~n8561 & ~n8562;
  assign n3142 = n8555 | ~n8563;
  assign n8565 = ~Pg35 & Ng164;
  assign n8566 = Ng150 & n7270;
  assign n8567 = ~n7266 & ~n8566;
  assign n8568 = ~n7267 & ~n8567;
  assign n3147 = n8565 | n8568;
  assign n8570 = Pg35 & ~n6249;
  assign n8571 = ~Ng1624 & Ng1648;
  assign n8572 = Pg35 & ~n8571;
  assign n8573 = ~n8570 & ~n8572;
  assign n8574 = ~Ng1696 & ~n8573;
  assign n8575 = Pg35 & Ng1687;
  assign n8576 = Ng1691 & n8575;
  assign n8577 = ~Ng1691 & ~n8575;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = n8573 & ~n8578;
  assign n3152_1 = ~n8574 & ~n8579;
  assign n8581 = ~Pg35 & Ng6549;
  assign n8582 = Ng6549 & ~Ng6555;
  assign n8583 = ~n7103 & ~n8582;
  assign n8584 = n7714 & ~n8583;
  assign n3157_1 = n8581 | n8584;
  assign n3162 = Pg35 & \[4431] ;
  assign n8587 = ~Pg35 & Ng3873;
  assign n8588 = n1336_1 & ~n6213;
  assign n8589 = ~n6214 & ~n8588;
  assign n8590 = ~n8021 & ~n8589;
  assign n3166 = n8587 | n8590;
  assign n8592 = n4713 & n8582;
  assign n8593 = Pg35 & ~n8592;
  assign n8594 = Ng6621 & n8593;
  assign n8595 = ~Pg35 & Ng6601;
  assign n8596 = ~n5083 & ~n8595;
  assign n8597 = ~n8593 & ~n8596;
  assign n3171_1 = n8594 | n8597;
  assign n8599 = ~Ng3470 & n5213;
  assign n8600 = Pg35 & ~Ng3470;
  assign n8601 = ~Pg35 & Ng3466;
  assign n8602 = ~n8600 & ~n8601;
  assign n8603 = ~n5213 & n8602;
  assign n3176_1 = ~n8599 & ~n8603;
  assign n8605 = Ng3869 & n6919;
  assign n8606 = Pg35 & ~n8605;
  assign n8607 = ~Pg35 & ~Ng3949;
  assign n8608 = ~n5018 & ~n8607;
  assign n8609 = ~n8606 & ~n8608;
  assign n8610 = ~Ng3897 & n8606;
  assign n3181_1 = ~n8609 & ~n8610;
  assign n8612 = Ng518 & n7910;
  assign n8613 = Ng513 & n7912;
  assign n3186 = n8612 | n8613;
  assign n8615 = ~Ng538 & ~Ng209;
  assign n3191 = Pg35 & ~n8615;
  assign n8617 = ~Pg35 & Ng2555;
  assign n8618 = ~Ng112 & ~n4568;
  assign n8619 = Ng112 & n4568;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = n4567 & n5528;
  assign n8622 = n8620 & n8621;
  assign n8623 = n5842 & n8622;
  assign n8624 = ~n8617 & ~n8623;
  assign n8625 = n4928 & n8621;
  assign n8626 = Ng2606 & ~n8625;
  assign n8627 = Pg35 & n8626;
  assign n3196 = ~n8624 | n8627;
  assign n8629 = ~Pg35 & Ng1467;
  assign n8630 = Ng1467 & n7776;
  assign n8631 = n7677 & n8630;
  assign n8632 = Ng1472 & n8631;
  assign n8633 = Pg35 & Ng1472;
  assign n8634 = ~n8631 & ~n8633;
  assign n8635 = ~n8632 & ~n8634;
  assign n3201 = n8629 | n8635;
  assign n8637 = ~Ng542 & Ng691;
  assign n8638 = n5145 & ~n8637;
  assign n8639 = ~Pg35 & Ng546;
  assign n3206 = n8638 | n8639;
  assign n8641 = ~Pg35 & Ng5180;
  assign n8642 = Ng5180 & Ng5176;
  assign n3525_1 = Pg35 & Ng5188;
  assign n8644 = ~n8642 & ~n3525_1;
  assign n8645 = ~Pg32975 & ~n5594_1;
  assign n8646 = ~n8644 & n8645;
  assign n3211_1 = n8641 | n8646;
  assign n8648 = ~Pg35 & Ng5685;
  assign n8649 = Pg17711 & n5341;
  assign n8650 = Pg17580 & n8649;
  assign n8651 = ~Ng5689 & ~n8650;
  assign n8652 = Ng5689 & n8650;
  assign n8653 = Pg35 & ~n8652;
  assign n8654 = ~n8651 & n8653;
  assign n3216 = n8648 | n8654;
  assign n8656 = Ng405 & n5151;
  assign n8657 = Ng392 & ~n5151;
  assign n3224 = n8656 | n8657;
  assign n8659 = n4708_1 & n7616;
  assign n8660 = Pg35 & ~n8659;
  assign n8661 = ~Pg35 & ~Ng5220;
  assign n8662 = ~n5018 & ~n8661;
  assign n8663 = ~n8660 & ~n8662;
  assign n8664 = ~Ng5216 & n8660;
  assign n3229_1 = ~n8663 & ~n8664;
  assign n8666 = Ng4669 & n7978;
  assign n8667 = n7977 & n7979;
  assign n8668 = ~Pg35 & Ng4664;
  assign n8669 = ~n8667 & ~n8668;
  assign n3238_1 = n8666 | ~n8669;
  assign n8671 = ~Pg35 & Ng1236;
  assign n3243_1 = n6167 | n8671;
  assign n8673 = ~Pg35 & \[4507] ;
  assign n8674 = ~Ng4311 & n4537;
  assign n8675 = Pg35 & n5189;
  assign n8676 = n8674 & n8675;
  assign n8677 = Ng4643 & ~Ng4340;
  assign n8678 = n8676 & n8677;
  assign n3248 = n8673 | n8678;
  assign n8680 = Pg35 & Ng2860;
  assign n8681 = ~Pg35 & Ng2852;
  assign n3253_1 = n8680 | n8681;
  assign n8683 = ~n6513_1 & n6903;
  assign n8684 = Pg35 & ~n8683;
  assign n8685 = ~Ng4749 & ~n8684;
  assign n8686 = ~Ng4743 & ~n6903;
  assign n8687 = ~n5669 & ~n8686;
  assign n8688 = n6519 & ~n8687;
  assign n3258 = ~n8685 & ~n8688;
  assign n8690 = ~Ng6549 & ~Ng6561;
  assign n8691 = ~Ng6555 & n8690;
  assign n8692 = n7557 & n8691;
  assign n8693 = n5083 & n8692;
  assign n8694 = ~Pg35 & Ng6597;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = Pg35 & Ng6593;
  assign n8697 = ~n8692 & n8696;
  assign n3263_1 = ~n8695 | n8697;
  assign n8699 = Pg35 & Ng218;
  assign n8700 = ~Pg35 & ~Ng209;
  assign n3268 = ~n8699 & ~n8700;
  assign n8702 = ~Pg35 & Ng1542;
  assign n8703 = Ng1339 & Ng1521;
  assign n8704 = ~Ng1532 & n8703;
  assign n8705 = Pg7946 & ~n8704;
  assign n8706 = n6435 & n8705;
  assign n8707 = Ng1542 & n8706;
  assign n8708 = Pg35 & Ng1413;
  assign n8709 = ~n8707 & ~n8708;
  assign n8710 = Ng1345 & Ng1379;
  assign n8711 = Ng1367 & n8710;
  assign n8712 = ~n5509 & n8711;
  assign n8713 = n4822 & ~n8712;
  assign n8714 = Pg7946 & ~n8713;
  assign n8715 = n8704 & n8714;
  assign n8716 = Ng1536 & ~n6435;
  assign n8717 = n8715 & ~n8716;
  assign n8718 = Ng1413 & n8707;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n8709 & n8719;
  assign n3276_1 = n8702 | n8720;
  assign n8722 = n7556 & n7753;
  assign n8723 = n5018 & n8722;
  assign n8724 = ~Pg35 & ~Ng6625;
  assign n8725 = ~n8723 & ~n8724;
  assign n8726 = Pg35 & ~n8722;
  assign n8727 = ~Ng6641 & n8726;
  assign n3287_1 = n8725 & ~n8727;
  assign n8729 = Ng1936 & n5873;
  assign n8730 = Pg35 & n5875;
  assign n8731 = Ng1906 & ~n8730;
  assign n8732 = ~n5873 & n8731;
  assign n3292_1 = n8729 | n8732;
  assign n8734 = ~Ng499 & n7912;
  assign n8735 = ~Ng504 & n7910;
  assign n3302_1 = ~n8734 & ~n8735;
  assign n8737 = ~Pg35 & Ng2595;
  assign n8738 = n5332 & n8111;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = Ng2587 & n5330;
  assign n8741 = ~n6422 & ~n8740;
  assign n3307 = ~n8739 | ~n8741;
  assign n8743 = ~Pg35 & Ng4477;
  assign n8744 = Ng4581 & n6134;
  assign n8745 = ~Ng4372 & ~Ng4581;
  assign n8746 = Pg35 & ~n8745;
  assign n8747 = ~n8744 & n8746;
  assign n8748 = ~n7451 & ~n8747;
  assign n3312 = n8743 | ~n8748;
  assign n8750 = ~Pg35 & ~Ng2315;
  assign n8751 = ~Ng2287 & Ng2331;
  assign n8752 = ~n4978 & n8751;
  assign n8753 = ~n4985 & n8752;
  assign n8754 = Ng2311 & ~n8752;
  assign n8755 = Pg35 & ~n8754;
  assign n8756 = ~n8753 & n8755;
  assign n3317_1 = ~n8750 & ~n8756;
  assign n8758 = ~Pg35 & ~Ng3586;
  assign n8759 = n5032_1 & n5634;
  assign n8760 = ~n5018 & n8759;
  assign n8761 = Pg35 & ~Ng3602;
  assign n8762 = ~n8759 & ~n8761;
  assign n8763 = ~n8760 & ~n8762;
  assign n3322_1 = ~n8758 & ~n8763;
  assign n8765 = n5374 & n7624;
  assign n8766 = n5018 & n8765;
  assign n8767 = ~Pg35 & ~Ng5543;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = Pg35 & ~n8765;
  assign n8770 = ~Ng5571 & n8769;
  assign n3327_1 = n8768 & ~n8770;
  assign n8772 = n4705 & n5200;
  assign n8773 = n5083 & n8772;
  assign n8774 = ~Pg35 & Ng3558;
  assign n8775 = ~n8773 & ~n8774;
  assign n8776 = Pg35 & Ng3578;
  assign n8777 = ~n8772 & n8776;
  assign n3332 = ~n8775 | n8777;
  assign n8779 = Ng5827 & n6560;
  assign n8780 = Ng5821 & ~n6560;
  assign n3341_1 = n8779 | n8780;
  assign n8782 = n5201 & n5635;
  assign n8783 = n5018 & n8782;
  assign n8784 = ~Pg35 & ~Ng3566;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = Pg35 & ~n8782;
  assign n8787 = ~Ng3582 & n8786;
  assign n3346_1 = n8785 & ~n8787;
  assign n8789 = ~Pg35 & ~Ng6247;
  assign n8790 = n5498 & n6386;
  assign n8791 = Pg35 & ~Ng6271;
  assign n8792 = ~n8790 & n8791;
  assign n8793 = n5018 & n8790;
  assign n8794 = ~n8792 & ~n8793;
  assign n3351_1 = ~n8789 & n8794;
  assign n3356 = Ng4681 & ~n5864;
  assign n8797 = Ng2380 & n4981;
  assign n8798 = Ng2375 & ~n4981;
  assign n3361_1 = n8797 | n8798;
  assign n8800 = ~Pg35 & Ng5188;
  assign n8801 = n5820 & n7616;
  assign n8802 = n5083 & n8801;
  assign n8803 = Pg35 & Ng5196;
  assign n8804 = ~n8801 & n8803;
  assign n8805 = ~n8802 & ~n8804;
  assign n3366 = n8800 | ~n8805;
  assign n8807 = Ng3155 & ~Ng3161;
  assign n8808 = n4730 & n8807;
  assign n8809 = n5083 & n8808;
  assign n8810 = ~Pg35 & Ng3207;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = Pg35 & Ng3227;
  assign n8813 = ~n8808 & n8812;
  assign n3371_1 = ~n8811 | n8813;
  assign n8815 = ~Pg35 & ~Ng2024;
  assign n8816 = Ng2040 & ~Ng1996;
  assign n8817 = ~n5660 & n8816;
  assign n8818 = ~n6911 & n8817;
  assign n8819 = Ng2020 & ~n8817;
  assign n8820 = Pg35 & ~n8819;
  assign n8821 = ~n8818 & n8820;
  assign n3376 = ~n8815 & ~n8821;
  assign n8823 = Ng6541 & ~n4714;
  assign n8824 = n5018 & n8823;
  assign n8825 = n5083 & ~n8823;
  assign n3387 = n8824 | n8825;
  assign n8827 = ~Ng3179 & n6988;
  assign n8828 = Pg35 & ~n8827;
  assign n8829 = Ng3203 & n8828;
  assign n8830 = ~Pg35 & Ng3251;
  assign n8831 = ~n5083 & ~n8830;
  assign n8832 = ~n8828 & ~n8831;
  assign n3392_1 = n8829 | n8832;
  assign n8834 = Ng1668 & n5244;
  assign n8835 = n4575_1 & n5089;
  assign n8836 = Pg35 & n8835;
  assign n8837 = Ng1636 & ~n8836;
  assign n8838 = ~n5244 & n8837;
  assign n3397_1 = n8834 | n8838;
  assign n8840 = Ng4760 & n6856;
  assign n8841 = ~Ng6040 & ~Ng6049;
  assign n8842 = ~Ng6044 & Ng6049;
  assign n8843 = ~n8841 & ~n8842;
  assign n8844 = Ng5990 & n8843;
  assign n8845 = ~Ng5990 & ~n8843;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = n6556_1 & ~n8846;
  assign n8848 = ~Ng4760 & ~n8847;
  assign n8849 = Pg35 & n6512;
  assign n8850 = ~n8848 & n8849;
  assign n3402_1 = n8840 | n8850;
  assign n8852 = Pg14096 & n7390;
  assign n8853 = ~Pg35 & Ng232;
  assign n8854 = Ng262 & n7393;
  assign n8855 = ~n8853 & ~n8854;
  assign n3407 = n8852 | ~n8855;
  assign n8857 = Pg35 & ~n7848;
  assign n8858 = ~n5087 & ~n8857;
  assign n8859 = Ng1834 & n8858;
  assign n8860 = Ng1840 & ~n8858;
  assign n3412_1 = n8859 | n8860;
  assign n8862 = Ng5467 & n7205;
  assign n8863 = Ng5503 & ~n7205;
  assign n3417_1 = n8862 | n8863;
  assign n8865 = ~Ng370 & n6740;
  assign n8866 = Ng246 & n8865;
  assign n8867 = Ng460 & n5027_1;
  assign n8868 = ~Pg35 & Ng168;
  assign n8869 = ~n8867 & ~n8868;
  assign n3422 = n8866 | ~n8869;
  assign n8871 = ~Pg35 & Ng6203;
  assign n8872 = ~n5497 & ~n6386;
  assign n8873 = n5110 & ~n8872;
  assign n3427_1 = n8871 | n8873;
  assign n8875 = ~\[4436]  & n7128;
  assign n8876 = Pg35 & Ng333;
  assign n8877 = ~n7128 & ~n8876;
  assign n8878 = ~Ng355 & n8877;
  assign n3432 = ~n8875 & ~n8878;
  assign n8880 = Ng655 & n6095;
  assign n8881 = Ng650 & ~n6095;
  assign n3440_1 = n8880 | n8881;
  assign n3445 = Pg35 & Ng3502;
  assign n8884 = n4589 & n6494;
  assign n8885 = n4928 & n8884;
  assign n8886 = Pg35 & Ng2204;
  assign n8887 = ~n8885 & n8886;
  assign n8888 = Ng112 & n4590;
  assign n8889 = ~Ng112 & ~n4590;
  assign n8890 = ~n8888 & ~n8889;
  assign n8891 = n5842 & n8890;
  assign n8892 = n8884 & n8891;
  assign n8893 = ~Pg35 & Ng2153;
  assign n8894 = ~n8892 & ~n8893;
  assign n3450_1 = n8887 | ~n8894;
  assign n8896 = n5820 & n6412;
  assign n8897 = Pg35 & ~n8896;
  assign n8898 = Ng5256 & n8897;
  assign n8899 = ~Pg35 & Ng5240;
  assign n8900 = ~n5083 & ~n8899;
  assign n8901 = ~n8897 & ~n8900;
  assign n3455_1 = n8898 | n8901;
  assign n8903 = Ng4601 & n5569;
  assign n8904 = n5568 & n8903;
  assign n8905 = ~Ng4608 & n8904;
  assign n8906 = n7476 & ~n8903;
  assign n8907 = Ng4608 & n8906;
  assign n8908 = ~Pg35 & Ng4601;
  assign n8909 = ~n8907 & ~n8908;
  assign n3460 = n8905 | ~n8909;
  assign n8911 = ~Pg35 & Ng790;
  assign n8912 = Ng794 & n5145;
  assign n8913 = ~n5142 & ~n8912;
  assign n8914 = ~n5143 & ~n8913;
  assign n3465_1 = n8911 | n8914;
  assign n8916 = ~Pg35 & Ng3680;
  assign n8917 = ~Ng3689 & ~n5284;
  assign n8918 = Pg35 & ~n5285;
  assign n8919 = ~n8917 & n8918;
  assign n3477_1 = n8916 | n8919;
  assign n8921 = Pg35 & ~Ng703;
  assign n8922 = n6741 & n7042;
  assign n8923 = Ng837 & n8922;
  assign n8924 = ~n8921 & ~n8923;
  assign n8925 = Ng822 & Ng723;
  assign n8926 = n7038 & n8925;
  assign n8927 = ~Ng847 & n8926;
  assign n8928 = ~n8924 & ~n8927;
  assign n8929 = ~Pg35 & ~Ng847;
  assign n3486 = ~n8928 & ~n8929;
  assign n8931 = ~Pg35 & Ng890;
  assign n8932 = Ng890 & Ng896;
  assign n8933 = Pg35 & ~n8932;
  assign n8934 = ~n7388 & n8933;
  assign n3491_1 = n8931 | n8934;
  assign n8936 = ~Pg35 & ~Ng3231;
  assign n8937 = n5396 & n7522;
  assign n8938 = Pg35 & ~Ng3247;
  assign n8939 = ~n8937 & n8938;
  assign n8940 = n5018 & n8937;
  assign n8941 = ~n8939 & ~n8940;
  assign n3496 = ~n8936 & n8941;
  assign n8943 = ~Pg35 & Ng2047;
  assign n8944 = Ng2040 & n5661;
  assign n8945 = n4595 & n5089;
  assign n8946 = Pg35 & ~n8945;
  assign n8947 = n8013 & n8946;
  assign n8948 = ~n8944 & ~n8947;
  assign n3501_1 = n8943 | ~n8948;
  assign n8950 = ~Pg35 & ~Ng4176;
  assign n8951 = Pg35 & ~Ng4146;
  assign n3506 = ~n8950 & ~n8951;
  assign n8953 = n5310 & n5312;
  assign n8954 = ~Ng4633 & n8953;
  assign n8955 = Pg35 & ~n8954;
  assign n8956 = Ng4628 & ~n8955;
  assign n8957 = Ng4628 & ~n5313;
  assign n8958 = n5311 & ~n8957;
  assign n8959 = Ng4633 & n8958;
  assign n3511_1 = n8956 | n8959;
  assign n8961 = n4824 & n7062;
  assign n8962 = Ng979 & Ng1236;
  assign n8963 = ~Ng979 & ~Ng1236;
  assign n8964 = Pg35 & ~n8963;
  assign n8965 = ~n8962 & n8964;
  assign n8966 = n8961 & n8965;
  assign n8967 = ~Pg8416 & n6939;
  assign n8968 = ~Pg13259 & n8967;
  assign n8969 = n8966 & n8968;
  assign n8970 = Pg35 & n8968;
  assign n8971 = ~Pg35 & Ng996;
  assign n8972 = ~n8970 & ~n8971;
  assign n8973 = ~n8966 & n8972;
  assign n3516_1 = ~n8969 & ~n8973;
  assign n8975 = Pg35 & Ng4732;
  assign n8976 = ~Pg35 & Ng4727;
  assign n3520_1 = n8975 | n8976;
  assign n8978 = Ng5817 & n6560;
  assign n8979 = Pg35 & Ng5813;
  assign n8980 = ~Ng5808 & n8979;
  assign n8981 = Ng5808 & ~n8979;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = ~n6560 & ~n8982;
  assign n3529_1 = n8978 | n8983;
  assign n8985 = ~Pg35 & Ng2357;
  assign n8986 = Ng2342 & n7690;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = Ng2351 & n7142;
  assign n8989 = ~n7146 & ~n8988;
  assign n3534_1 = ~n8987 | ~n8989;
  assign n8991 = ~Ng2629 & ~Ng2555;
  assign n8992 = Pg35 & ~n8991;
  assign n8993 = ~n7668 & ~n8992;
  assign n8994 = Ng2643 & n8993;
  assign n8995 = Ng2648 & ~n8993;
  assign n3539_1 = n8994 | n8995;
  assign n8997 = Pg35 & n6465;
  assign n3544 = Ng6732 & ~n8997;
  assign n8999 = ~n5670 & n8523;
  assign n9000 = Pg35 & ~n8999;
  assign n9001 = ~Ng4950 & ~n9000;
  assign n9002 = ~Ng4944 & ~n8523;
  assign n9003 = ~n5669 & ~n9002;
  assign n9004 = n5677 & ~n9003;
  assign n3549 = ~n9001 & ~n9004;
  assign n9006 = ~Pg35 & Ng4125;
  assign n9007 = n4521 & n4527;
  assign n9008 = Ng4076 & Ng4087;
  assign n9009 = n4712 & n9008;
  assign n9010 = n9007 & n9009;
  assign n9011 = n6197_1 & ~n9010;
  assign n3554_1 = n9006 | n9011;
  assign n9013 = ~Pg35 & ~Ng333;
  assign n3559 = ~n6750 & ~n9013;
  assign n9015 = Pg35 & Ng3462;
  assign n9016 = ~Ng3457 & ~n9015;
  assign n9017 = Ng3457 & n9015;
  assign n9018 = ~n9016 & ~n9017;
  assign n9019 = ~n7361 & n9018;
  assign n9020 = Ng3466 & n7361;
  assign n3567_1 = n9019 | n9020;
  assign n9022 = ~Ng4076 & n4523;
  assign n9023 = n4521 & n9022;
  assign n9024 = Ng4064 & ~Ng4057;
  assign n9025 = n9023 & n9024;
  assign n9026 = Pg35 & ~n9025;
  assign n9027 = Ng4116 & n9026;
  assign n9028 = ~Pg35 & Ng4112;
  assign n9029 = Pg35 & Ng4145;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = ~n9026 & ~n9030;
  assign n3572_1 = n9027 | n9031;
  assign n9033 = ~n4903 & ~n4910;
  assign n9034 = Pg35 & ~Ng5041;
  assign n9035 = ~n9033 & n9034;
  assign n9036 = ~Pg35 & Ng5037;
  assign n9037 = ~n9035 & ~n9036;
  assign n9038 = n7591 & n9033;
  assign n9039 = Ng5041 & n9038;
  assign n3577_1 = ~n9037 | n9039;
  assign n9041 = n6864 & n7403;
  assign n9042 = Ng4430 & n9041;
  assign n3582 = Ng4452 | n9042;
  assign n9044 = Ng3827 & n7017;
  assign n9045 = Ng3821 & ~n7017;
  assign n3587_1 = n9044 | n9045;
  assign n9047 = ~Pg35 & Ng6505;
  assign n9048 = ~Ng6682 & ~Ng6741;
  assign n9049 = Ng6645 & Pg17688;
  assign n9050 = n9048 & n9049;
  assign n9051 = ~Ng6727 & ~Pg12470;
  assign n9052 = Ng6727 & Pg12470;
  assign n9053 = ~n9051 & ~n9052;
  assign n9054 = Ng6682 & ~Ng6741;
  assign n9055 = Ng6613 & Pg14828;
  assign n9056 = n9054 & n9055;
  assign n9057 = ~n9053 & ~n9056;
  assign n9058 = Pg17778 & n4538;
  assign n9059 = Ng6629 & n9058;
  assign n9060 = n9057 & ~n9059;
  assign n9061 = ~n9050 & n9060;
  assign n9062 = ~Ng6682 & Ng6741;
  assign n9063 = Ng6637 & Pg17778;
  assign n9064 = n9062 & n9063;
  assign n9065 = Pg17688 & n9054;
  assign n9066 = Ng6653 & n9065;
  assign n9067 = Ng6621 & Pg14828;
  assign n9068 = n9048 & n9067;
  assign n9069 = ~n9066 & ~n9068;
  assign n9070 = n9053 & n9069;
  assign n9071 = ~n9064 & n9070;
  assign n9072 = ~n9061 & ~n9071;
  assign n9073 = Pg13099 & Ng6593;
  assign n9074 = Ng6723 & Ng6605;
  assign n9075 = ~n9073 & ~n9074;
  assign n9076 = n9054 & ~n9075;
  assign n9077 = Ng6633 & n9048;
  assign n9078 = Pg14749 & n9077;
  assign n9079 = ~n9076 & ~n9078;
  assign n9080 = Ng6649 & Pg17764;
  assign n9081 = Ng6597 & Pg17722;
  assign n9082 = ~n9080 & ~n9081;
  assign n9083 = n9062 & ~n9082;
  assign n9084 = Pg17871 & Ng6617;
  assign n9085 = Pg12470 & Ng6601;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = n4538 & ~n9086;
  assign n9088 = ~Ng6727 & ~n9087;
  assign n9089 = ~n9083 & n9088;
  assign n9090 = n9079 & n9089;
  assign n9091 = Pg13099 & Ng6581;
  assign n9092 = Ng6589 & Ng6723;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = n9048 & ~n9093;
  assign n9095 = Ng6641 & Pg17764;
  assign n9096 = n4538 & n9095;
  assign n9097 = Ng6727 & ~n9096;
  assign n9098 = Ng6609 & Pg17871;
  assign n9099 = Ng6585 & Pg12470;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = n9062 & ~n9100;
  assign n9102 = Pg14749 & n9054;
  assign n9103 = Ng6625 & n9102;
  assign n9104 = ~n9101 & ~n9103;
  assign n9105 = n9097 & n9104;
  assign n9106 = ~n9094 & n9105;
  assign n9107 = ~n9090 & ~n9106;
  assign n9108 = ~n9072 & ~n9107;
  assign n9109 = ~Ng6657 & n9108;
  assign n9110 = n7838 & ~n9109;
  assign n9111 = n7836 & ~n9108;
  assign n9112 = ~n7839 & ~n9111;
  assign n9113 = ~n9110 & ~n9112;
  assign n9114 = Pg35 & ~n9113;
  assign n9115 = Ng6500 & n9114;
  assign n9116 = Pg35 & ~n9112;
  assign n9117 = ~n9109 & n9116;
  assign n9118 = ~Ng6500 & n9117;
  assign n9119 = ~n9115 & ~n9118;
  assign n3592 = n9047 | ~n9119;
  assign n9121 = Ng3338 & n4532;
  assign n9122 = Pg16624 & n9121;
  assign n9123 = n7880 & n9122;
  assign n9124 = Pg35 & ~n9123;
  assign n9125 = ~Ng3133 & n9124;
  assign n9126 = ~Pg35 & Ng3129;
  assign n9127 = ~n6640 & ~n9126;
  assign n9128 = ~n9124 & n9127;
  assign n3600 = ~n9125 & ~n9128;
  assign n9130 = Pg35 & ~n7880;
  assign n9131 = Ng3333 & n9130;
  assign n9132 = Pg16718 & n4532;
  assign n9133 = Ng3235 & n9132;
  assign n9134 = Ng3288 & ~Ng3352;
  assign n9135 = Pg13895 & Ng3219;
  assign n9136 = n9134 & n9135;
  assign n9137 = ~n9133 & ~n9136;
  assign n9138 = ~Ng3288 & ~Ng3352;
  assign n9139 = Pg16603 & Ng3251;
  assign n9140 = n9138 & n9139;
  assign n9141 = Ng3338 & ~Pg11349;
  assign n9142 = ~Ng3338 & Pg11349;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 = ~n9140 & n9143;
  assign n9145 = n9137 & n9144;
  assign n9146 = ~Ng3288 & Ng3352;
  assign n9147 = Ng3243 & Pg16718;
  assign n9148 = n9146 & n9147;
  assign n9149 = Ng3259 & Pg16603;
  assign n9150 = n9134 & n9149;
  assign n9151 = ~n9143 & ~n9150;
  assign n9152 = Ng3227 & n9138;
  assign n9153 = Pg13895 & n9152;
  assign n9154 = n9151 & ~n9153;
  assign n9155 = ~n9148 & n9154;
  assign n9156 = ~n9145 & ~n9155;
  assign n9157 = Ng3247 & n4532;
  assign n9158 = Pg16686 & n9157;
  assign n9159 = Ng3231 & n9134;
  assign n9160 = Pg13865 & n9159;
  assign n9161 = ~n9158 & ~n9160;
  assign n9162 = Pg16874 & Ng3215;
  assign n9163 = Pg11349 & Ng3191;
  assign n9164 = ~n9162 & ~n9163;
  assign n9165 = n9146 & ~n9164;
  assign n9166 = Pg14421 & Ng3187;
  assign n9167 = Ng3195 & Ng3329;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = n9138 & ~n9168;
  assign n9170 = Ng3338 & ~n9169;
  assign n9171 = ~n9165 & n9170;
  assign n9172 = n9161 & n9171;
  assign n9173 = Ng3239 & n9138;
  assign n9174 = Pg13865 & n9173;
  assign n9175 = Pg16874 & Ng3223;
  assign n9176 = Pg11349 & Ng3207;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = n4532 & ~n9177;
  assign n9179 = ~Ng3338 & ~n9178;
  assign n9180 = Pg14421 & Ng3199;
  assign n9181 = Ng3329 & Ng3211;
  assign n9182 = ~n9180 & ~n9181;
  assign n9183 = n9134 & ~n9182;
  assign n9184 = Ng3255 & Pg16686;
  assign n9185 = Ng3203 & Pg16624;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = n9146 & ~n9186;
  assign n9188 = ~n9183 & ~n9187;
  assign n9189 = n9179 & n9188;
  assign n9190 = ~n9174 & n9189;
  assign n9191 = ~n9172 & ~n9190;
  assign n9192 = ~n9156 & ~n9191;
  assign n9193 = ~Ng3263 & n9192;
  assign n9194 = ~n9122 & n9192;
  assign n9195 = Pg35 & n7880;
  assign n9196 = ~n9194 & n9195;
  assign n9197 = ~n9193 & n9196;
  assign n9198 = ~Pg35 & Ng3263;
  assign n9199 = ~n9197 & ~n9198;
  assign n3605 = n9131 | ~n9199;
  assign n3614 = Ng4674 & ~n5864;
  assign n9202 = ~Pg35 & Ng294;
  assign n9203 = Ng298 & n5713;
  assign n9204 = ~n5712 & ~n9203;
  assign n9205 = ~n6927 & ~n9204;
  assign n3619_1 = n9202 | n9205;
  assign n9207 = Ng2661 & n8993;
  assign n9208 = Ng2667 & ~n8993;
  assign n3624_1 = n9207 | n9208;
  assign n9210 = ~Pg35 & Ng1902;
  assign n9211 = Ng1917 & ~Ng1894;
  assign n9212 = Pg35 & ~n9211;
  assign n9213 = n5297 & n9212;
  assign n9214 = ~Ng1926 & n9213;
  assign n9215 = ~n9210 & ~n9214;
  assign n9216 = Ng1894 & n5838;
  assign n9217 = ~n5844 & ~n9216;
  assign n3632 = ~n9215 | ~n9217;
  assign n9219 = Pg35 & Ng2988;
  assign n9220 = ~Pg35 & Ng2994;
  assign n3637 = n9219 | n9220;
  assign n9222 = n5034 & n5635;
  assign n9223 = n5083 & n9222;
  assign n9224 = ~Pg35 & Ng3530;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = Pg35 & Ng3538;
  assign n9227 = ~n9222 & n9226;
  assign n3642_1 = ~n9225 | n9227;
  assign n9229 = Pg35 & ~n7269;
  assign n3647_1 = Ng160 & ~n9229;
  assign n9231 = Pg35 & Ng316;
  assign n9232 = ~Pg35 & \[4431] ;
  assign n3652_1 = n9231 | n9232;
  assign n9234 = Ng827 & n7046;
  assign n9235 = n7039 & n7044;
  assign n9236 = ~Ng827 & n9235;
  assign n9237 = Pg35 & ~n9236;
  assign n9238 = Ng822 & ~n9237;
  assign n3657_1 = n9234 | n9238;
  assign n9240 = n7502 & ~n8961;
  assign n9241 = Pg35 & ~Pg17291;
  assign n9242 = ~Pg17316 & ~Pg17400;
  assign n9243 = n9241 & n9242;
  assign n3662 = ~n9240 & n9243;
  assign n9245 = Ng2555 & n7668;
  assign n9246 = ~Ng2555 & ~n5534;
  assign n9247 = ~Ng2629 & n7672;
  assign n9248 = ~n9246 & n9247;
  assign n3666 = n9245 | n9248;
  assign n9250 = Pg35 & ~n7836;
  assign n9251 = Ng5011 & n9250;
  assign n9252 = ~Pg35 & Ng6657;
  assign n9253 = ~n9251 & ~n9252;
  assign n3671 = n9117 | ~n9253;
  assign n9255 = ~Ng222 & ~Ng199;
  assign n9256 = Pg35 & n9255;
  assign n9257 = ~Pg35 & ~\[4426] ;
  assign n3676_1 = ~n9256 & ~n9257;
  assign n9259 = Ng6523 & n7840;
  assign n9260 = Pg35 & ~Ng6513;
  assign n9261 = n7839 & n9260;
  assign n9262 = ~Ng6519 & n9261;
  assign n9263 = ~n9259 & ~n9262;
  assign n9264 = Ng6519 & ~n9260;
  assign n9265 = ~n7840 & n9264;
  assign n3681_1 = ~n9263 | n9265;
  assign n9267 = Pg7946 & Ng1514;
  assign n9268 = Ng1526 & ~n9267;
  assign n9269 = ~n8717 & ~n9268;
  assign n9270 = Pg35 & ~n9269;
  assign n9271 = Pg7946 & ~Ng1526;
  assign n9272 = Pg35 & ~n9271;
  assign n9273 = Ng1514 & ~n9272;
  assign n3686_1 = n9270 | n9273;
  assign n9275 = ~Ng4601 & ~n5569;
  assign n9276 = n8906 & ~n9275;
  assign n9277 = ~Pg35 & Ng4593;
  assign n3691 = n9276 | n9277;
  assign n9279 = ~Ng437 & ~Ng405;
  assign n9280 = ~Ng401 & Ng405;
  assign n9281 = Ng392 & ~n9280;
  assign n9282 = ~n9279 & n9281;
  assign n9283 = ~Ng405 & ~Ng424;
  assign n9284 = ~Ng437 & Ng405;
  assign n9285 = ~n9283 & ~n9284;
  assign n9286 = ~Ng392 & n9285;
  assign n9287 = ~n9282 & ~n9286;
  assign n9288 = Ng417 & n9287;
  assign n9289 = Ng370 & n5807_1;
  assign n9290 = ~Ng385 & n9289;
  assign n9291 = ~n9288 & n9290;
  assign n9292 = Ng441 & Ng392;
  assign n9293 = ~Ng392 & Ng411;
  assign n9294 = ~Ng691 & ~n9293;
  assign n9295 = ~n9292 & n9294;
  assign n9296 = Ng452 & Ng392;
  assign n9297 = Ng174 & ~Ng392;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = ~Ng182 & n9298;
  assign n9300 = Ng182 & ~n9298;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = n9295 & n9301;
  assign n9303 = ~Ng417 & ~n9287;
  assign n9304 = ~n9302 & n9303;
  assign n9305 = n9291 & ~n9304;
  assign n9306 = Ng854 & ~n9290;
  assign n9307 = ~n9305 & ~n9306;
  assign n3696 = Pg35 & ~n9307;
  assign n9309 = ~Ng1484 & ~n6276_1;
  assign n9310 = Pg35 & n6265;
  assign n9311 = ~Ng1300 & n6271_1;
  assign n9312 = Ng1300 & ~n6271_1;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = n9310 & ~n9313;
  assign n9315 = ~n9309 & n9314;
  assign n9316 = ~Pg35 & Ng1472;
  assign n9317 = Ng1484 & n6266_1;
  assign n9318 = ~n9316 & ~n9317;
  assign n3701 = n9315 | ~n9318;
  assign n9320 = Pg35 & Ng4922;
  assign n9321 = ~Pg35 & Ng4917;
  assign n3706_1 = n9320 | n9321;
  assign n9323 = ~Pg35 & Ng5077;
  assign n9324 = Ng5077 & ~Ng5069;
  assign n9325 = Ng5084 & ~n9324;
  assign n9326 = Ng5077 & ~Ng5073;
  assign n9327 = ~Ng5084 & ~n9326;
  assign n9328 = ~n9325 & ~n9327;
  assign n3711 = n9323 | n9328;
  assign n9330 = ~Pg35 & Ng5857;
  assign n9331 = ~n6426 & ~n7650;
  assign n9332 = n7580 & ~n9331;
  assign n3716_1 = n9330 | n9332;
  assign n9334 = ~Ng10384 & n7858;
  assign n9335 = ~Pg35 & Ng4462;
  assign n3721_1 = n9334 | n9335;
  assign n9337 = Ng2504 & ~n6149;
  assign n9338 = Ng2476 & ~Ng2453;
  assign n9339 = Pg35 & ~n9338;
  assign n9340 = ~n6149 & ~n9339;
  assign n9341 = Ng2518 & ~n9340;
  assign n9342 = ~n9337 & n9341;
  assign n9343 = n9337 & ~n9341;
  assign n3726 = n9342 | n9343;
  assign n9345 = ~Pg35 & Ng2648;
  assign n9346 = ~n5543 & ~n9345;
  assign n9347 = n8993 & n9346;
  assign n9348 = ~Ng2567 & ~n8993;
  assign n3731_1 = ~n9347 & ~n9348;
  assign n9350 = ~Pg35 & Ng562;
  assign n9351 = Ng568 & n5737;
  assign n9352 = ~n5747 & ~n9351;
  assign n9353 = ~n5748 & ~n9352;
  assign n3736_1 = n9350 | n9353;
  assign n9355 = Ng3263 & n5955;
  assign n9356 = ~Pg35 & Ng3259;
  assign n9357 = ~n5083 & ~n9356;
  assign n9358 = ~n5955 & ~n9357;
  assign n3741_1 = n9355 | n9358;
  assign n9360 = n7380 & n8582;
  assign n9361 = Pg35 & ~n9360;
  assign n9362 = ~Pg35 & ~Ng6585;
  assign n9363 = ~n5018 & ~n9362;
  assign n9364 = ~n9361 & ~n9363;
  assign n9365 = ~Ng6613 & n9361;
  assign n3746 = ~n9364 & ~n9365;
  assign n9367 = Pg35 & n8327;
  assign n3751 = Ng6040 & ~n9367;
  assign n9369 = ~Ng6494 & Pg9743;
  assign n9370 = ~Ng6444 & ~n9369;
  assign n9371 = Pg35 & ~Pg9817;
  assign n9372 = ~n9370 & n9371;
  assign n9373 = ~Pg35 & Ng6494;
  assign n3756 = n9372 | n9373;
  assign n9375 = ~Pg35 & ~Ng2955;
  assign n9376 = n4863 & ~n4871;
  assign n9377 = Pg91 & Pg35;
  assign n9378 = ~Ng2965 & n9377;
  assign n9379 = n9376 & n9378;
  assign n3761_1 = ~n9375 & ~n9379;
  assign n3766_1 = ~Ng5857 & n7581;
  assign n9382 = ~Pg35 & Ng1620;
  assign n9383 = Pg35 & ~n6253;
  assign n9384 = ~n5244 & ~n9383;
  assign n9385 = n5237 & n9384;
  assign n9386 = Ng1616 & ~n9384;
  assign n9387 = ~n9385 & ~n9386;
  assign n3771_1 = n9382 | ~n9387;
  assign n9389 = ~Pg35 & ~Ng446;
  assign n9390 = ~Ng703 & n9305;
  assign n9391 = ~n5808 & ~n9390;
  assign n9392 = Ng896 & ~n9391;
  assign n9393 = Ng862 & ~n9392;
  assign n9394 = n8933 & ~n9393;
  assign n3776_1 = ~n9389 & ~n9394;
  assign n9396 = Ng3518 & n5828;
  assign n9397 = Pg35 & ~n9396;
  assign n9398 = ~Pg35 & ~Ng3606;
  assign n9399 = ~n5018 & ~n9398;
  assign n9400 = ~n9397 & ~n9399;
  assign n9401 = ~Ng3562 & n9397;
  assign n3784_1 = ~n9400 & ~n9401;
  assign n9403 = ~Ng4297 & ~Pg10122;
  assign n9404 = Pg35 & n9403;
  assign n9405 = ~Pg35 & Ng4239;
  assign n3789_1 = n9404 | n9405;
  assign n9407 = ~Pg35 & Ng1395;
  assign n9408 = Pg35 & ~Ng1322;
  assign n9409 = Pg12923 & ~n5518;
  assign n9410 = Ng1395 & n9409;
  assign n9411 = ~Ng1404 & n9410;
  assign n9412 = Ng1404 & ~n9410;
  assign n9413 = ~n9411 & ~n9412;
  assign n9414 = n9408 & ~n9413;
  assign n3793_1 = n9407 | n9414;
  assign n9416 = Pg35 & Ng3813;
  assign n9417 = Ng3808 & n9416;
  assign n9418 = ~Ng3808 & ~n9416;
  assign n9419 = ~n9417 & ~n9418;
  assign n9420 = ~n7017 & ~n9419;
  assign n9421 = ~Ng3817 & n7017;
  assign n3798_1 = ~n9420 & ~n9421;
  assign n9423 = Ng4498 & ~n5406;
  assign n9424 = ~n6976 & ~n9423;
  assign n3808 = n7572 | ~n9424;
  assign n9426 = ~Ng287 & n5708;
  assign n9427 = Pg35 & ~n9426;
  assign n9428 = Ng283 & ~n9427;
  assign n9429 = ~Ng283 & n5713;
  assign n9430 = Ng287 & n9429;
  assign n3813_1 = n9428 | n9430;
  assign n9432 = ~Pg35 & Ng2719;
  assign n9433 = Ng2841 & ~Ng2724;
  assign n9434 = n5327 & n9433;
  assign n9435 = ~n9432 & ~n9434;
  assign n9436 = Ng2724 & n7718;
  assign n9437 = ~n5327 & n9436;
  assign n3818_1 = ~n9435 | n9437;
  assign n9439 = Ng4704 & n6069;
  assign n9440 = ~Ng5357 & ~Ng5348;
  assign n9441 = Ng5357 & ~Ng5352;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = Ng5297 & n9442;
  assign n9444 = ~Ng5297 & ~n9442;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = Pg33959 & ~n9445;
  assign n9447 = ~Ng4704 & ~n9446;
  assign n9448 = Pg35 & n4616;
  assign n9449 = ~n9447 & n9448;
  assign n3823_1 = n9439 | n9449;
  assign n9451 = ~Ng2878 & n9377;
  assign n9452 = ~Pg35 & ~Ng2882;
  assign n3833_1 = ~n9451 & ~n9452;
  assign n9454 = Ng5176 & n5041;
  assign n9455 = n5018 & n9454;
  assign n9456 = ~Pg35 & ~Ng5264;
  assign n9457 = ~n9455 & ~n9456;
  assign n9458 = Pg35 & ~n9454;
  assign n9459 = ~Ng5220 & n9458;
  assign n3838_1 = n9457 & ~n9459;
  assign n9461 = ~Pg35 & Ng613;
  assign n9462 = Ng617 & n5737;
  assign n9463 = ~n5943 & ~n9462;
  assign n9464 = ~n5944 & ~n9463;
  assign n3843_1 = n9461 | n9464;
  assign n9466 = ~Pg35 & Ng324;
  assign n3852_1 = n8277 | n9466;
  assign n9468 = Ng1270 & n7939;
  assign n9469 = ~n4823 & n9468;
  assign n9470 = Pg35 & ~n9469;
  assign n3857 = Ng1274 & ~n9470;
  assign n9472 = ~Ng6513 & n7313;
  assign n9473 = ~Pg35 & Ng6509;
  assign n9474 = ~n9260 & ~n9473;
  assign n9475 = ~n7313 & n9474;
  assign n3862_1 = ~n9472 & ~n9475;
  assign n9477 = n8268 & n8275;
  assign n9478 = ~Pg35 & ~Ng311;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = Pg35 & n8276;
  assign n9481 = ~Ng336 & n9480;
  assign n3867_1 = n9479 & ~n9481;
  assign n9483 = Pg35 & ~Ng2882;
  assign n9484 = n9376 & n9483;
  assign n9485 = ~Pg35 & ~Ng2898;
  assign n3872_1 = ~n9484 & ~n9485;
  assign n9487 = Pg35 & n4825;
  assign n9488 = Pg35 & ~n6166_1;
  assign n9489 = Ng930 & ~n9488;
  assign n3877_1 = ~n9487 & n9489;
  assign n9491 = ~Pg35 & Ng1913;
  assign n9492 = Ng1906 & n5873;
  assign n9493 = n4951 & n5876;
  assign n9494 = ~n9492 & ~n9493;
  assign n3882_1 = n9491 | ~n9494;
  assign n3887_1 = Pg6745 & Pg35;
  assign n9497 = ~Ng2193 & n8039;
  assign n9498 = ~Pg35 & \[4428] ;
  assign n9499 = Ng2799 & n8036;
  assign n9500 = ~n9498 & ~n9499;
  assign n3897 = n9497 | ~n9500;
  assign n9502 = Pg35 & Ng4912;
  assign n9503 = ~Pg35 & Ng4907;
  assign n3908 = n9502 | n9503;
  assign n9505 = ~Pg35 & Ng4146;
  assign n3913 = n7055 | n9505;
  assign n9507 = ~Pg35 & Ng2537;
  assign n9508 = Pg35 & ~Ng2541;
  assign n9509 = ~n9507 & ~n9508;
  assign n9510 = n7009 & n9509;
  assign n9511 = ~Ng2541 & ~n7009;
  assign n3918_1 = ~n9510 & ~n9511;
  assign n9513 = Pg35 & n6498_1;
  assign n9514 = Ng2153 & n9513;
  assign n9515 = n4589 & n5089;
  assign n9516 = Pg35 & ~n9515;
  assign n9517 = ~Ng2227 & n9516;
  assign n9518 = ~n9514 & ~n9517;
  assign n9519 = ~Ng2197 & ~n6498_1;
  assign n9520 = ~Ng2153 & ~n9519;
  assign n3923_1 = ~n9518 & ~n9520;
  assign n9522 = ~Ng550 & \[4435] ;
  assign n9523 = Pg35 & n9522;
  assign n9524 = ~Pg35 & ~Ng534;
  assign n3928 = ~n9523 & ~n9524;
  assign n9526 = Ng255 & n7393;
  assign n9527 = Pg14201 & n7390;
  assign n9528 = ~Pg35 & Ng225;
  assign n9529 = ~n9527 & ~n9528;
  assign n3933_1 = n9526 | ~n9529;
  assign n9531 = Ng1874 & n5299;
  assign n9532 = Pg35 & n9531;
  assign n9533 = ~Pg35 & Ng1926;
  assign n9534 = Ng1945 & n5838;
  assign n9535 = Ng1890 & n4654;
  assign n9536 = Ng1926 & ~Ng1917;
  assign n9537 = Ng1878 & n9536;
  assign n9538 = Ng1870 & n9211;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = ~Ng1917 & Ng1894;
  assign n9541 = Ng1886 & n9540;
  assign n9542 = Ng1882 & ~Ng1926;
  assign n9543 = ~Ng1894 & n9542;
  assign n9544 = ~n9541 & ~n9543;
  assign n9545 = n9539 & n9544;
  assign n9546 = ~n9535 & n9545;
  assign n9547 = n5836 & ~n9546;
  assign n9548 = ~n9534 & ~n9547;
  assign n9549 = ~n9533 & n9548;
  assign n3938 = n9532 | ~n9549;
  assign n9551 = ~Ng5164 & Ng5170;
  assign n9552 = n5820 & n9551;
  assign n9553 = n5083 & n9552;
  assign n9554 = ~Pg35 & Ng5224;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = Pg35 & Ng5240;
  assign n9557 = ~n9552 & n9556;
  assign n3943_1 = ~n9555 | n9557;
  assign n9559 = ~Pg35 & Ng1437;
  assign n9560 = Ng1437 & n6270;
  assign n9561 = n7677 & n9560;
  assign n9562 = Ng1478 & n9561;
  assign n9563 = Pg35 & Ng1478;
  assign n9564 = ~n9561 & ~n9563;
  assign n9565 = ~n9562 & ~n9564;
  assign n3948_1 = n9559 | n9565;
  assign n9567 = ~Pg35 & Ng3857;
  assign n9568 = ~n6918 & ~n8079;
  assign n9569 = n8025 & ~n9568;
  assign n3953_1 = n9567 | n9569;
  assign n9571 = Ng1945 & ~n5838;
  assign n9572 = ~n5838 & ~n9212;
  assign n9573 = Ng1959 & ~n9572;
  assign n9574 = ~n9571 & n9573;
  assign n9575 = n9571 & ~n9573;
  assign n3958 = n9574 | n9575;
  assign n9577 = Ng3480 & n7361;
  assign n9578 = ~Ng3476 & n8600;
  assign n9579 = Ng3476 & ~n8600;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = ~n7361 & ~n9580;
  assign n3963_1 = n9577 | n9581;
  assign n9583 = n4713 & n7556;
  assign n9584 = n5083 & n9583;
  assign n9585 = ~Pg35 & Ng6637;
  assign n9586 = ~n9584 & ~n9585;
  assign n9587 = Pg35 & Ng6653;
  assign n9588 = ~n9583 & n9587;
  assign n3968 = ~n9586 | n9588;
  assign n9590 = Pg35 & ~Ng2864;
  assign n9591 = n5802_1 & n9590;
  assign n9592 = ~Pg35 & ~Ng2856;
  assign n3976_1 = ~n9591 & ~n9592;
  assign n9594 = Ng4894 & n9250;
  assign n9595 = ~Ng6741 & ~Ng6732;
  assign n9596 = ~Ng6736 & Ng6741;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = Ng6682 & n9597;
  assign n9599 = ~Ng6682 & ~n9597;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = n7836 & ~n9600;
  assign n9602 = ~Ng4894 & ~n9601;
  assign n9603 = Pg35 & n4610;
  assign n9604 = ~n9602 & n9603;
  assign n3981 = n9594 | n9604;
  assign n3989 = ~Ng3857 & n8026;
  assign n9607 = Ng513 & n5351;
  assign n9608 = Ng499 & ~n9607;
  assign n9609 = Ng518 & ~n5348;
  assign n9610 = n5351 & ~n9609;
  assign n9611 = ~n9608 & ~n9610;
  assign n3997_1 = Pg35 & ~n9611;
  assign n9613 = ~Ng1002 & n5606;
  assign n9614 = Pg35 & ~n9613;
  assign n9615 = ~n5618 & n9614;
  assign n9616 = ~Pg35 & Ng1008;
  assign n4002 = n9615 | n9616;
  assign n9618 = ~Pg35 & Ng772;
  assign n9619 = Ng776 & n5145;
  assign n9620 = ~n5138 & ~n9619;
  assign n9621 = ~n5139 & ~n9620;
  assign n4007 = n9618 | n9621;
  assign n4016 = n7422 & n7978;
  assign n9624 = Ng2453 & ~n6149;
  assign n9625 = Ng2476 & n6149;
  assign n9626 = ~n6153_1 & ~n9625;
  assign n4021_1 = n9624 | ~n9626;
  assign n9628 = Pg35 & n6249;
  assign n9629 = Ng1648 & n9628;
  assign n9630 = ~Pg35 & Ng1664;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = n5843 & n7365;
  assign n9633 = Ng1657 & n8570;
  assign n9634 = ~n9632 & ~n9633;
  assign n4026 = ~n9631 | ~n9634;
  assign n9636 = ~Pg35 & Ng2361;
  assign n9637 = ~Ng2375 & n4978;
  assign n9638 = ~Ng1589 & ~n4976;
  assign n9639 = ~n4984 & ~n9638;
  assign n9640 = Ng2375 & ~n4979_1;
  assign n9641 = n9639 & n9640;
  assign n9642 = ~n9639 & ~n9640;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = ~n4978 & n9643;
  assign n9645 = Pg35 & ~n9644;
  assign n9646 = ~n9637 & n9645;
  assign n4031_1 = n9636 | n9646;
  assign n9648 = Pg35 & ~Ng890;
  assign n9649 = Ng862 & ~n9648;
  assign n9650 = ~Ng862 & n9648;
  assign n4048_1 = n9649 | n9650;
  assign n9652 = ~Pg35 & Ng278;
  assign n4053 = n9429 | n9652;
  assign n9654 = ~Pg35 & Ng3155;
  assign n9655 = ~n5015 & ~n8807;
  assign n9656 = n5252 & ~n9655;
  assign n4058_1 = n9654 | n9656;
  assign n9658 = Ng2370 & ~n7142;
  assign n9659 = ~n7142 & ~n7599;
  assign n9660 = Ng2384 & ~n9659;
  assign n9661 = ~n9658 & n9660;
  assign n9662 = n9658 & ~n9660;
  assign n4063_1 = n9661 | n9662;
  assign n9664 = Ng4616 & n7476;
  assign n9665 = Pg35 & ~n8904;
  assign n9666 = Ng4608 & ~n9665;
  assign n4071_1 = n9664 | n9666;
  assign n9668 = ~Pg35 & Ng4558;
  assign n9669 = Pg6749 & Pg35;
  assign n4076_1 = n9668 | n9669;
  assign n9671 = ~Pg35 & ~Ng2012;
  assign n9672 = n4596 & ~n5660;
  assign n9673 = ~n6911 & n9672;
  assign n9674 = Ng2024 & ~n9672;
  assign n9675 = Pg35 & ~n9674;
  assign n9676 = ~n9673 & n9675;
  assign n4081 = ~n9671 & ~n9676;
  assign n9678 = Ng2795 & n8036;
  assign n9679 = ~Ng2036 & n8039;
  assign n9680 = ~Pg35 & Ng2791;
  assign n9681 = ~n9679 & ~n9680;
  assign n4090 = n9678 | ~n9681;
  assign n9683 = ~Pg35 & Ng608;
  assign n9684 = Ng613 & n5737;
  assign n9685 = ~n5757 & ~n9684;
  assign n9686 = ~n5943 & ~n9685;
  assign n4095_1 = n9683 | n9686;
  assign n9688 = Pg35 & ~Ng4521;
  assign n9689 = n5180 & n9688;
  assign n9690 = Ng4489 & Ng4483;
  assign n9691 = Ng4492 & Ng4486;
  assign n9692 = n9690 & n9691;
  assign n9693 = Ng4527 & ~n9692;
  assign n9694 = ~Ng4527 & n9692;
  assign n9695 = Pg35 & ~n9694;
  assign n9696 = ~n9693 & n9695;
  assign n9697 = Ng4521 & ~n9696;
  assign n4100_1 = n9689 | n9697;
  assign n9699 = Pg35 & ~Ng1834;
  assign n9700 = Ng1840 & n9699;
  assign n9701 = ~Ng1840 & ~n9699;
  assign n9702 = ~n9700 & ~n9701;
  assign n9703 = n8858 & n9702;
  assign n9704 = Ng1844 & ~n8858;
  assign n4105 = n9703 | n9704;
  assign n9706 = Ng5873 & ~Ng5881;
  assign n9707 = n6426 & n9706;
  assign n9708 = Pg35 & ~Ng5937;
  assign n9709 = ~n9707 & n9708;
  assign n9710 = n5018 & n9707;
  assign n9711 = ~Pg35 & ~Ng5921;
  assign n9712 = ~n9710 & ~n9711;
  assign n4110_1 = ~n9709 & n9712;
  assign n9714 = Ng4567 & ~n5406;
  assign n9715 = ~n6666_1 & ~n9714;
  assign n4115_1 = n7572 | ~n9715;
  assign n9717 = ~Ng2523 & ~n9340;
  assign n9718 = Pg35 & Ng2514;
  assign n9719 = Ng2518 & n9718;
  assign n9720 = ~Ng2518 & ~n9718;
  assign n9721 = ~n9719 & ~n9720;
  assign n9722 = n9340 & ~n9721;
  assign n4120_1 = ~n9717 & ~n9722;
  assign n9724 = ~Pg13895 & ~Pg16718;
  assign n9725 = ~n6651 & ~n9724;
  assign n9726 = Pg35 & ~Pg16603;
  assign n9727 = ~Pg14421 & ~Pg16624;
  assign n9728 = n9726 & n9727;
  assign n4125 = ~n9725 & n9728;
  assign n9730 = ~Pg35 & Ng2629;
  assign n9731 = ~Ng2643 & n5533;
  assign n9732 = ~Ng1589 & ~n5531;
  assign n9733 = ~n5541 & ~n9732;
  assign n9734 = Ng2643 & ~n8991;
  assign n9735 = n9733 & n9734;
  assign n9736 = ~n9733 & ~n9734;
  assign n9737 = ~n9735 & ~n9736;
  assign n9738 = ~n5533 & n9737;
  assign n9739 = Pg35 & ~n9738;
  assign n9740 = ~n9731 & n9739;
  assign n4129_1 = n9730 | n9740;
  assign n9742 = ~Ng1442 & n9310;
  assign n9743 = Ng1495 & n6265;
  assign n9744 = Pg35 & Ng1489;
  assign n9745 = ~n9743 & n9744;
  assign n4134_1 = n9742 | n9745;
  assign n9747 = Pg8291 & Ng218;
  assign n9748 = Ng191 & n9747;
  assign n9749 = ~Pg8358 & ~n9747;
  assign n9750 = ~n9748 & ~n9749;
  assign n9751 = Pg35 & n9750;
  assign n9752 = ~Pg35 & Ng222;
  assign n4139_1 = n9751 | n9752;
  assign n9754 = Ng2547 & n9508;
  assign n9755 = ~Ng2547 & ~n9508;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = ~n5010 & ~n9756;
  assign n9758 = ~Ng2551 & n5010;
  assign n4143 = ~n9757 & ~n9758;
  assign n9760 = Ng5156 & ~Pg32975;
  assign n9761 = n5018 & n9760;
  assign n9762 = n5083 & ~n9760;
  assign n4148 = n9761 | n9762;
  assign n9764 = Pg35 & Ng4281;
  assign n9765 = ~Pg35 & ~Ng4245;
  assign n4161 = ~n9764 & ~n9765;
  assign n9767 = Pg35 & ~n7948;
  assign n9768 = ~n5873 & ~n9767;
  assign n9769 = Ng1950 & n9768;
  assign n9770 = Ng1955 & ~n9768;
  assign n4165_1 = n9769 | n9770;
  assign n9772 = ~Pg35 & Ng6044;
  assign n9773 = n6791 & ~n7810;
  assign n9774 = ~Ng6049 & ~n9773;
  assign n9775 = ~n7807 & ~n9774;
  assign n4170_1 = n9772 | n9775;
  assign n9777 = ~Pg35 & Ng2269;
  assign n9778 = Pg35 & ~Ng2273;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = Pg35 & ~n7537;
  assign n9781 = ~n9513 & ~n9780;
  assign n9782 = n9779 & n9781;
  assign n9783 = ~Ng2273 & ~n9781;
  assign n4175 = ~n9782 & ~n9783;
  assign n9785 = ~Ng6395 & ~Ng6386;
  assign n9786 = Ng6395 & ~Ng6390;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = Ng6336 & n9787;
  assign n9789 = ~Ng6336 & ~n9787;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = n5385 & ~n9790;
  assign n9792 = ~Ng4771 & ~n9791;
  assign n9793 = Ng4771 & n5937;
  assign n9794 = n4615 & n4744;
  assign n9795 = Pg35 & n9794;
  assign n9796 = ~n9793 & ~n9795;
  assign n4183_1 = ~n9792 & ~n9796;
  assign n9798 = ~Ng6148 & Pg9682;
  assign n9799 = ~Ng6098 & ~n9798;
  assign n9800 = Pg35 & ~Pg9741;
  assign n9801 = ~n9799 & n9800;
  assign n9802 = ~Pg35 & Ng6148;
  assign n4188 = n9801 | n9802;
  assign n9804 = Ng3147 & ~n4731;
  assign n9805 = n5018 & n9804;
  assign n9806 = n5083 & ~n9804;
  assign n4193 = n9805 | n9806;
  assign n9808 = Pg35 & n6654;
  assign n4198_1 = Ng3343 & ~n9808;
  assign n9810 = Ng2265 & n6709;
  assign n9811 = ~Ng2265 & ~n6709;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = n9781 & n9812;
  assign n9814 = Ng2269 & ~n9781;
  assign n4203_1 = n9813 | n9814;
  assign n9816 = Pg35 & Ng26936;
  assign n9817 = ~Ng2712 & n9816;
  assign n9818 = ~Pg35 & Ng2841;
  assign n4212_1 = n9817 | n9818;
  assign n9820 = ~Pg35 & Ng622;
  assign n9821 = Ng626 & n5737;
  assign n9822 = ~n5945 & ~n9821;
  assign n9823 = ~n7345 & ~n9822;
  assign n4217_1 = n9820 | n9823;
  assign n9825 = ~Ng2729 & ~n7797;
  assign n9826 = ~n7798 & ~n9825;
  assign n9827 = n7718 & ~n9826;
  assign n9828 = ~Pg35 & ~Ng2724;
  assign n4222_1 = ~n9827 & ~n9828;
  assign n9830 = ~Pg35 & ~Ng5352;
  assign n9831 = Ng5357 & ~Pg33959;
  assign n9832 = ~Ng5357 & Pg33959;
  assign n9833 = ~n7916 & n9832;
  assign n9834 = Pg35 & ~n9833;
  assign n9835 = ~n9831 & n9834;
  assign n4227_1 = ~n9830 & ~n9835;
  assign n9837 = n6592 & n6594;
  assign n9838 = ~Ng4991 & n9837;
  assign n9839 = Ng4991 & n6596_1;
  assign n9840 = ~Pg35 & Ng4983;
  assign n9841 = ~n9839 & ~n9840;
  assign n4232 = n9838 | ~n9841;
  assign n9843 = Ng4709 & n5552;
  assign n9844 = Pg35 & n4744;
  assign n9845 = n4747 & n5550;
  assign n9846 = ~n9844 & ~n9845;
  assign n9847 = ~n5548 & ~n9846;
  assign n9848 = ~Pg35 & Ng4785;
  assign n9849 = ~n9847 & ~n9848;
  assign n4240 = n9843 | ~n9849;
  assign n9851 = ~Pg35 & ~Ng2917;
  assign n9852 = Pg44 & Pg35;
  assign n9853 = ~Ng2932 & ~Ng2927;
  assign n9854 = n9852 & n9853;
  assign n4245_1 = ~n9851 & ~n9854;
  assign n9856 = Ng4628 & n5559;
  assign n9857 = ~Ng4340 & ~n9856;
  assign n9858 = ~n5561 & ~n9857;
  assign n9859 = Pg35 & ~n9858;
  assign n9860 = ~n5309 & n9859;
  assign n9861 = ~Pg35 & ~Ng4643;
  assign n4250 = ~n9860 & ~n9861;
  assign n9863 = ~Pg35 & ~Ng5909;
  assign n9864 = n4717 & n7650;
  assign n9865 = n5018 & n9864;
  assign n9866 = Pg35 & ~Ng5929;
  assign n9867 = ~n9864 & n9866;
  assign n9868 = ~n9865 & ~n9867;
  assign n4255 = ~n9863 & n9868;
  assign n9870 = Pg35 & Ng4907;
  assign n9871 = ~Pg35 & Ng4922;
  assign n4260 = n9870 | n9871;
  assign n9873 = Ng4035 & n6698;
  assign n9874 = ~Pg35 & Ng3965;
  assign n9875 = ~n9873 & ~n9874;
  assign n4268_1 = n8406 | ~n9875;
  assign n9877 = Pg35 & Pg9019;
  assign n9878 = Ng4291 & ~n9877;
  assign n9879 = ~Ng4291 & n9877;
  assign n4273 = n9878 | n9879;
  assign n9881 = ~Pg35 & Ng914;
  assign n9882 = Ng918 & n6167;
  assign n9883 = ~n6164 & ~n9882;
  assign n9884 = ~n6165 & ~n9883;
  assign n4278 = n9881 | n9884;
  assign n9886 = ~Ng4082 & ~n6201;
  assign n9887 = ~n6202_1 & ~n9886;
  assign n9888 = n7718 & ~n9887;
  assign n9889 = ~Pg35 & ~Ng4141;
  assign n4283_1 = ~n9888 & ~n9889;
  assign n4288_1 = Pg35 & Ng6573;
  assign n9892 = ~Pg35 & Ng2016;
  assign n9893 = n4639 & n6947;
  assign n9894 = n8816 & n9893;
  assign n9895 = ~Ng2036 & ~n9893;
  assign n9896 = Pg35 & ~n9895;
  assign n9897 = ~n9894 & n9896;
  assign n4292_1 = n9892 | n9897;
  assign n9899 = ~Pg35 & Ng586;
  assign n9900 = Ng577 & n5737;
  assign n9901 = ~n5750 & ~n9900;
  assign n9902 = ~n5751 & ~n9901;
  assign n4297_1 = n9899 | n9902;
  assign n9904 = ~Pg35 & Ng1608;
  assign n9905 = Pg31862 & ~n5227;
  assign n9906 = Pg35 & ~n9905;
  assign n9907 = ~n5237 & ~n9906;
  assign n9908 = ~n9904 & n9907;
  assign n9909 = ~Ng1620 & n9906;
  assign n4302_1 = ~n9908 & ~n9909;
  assign n9911 = Ng2775 & n5961;
  assign n9912 = Ng2783 & n5001;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = Ng2771 & n5256;
  assign n9915 = Ng2787 & n5327;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = n9913 & n9916;
  assign n9918 = n5959 & ~n9917;
  assign n9919 = ~Ng1811 & n5961;
  assign n9920 = ~Ng1945 & n5001;
  assign n9921 = ~Ng1677 & n5256;
  assign n9922 = ~Ng2079 & n5327;
  assign n9923 = ~n9921 & ~n9922;
  assign n9924 = ~n9920 & n9923;
  assign n9925 = ~n9919 & n9924;
  assign n9926 = ~n5959 & ~n9925;
  assign n9927 = Pg35 & ~n9926;
  assign n9928 = ~n9918 & n9927;
  assign n9929 = ~Pg35 & Ng2771;
  assign n4307_1 = n9928 | n9929;
  assign n9931 = Ng667 & n7910;
  assign n9932 = Ng686 & ~n7910;
  assign n4312_1 = n9931 | n9932;
  assign n9934 = ~Ng930 & n6165;
  assign n9935 = Pg35 & ~n9934;
  assign n9936 = Ng925 & ~n9935;
  assign n9937 = ~n6166_1 & n6167;
  assign n9938 = Ng930 & n9937;
  assign n4317_1 = n9936 | n9938;
  assign n9940 = Ng3873 & ~Ng3881;
  assign n9941 = n6918 & n9940;
  assign n9942 = n5018 & n9941;
  assign n9943 = ~Pg35 & ~Ng3921;
  assign n9944 = ~n9942 & ~n9943;
  assign n9945 = Pg35 & ~n9941;
  assign n9946 = ~Ng3937 & n9945;
  assign n4322_1 = n9944 & ~n9946;
  assign n9948 = ~Pg35 & Ng812;
  assign n9949 = ~Ng817 & ~n5150;
  assign n9950 = n8249 & ~n9949;
  assign n4327_1 = n9948 | n9950;
  assign n4332_1 = ~Ng1249 & n5591;
  assign n9953 = Ng832 & Ng827;
  assign n9954 = Pg35 & ~n7042;
  assign n9955 = ~n9953 & n9954;
  assign n9956 = ~n5151 & ~n9955;
  assign n9957 = Ng837 & ~n9956;
  assign n9958 = Pg35 & ~n7043;
  assign n9959 = Ng703 & ~n9958;
  assign n9960 = ~n5151 & n9959;
  assign n4337_1 = n9957 | n9960;
  assign n9962 = ~Pg35 & Ng595;
  assign n9963 = Ng599 & n5737;
  assign n9964 = ~n5754 & ~n9963;
  assign n9965 = ~n5755 & ~n9964;
  assign n4345_1 = n9962 | n9965;
  assign n9967 = ~Ng5475 & n7205;
  assign n9968 = Pg35 & ~Ng5475;
  assign n9969 = ~Pg35 & Ng5471;
  assign n9970 = ~n9968 & ~n9969;
  assign n9971 = ~n7205 & n9970;
  assign n4350_1 = ~n9967 & ~n9971;
  assign n9973 = ~Pg35 & Ng736;
  assign n9974 = ~Ng739 & ~n5130;
  assign n9975 = ~n5131 & n5145;
  assign n9976 = ~n9974 & n9975;
  assign n4355_1 = n9973 | n9976;
  assign n9978 = ~Pg35 & ~Ng5933;
  assign n9979 = n6427 & n7328;
  assign n9980 = Pg35 & ~Ng5949;
  assign n9981 = ~n9979 & n9980;
  assign n9982 = n5018 & n9979;
  assign n9983 = ~n9981 & ~n9982;
  assign n4360_1 = ~n9978 & n9983;
  assign n9985 = n4537 & n7836;
  assign n9986 = n7083 & n9985;
  assign n9987 = Ng6682 & ~n7836;
  assign n9988 = ~n4538 & n7836;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = ~n9986 & ~n9989;
  assign n9991 = Pg35 & ~n9990;
  assign n9992 = Pg35 & Ng6682;
  assign n9993 = ~Ng6741 & ~n9992;
  assign n4365_1 = ~n9991 & ~n9993;
  assign n4370 = ~Ng904 & n6167;
  assign n9996 = Pg35 & Ng2873;
  assign n9997 = ~Pg35 & Ng2868;
  assign n4375 = n9996 | n9997;
  assign n9999 = Ng1760 & n6185;
  assign n10000 = Ng1792 & n9999;
  assign n10001 = Pg35 & ~n10000;
  assign n10002 = Ng1854 & n10001;
  assign n10003 = Ng1848 & ~n10001;
  assign n4380_1 = n10002 | n10003;
  assign n10005 = Pg35 & n9327;
  assign n10006 = Ng5080 & ~n10005;
  assign n10007 = ~Ng5084 & ~n9324;
  assign n10008 = ~n9326 & ~n10007;
  assign n10009 = Pg35 & ~Ng5080;
  assign n10010 = ~n10008 & n10009;
  assign n4385_1 = n10006 | n10010;
  assign n10012 = n5318 & n5374;
  assign n10013 = n5083 & n10012;
  assign n10014 = ~Pg35 & Ng5587;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = Pg35 & Ng5603;
  assign n10017 = ~n10012 & n10016;
  assign n4390 = ~n10015 | n10017;
  assign n10019 = Ng2495 & n6965;
  assign n10020 = Pg35 & n6961;
  assign n10021 = Ng2465 & ~n10020;
  assign n10022 = ~n6965 & n10021;
  assign n4398_1 = n10019 | n10022;
  assign n10024 = Ng2465 & ~n6959;
  assign n10025 = ~Ng2495 & n10024;
  assign n10026 = n7004 & n10025;
  assign n10027 = ~Pg35 & Ng2429;
  assign n10028 = Pg35 & Ng2437;
  assign n10029 = ~n10025 & n10028;
  assign n10030 = ~n10027 & ~n10029;
  assign n4403_1 = n10026 | ~n10030;
  assign n10032 = ~Ng2102 & n6950;
  assign n10033 = ~Pg35 & Ng2098;
  assign n10034 = ~n7292 & ~n10033;
  assign n10035 = ~n6950 & n10034;
  assign n4408 = ~n10032 & ~n10035;
  assign n10037 = Ng2185 & ~n5259;
  assign n10038 = Ng2208 & n5259;
  assign n10039 = n5843 & n7984;
  assign n10040 = ~n10038 & ~n10039;
  assign n4413 = n10037 | ~n10040;
  assign n10042 = ~Pg35 & ~Ng2583;
  assign n10043 = ~n5533 & n8113;
  assign n10044 = ~n5542_1 & n10043;
  assign n10045 = Ng2579 & ~n10043;
  assign n10046 = Pg35 & ~n10045;
  assign n10047 = ~n10044 & n10046;
  assign n4418_1 = ~n10042 & ~n10047;
  assign n10049 = ~Pg35 & ~Ng4072;
  assign n10050 = Ng4064 & n7718;
  assign n4423 = ~n10049 & ~n10050;
  assign n10052 = Ng4899 & n6595;
  assign n10053 = n4688_1 & n6593;
  assign n10054 = Pg35 & n4686;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = ~n5817 & ~n10055;
  assign n10057 = ~Pg35 & Ng4975;
  assign n10058 = ~n10056 & ~n10057;
  assign n4428_1 = n10052 | ~n10058;
  assign n10060 = ~Pg35 & ~Ng2715;
  assign n10061 = ~n5256 & ~n5327;
  assign n10062 = n7718 & ~n10061;
  assign n4433_1 = ~n10060 & ~n10062;
  assign n10064 = Ng4785 & n5552;
  assign n10065 = ~Pg35 & Ng4776;
  assign n10066 = ~n5548 & n5550;
  assign n10067 = ~Ng4785 & n10066;
  assign n10068 = ~n10065 & ~n10067;
  assign n4438 = n10064 | ~n10068;
  assign n10070 = ~Pg35 & ~Ng5563;
  assign n10071 = n4726 & n7624;
  assign n10072 = ~n5018 & n10071;
  assign n10073 = Pg35 & ~Ng5583;
  assign n10074 = ~n10071 & ~n10073;
  assign n10075 = ~n10072 & ~n10074;
  assign n4443_1 = ~n10070 & ~n10075;
  assign n10077 = ~Pg35 & Ng776;
  assign n10078 = Ng781 & n5145;
  assign n10079 = ~n5139 & ~n10078;
  assign n10080 = ~n5140 & ~n10079;
  assign n4448 = n10077 | n10080;
  assign n10082 = Ng6173 & n5387;
  assign n10083 = Ng6167 & ~n5387;
  assign n4453 = n10082 | n10083;
  assign n10085 = ~Pg35 & ~Ng2902;
  assign n10086 = ~Ng2917 & n4823;
  assign n10087 = n9487 & n10086;
  assign n4461 = ~n10085 & ~n10087;
  assign n10089 = ~Pg35 & Ng691;
  assign n10090 = ~Ng686 & ~n5351;
  assign n10091 = ~Ng691 & n5351;
  assign n10092 = Ng703 & n5894;
  assign n10093 = n10091 & n10092;
  assign n10094 = Pg35 & ~n10093;
  assign n10095 = ~n10090 & n10094;
  assign n4466 = n10089 | n10095;
  assign n10097 = ~Pg35 & Ng1280;
  assign n10098 = Ng1252 & n5591;
  assign n10099 = ~n7817 & ~n10098;
  assign n10100 = ~n7818 & ~n10099;
  assign n4471 = n10097 | n10100;
  assign n10102 = ~Pg35 & Ng667;
  assign n10103 = ~Ng671 & ~n5884;
  assign n10104 = n5900 & ~n10103;
  assign n4476 = n10102 | n10104;
  assign n10106 = Ng2259 & n9781;
  assign n10107 = Ng2265 & ~n9781;
  assign n4481 = n10106 | n10107;
  assign n10109 = n5497 & n6385;
  assign n10110 = n5083 & n10109;
  assign n10111 = ~Pg35 & Ng6267;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = Pg35 & Ng6283;
  assign n10114 = ~n10109 & n10113;
  assign n4486_1 = ~n10112 | n10114;
  assign n10116 = ~Ng5527 & ~n6773;
  assign n10117 = Pg35 & ~n10116;
  assign n10118 = Ng5523 & ~n10117;
  assign n10119 = Ng5527 & n6775;
  assign n4500 = n10118 | n10119;
  assign n10121 = ~Pg35 & Ng4486;
  assign n4505 = n9669 | n10121;
  assign n10123 = Ng1968 & n9768;
  assign n10124 = Ng1974 & ~n9768;
  assign n4510_1 = n10123 | n10124;
  assign n10126 = ~Pg35 & Ng1263;
  assign n10127 = Ng1270 & n5591;
  assign n10128 = ~n7939 & ~n10127;
  assign n10129 = ~n9468 & ~n10128;
  assign n4515_1 = n10126 | n10129;
  assign n10131 = Ng4966 & n6595;
  assign n10132 = Pg35 & ~n9837;
  assign n10133 = Ng4991 & ~n10132;
  assign n4520 = n10131 | n10133;
  assign n10135 = ~Pg35 & Ng6219;
  assign n6227 = Pg35 & Ng6227;
  assign n10137 = ~n7231 & n6227;
  assign n10138 = ~n7232 & ~n10137;
  assign n10139 = ~n5106 & ~n10138;
  assign n4525 = n10135 | n10139;
  assign n10141 = ~Pg35 & ~Ng3909;
  assign n10142 = n4733 & n8079;
  assign n10143 = n5018 & n10142;
  assign n10144 = Pg35 & ~Ng3929;
  assign n10145 = ~n10142 & n10144;
  assign n10146 = ~n10143 & ~n10145;
  assign n4530_1 = ~n10141 & n10146;
  assign n10148 = Ng5503 & ~n4727;
  assign n10149 = n5018 & n10148;
  assign n10150 = n5083 & ~n10148;
  assign n4535_1 = n10149 | n10150;
  assign n10152 = Ng4235 & Pg8870;
  assign n10153 = ~Pg8918 & ~Pg8916;
  assign n10154 = ~Pg11770 & ~Pg8920;
  assign n10155 = ~Pg8919 & ~Pg8917;
  assign n10156 = ~Pg8915 & n10155;
  assign n10157 = n10154 & n10156;
  assign n10158 = n10153 & n10157;
  assign n10159 = ~Ng4235 & ~Pg8870;
  assign n10160 = ~n10158 & n10159;
  assign n10161 = ~n10152 & ~n10160;
  assign n10162 = n7612 & n10161;
  assign n10163 = ~Pg35 & ~Ng4235;
  assign n10164 = Pg35 & ~n7611;
  assign n10165 = ~n10161 & n10164;
  assign n10166 = ~n10163 & ~n10165;
  assign n4540_1 = ~n10162 & n10166;
  assign n10168 = n6754 & n7650;
  assign n10169 = Pg35 & ~n10168;
  assign n10170 = Ng5925 & n10169;
  assign n10171 = ~Pg35 & Ng5901;
  assign n10172 = ~n5083 & ~n10171;
  assign n10173 = ~n10169 & ~n10172;
  assign n4545 = n10170 | n10173;
  assign n10175 = Pg13259 & n7745;
  assign n10176 = ~Ng976 & n4825;
  assign n10177 = ~Ng1129 & n10176;
  assign n10178 = Ng1129 & ~n10176;
  assign n10179 = ~n10177 & ~n10178;
  assign n10180 = n10175 & n10179;
  assign n10181 = ~Ng1099 & ~Ng1146;
  assign n10182 = n10175 & n10181;
  assign n10183 = ~Ng1124 & ~n10182;
  assign n10184 = Pg35 & ~n10183;
  assign n10185 = ~n10180 & n10184;
  assign n10186 = ~Pg35 & Ng1105;
  assign n4550_1 = n10185 | n10186;
  assign n10188 = ~Ng4955 & ~n6700;
  assign n10189 = ~n5669 & ~n10188;
  assign n10190 = n5677 & ~n10189;
  assign n10191 = ~n5670 & n6700;
  assign n10192 = Pg35 & ~n10191;
  assign n10193 = ~Ng4961 & ~n10192;
  assign n4555 = ~n10190 & ~n10193;
  assign n10195 = n5042_1 & n5820;
  assign n10196 = n5083 & n10195;
  assign n10197 = ~Pg35 & Ng5196;
  assign n10198 = ~n10196 & ~n10197;
  assign n10199 = Pg35 & Ng5224;
  assign n10200 = ~n10195 & n10199;
  assign n4560 = ~n10198 | n10200;
  assign n10202 = ~Pg35 & Ng2004;
  assign n10203 = Ng2040 & ~n5660;
  assign n10204 = ~Ng2070 & n10203;
  assign n10205 = n6912 & n10204;
  assign n10206 = Pg35 & Ng2012;
  assign n10207 = ~n10204 & n10206;
  assign n10208 = ~n10205 & ~n10207;
  assign n4565 = n10202 | ~n10208;
  assign n4570_1 = ~Ng6203 & n5111;
  assign n10211 = Pg35 & ~Pg32975;
  assign n10212 = Ng5120 & n10211;
  assign n10213 = Ng5156 & ~n10211;
  assign n4575 = n10212 | n10213;
  assign n10215 = ~Ng2389 & ~n9659;
  assign n10216 = Pg35 & Ng2380;
  assign n10217 = Ng2384 & n10216;
  assign n10218 = ~Ng2384 & ~n10216;
  assign n10219 = ~n10217 & ~n10218;
  assign n10220 = n9659 & ~n10219;
  assign n4583 = ~n10215 & ~n10220;
  assign n10222 = ~Ng2465 & ~n6959;
  assign n10223 = Ng2421 & n10222;
  assign n10224 = Pg35 & ~n10223;
  assign n10225 = Ng2429 & n10224;
  assign n10226 = ~Pg35 & Ng2433;
  assign n10227 = ~n7004 & ~n10226;
  assign n10228 = ~n10224 & ~n10227;
  assign n4593_1 = n10225 | n10228;
  assign n10230 = ~Pg35 & Ng2795;
  assign n10231 = Pg35 & ~Ng2795;
  assign n10232 = ~n5842 & ~n10231;
  assign n10233 = ~n4932 & n6718;
  assign n10234 = ~n10232 & n10233;
  assign n10235 = Pg35 & Ng2787;
  assign n10236 = ~n6718 & n10235;
  assign n10237 = ~n10234 & ~n10236;
  assign n4598 = n10230 | ~n10237;
  assign n10239 = Pg35 & ~Ng1287;
  assign n10240 = n4823 & n10239;
  assign n10241 = ~Pg35 & ~Ng1283;
  assign n4603 = ~n10240 & ~n10241;
  assign n10243 = ~Pg35 & Ng2671;
  assign n10244 = Pg35 & ~Ng2675;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = n8993 & n10245;
  assign n10247 = ~Ng2675 & ~n8993;
  assign n4608 = ~n10246 & ~n10247;
  assign n10249 = ~Pg35 & Ng4358;
  assign n10250 = ~Ng4593 & ~Ng4601;
  assign n10251 = Ng4633 & ~Ng4616;
  assign n10252 = ~Ng4584 & n10251;
  assign n10253 = n5560 & n10252;
  assign n10254 = ~Ng4608 & n10253;
  assign n10255 = n10250 & n10254;
  assign n10256 = n8676 & n10255;
  assign n4613 = n10249 | n10256;
  assign n10258 = ~n4606 & ~n5817;
  assign n10259 = Pg35 & n10258;
  assign n4618 = n6625_1 & n10259;
  assign n10261 = ~Ng1199 & ~n7030;
  assign n10262 = ~n7031 & ~n10261;
  assign n10263 = Pg35 & ~n10262;
  assign n10264 = ~Pg35 & ~Ng1193;
  assign n10265 = ~n10263 & ~n10264;
  assign n4623 = ~n6578 & n10265;
  assign n10267 = Ng1333 & ~n5516;
  assign n10268 = ~Ng1333 & n5516;
  assign n4628 = n10267 | n10268;
  assign n10270 = ~Pg35 & ~Ng5551;
  assign n10271 = n5317 & n6174;
  assign n10272 = Pg35 & ~Ng5547;
  assign n10273 = ~n10271 & n10272;
  assign n10274 = n5018 & n10271;
  assign n10275 = ~n10273 & ~n10274;
  assign n4632_1 = ~n10270 & n10275;
  assign n10277 = Pg35 & Ng2138;
  assign n10278 = ~Pg35 & Ng2130;
  assign n4637_1 = n10277 | n10278;
  assign n10280 = ~Pg35 & Ng2287;
  assign n10281 = n4586 & n4971;
  assign n10282 = Ng112 & n4587;
  assign n10283 = ~Ng112 & ~n4587;
  assign n10284 = ~n10282 & ~n10283;
  assign n10285 = n10281 & n10284;
  assign n10286 = n5842 & n10285;
  assign n10287 = ~n10280 & ~n10286;
  assign n10288 = n4928 & n10281;
  assign n10289 = Ng2338 & ~n10288;
  assign n10290 = Pg35 & n10289;
  assign n4645 = ~n10287 | n10290;
  assign n10292 = n5498 & n6227_1;
  assign n10293 = Pg35 & ~n10292;
  assign n10294 = ~Pg35 & ~Ng6251;
  assign n10295 = ~n5018 & ~n10294;
  assign n10296 = ~n10293 & ~n10295;
  assign n10297 = ~Ng6247 & n10293;
  assign n4653_1 = ~n10296 & ~n10297;
  assign n10299 = ~Ng1902 & n8039;
  assign n10300 = ~Pg35 & Ng2779;
  assign n10301 = ~n8036 & ~n10300;
  assign n10302 = ~n7279 & ~n10301;
  assign n4658 = n10299 | n10302;
  assign n10304 = n6919 & n7736;
  assign n10305 = Pg35 & ~n10304;
  assign n10306 = ~Pg35 & ~Ng3933;
  assign n10307 = ~n5018 & ~n10306;
  assign n10308 = ~n10305 & ~n10307;
  assign n10309 = ~Ng3949 & n10305;
  assign n4663_1 = ~n10308 & ~n10309;
  assign n4668 = Pg35 & Ng1291;
  assign n10312 = n4717 & n6426;
  assign n10313 = Pg35 & ~n10312;
  assign n10314 = ~Pg35 & ~Ng5929;
  assign n10315 = ~n5018 & ~n10314;
  assign n10316 = ~n10313 & ~n10315;
  assign n10317 = ~Ng5945 & n10313;
  assign n4673_1 = ~n10316 & ~n10317;
  assign n10319 = Ng5180 & ~Ng5188;
  assign n10320 = n9551 & n10319;
  assign n10321 = n5018 & n10320;
  assign n10322 = Pg35 & ~Ng5244;
  assign n10323 = ~n10320 & n10322;
  assign n10324 = ~Pg35 & ~Ng5228;
  assign n10325 = ~n10323 & ~n10324;
  assign n4678 = ~n10321 & n10325;
  assign n10327 = ~Ng2759 & ~n7799;
  assign n10328 = ~n7926 & ~n10327;
  assign n10329 = ~Pg35 & Ng2756;
  assign n10330 = ~n6197_1 & ~n10329;
  assign n4683 = n10328 | ~n10330;
  assign n10332 = Pg35 & n7836;
  assign n10333 = ~n9986 & n10332;
  assign n10334 = ~Ng6741 & n10333;
  assign n10335 = Ng6741 & n9250;
  assign n10336 = ~Pg35 & Ng6736;
  assign n10337 = ~n10335 & ~n10336;
  assign n4688 = n10334 | ~n10337;
  assign n10339 = ~Pg35 & Ng781;
  assign n10340 = Ng785 & n5145;
  assign n10341 = ~n5140 & ~n10340;
  assign n10342 = ~n5141 & ~n10341;
  assign n4693 = n10339 | n10342;
  assign n10344 = ~Pg35 & Ng1256;
  assign n10345 = Ng1259 & n5591;
  assign n10346 = ~n7819 & ~n10345;
  assign n10347 = ~n7938 & ~n10346;
  assign n4698 = n10344 | n10347;
  assign n10349 = ~Pg35 & Ng3480;
  assign n10350 = ~Ng3484 & ~n5487;
  assign n10351 = ~n6767 & ~n7361;
  assign n10352 = ~n10350 & ~n10351;
  assign n4703_1 = n10349 | n10352;
  assign n10354 = ~Pg8358 & n9747;
  assign n10355 = Pg35 & ~n10354;
  assign n10356 = ~Ng209 & ~n9747;
  assign n10357 = ~n9748 & ~n10356;
  assign n10358 = n10355 & ~n10357;
  assign n10359 = ~Ng191 & ~n10355;
  assign n4708 = ~n10358 & ~n10359;
  assign n10361 = n7753 & n8582;
  assign n10362 = n5018 & n10361;
  assign n10363 = ~Pg35 & ~Ng6581;
  assign n10364 = ~n10362 & ~n10363;
  assign n10365 = Pg35 & ~n10361;
  assign n10366 = ~Ng6609 & n10365;
  assign n4713_1 = n10364 & ~n10366;
  assign n10368 = ~Pg35 & Ng5511;
  assign n10369 = ~n5373 & ~n7624;
  assign n10370 = n6774 & ~n10369;
  assign n4718 = n10368 | n10370;
  assign n10372 = n4571 & ~n6959;
  assign n10373 = n7004 & n10372;
  assign n10374 = ~Pg35 & Ng2437;
  assign n10375 = Pg35 & Ng2449;
  assign n10376 = ~n10372 & n10375;
  assign n10377 = ~n10374 & ~n10376;
  assign n4723_1 = n10373 | ~n10377;
  assign n10379 = Ng2629 & n7670;
  assign n10380 = Pg35 & ~n10379;
  assign n10381 = Ng2575 & n10380;
  assign n10382 = ~Pg35 & Ng2579;
  assign n10383 = ~n5543 & ~n10382;
  assign n10384 = ~n10380 & ~n10383;
  assign n4728 = n10381 | n10384;
  assign n10386 = ~Pg35 & ~Ng2712;
  assign n10387 = Ng2715 & n7718;
  assign n4737_1 = ~n10386 & ~n10387;
  assign n10389 = ~Pg35 & Ng921;
  assign n10390 = Ng936 & n6167;
  assign n10391 = ~n6160 & ~n10390;
  assign n10392 = ~n6161_1 & ~n10391;
  assign n4742_1 = n10389 | n10392;
  assign n10394 = ~Pg35 & ~Ng2093;
  assign n10395 = ~Ng2028 & Ng2051;
  assign n10396 = n6947 & n10395;
  assign n10397 = Ng2098 & ~n10396;
  assign n10398 = Ng2089 & Ng2093;
  assign n10399 = ~Ng2089 & ~Ng2093;
  assign n10400 = ~n10398 & ~n10399;
  assign n10401 = n10396 & n10400;
  assign n10402 = Pg35 & ~n10401;
  assign n10403 = ~n10397 & n10402;
  assign n4747_1 = ~n10394 & ~n10403;
  assign n10405 = Pg35 & n7865;
  assign n10406 = Ng4643 & Ng4462;
  assign n10407 = Pg35 & n10406;
  assign n10408 = Ng4473 & ~n10407;
  assign n10409 = ~n8411 & ~n10408;
  assign n4752_1 = n10405 | ~n10409;
  assign n10411 = ~Pg35 & Ng599;
  assign n10412 = Ng604 & n5737;
  assign n10413 = ~n5755 & ~n10412;
  assign n10414 = ~n5756 & ~n10413;
  assign n4757_1 = n10411 | n10414;
  assign n10416 = Ng6561 & n7753;
  assign n10417 = n5083 & n10416;
  assign n10418 = ~Pg35 & Ng6641;
  assign n10419 = ~n10417 & ~n10418;
  assign n10420 = Pg35 & Ng6589;
  assign n10421 = ~n10416 & n10420;
  assign n4762 = ~n10419 | n10421;
  assign n10423 = ~Pg35 & ~Ng1890;
  assign n10424 = ~Ng1862 & Ng1906;
  assign n10425 = ~n4950 & n10424;
  assign n10426 = ~n4959 & n10425;
  assign n10427 = Ng1886 & ~n10425;
  assign n10428 = Pg35 & ~n10427;
  assign n10429 = ~n10426 & n10428;
  assign n4767_1 = ~n10423 & ~n10429;
  assign n10431 = Ng429 & n5151;
  assign n10432 = Ng433 & ~n5151;
  assign n4778_1 = n10431 | n10432;
  assign n10434 = ~Ng1906 & n4951;
  assign n10435 = Pg35 & ~n10434;
  assign n10436 = Ng1870 & n10435;
  assign n10437 = ~Pg35 & Ng1874;
  assign n10438 = ~n4960 & ~n10437;
  assign n10439 = ~n10435 & ~n10438;
  assign n4783_1 = n10436 | n10439;
  assign n10441 = Pg35 & Ng4249;
  assign n10442 = ~Pg35 & Ng4253;
  assign n4788 = n10441 | n10442;
  assign n10444 = Ng1811 & ~n8434;
  assign n10445 = ~n8429 & ~n8434;
  assign n10446 = Ng1825 & ~n10445;
  assign n10447 = ~n10444 & n10446;
  assign n10448 = n10444 & ~n10446;
  assign n4793_1 = n10447 | n10448;
  assign n10450 = Ng969 & ~n7063;
  assign n10451 = ~n5612 & ~n7065;
  assign n10452 = ~n5606 & ~n10451;
  assign n10453 = Pg35 & Ng1008;
  assign n10454 = ~n10452 & n10453;
  assign n4798 = n10450 | n10454;
  assign n10456 = Ng4392 & n6861;
  assign n10457 = ~n6866 & ~n10456;
  assign n10458 = ~Pg35 & Ng4417;
  assign n4803 = ~n10457 | n10458;
  assign n10460 = Ng3518 & n5635;
  assign n10461 = Pg35 & ~n10460;
  assign n10462 = Ng3546 & n10461;
  assign n10463 = ~Pg35 & Ng3598;
  assign n10464 = ~n5083 & ~n10463;
  assign n10465 = ~n10461 & ~n10464;
  assign n4808_1 = n10462 | n10465;
  assign n10467 = n4708_1 & n5042_1;
  assign n10468 = n5083 & n10467;
  assign n10469 = ~Pg35 & Ng5216;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = Pg35 & Ng5236;
  assign n10472 = ~n10467 & n10471;
  assign n4813_1 = ~n10470 | n10472;
  assign n10474 = Pg35 & ~n4659;
  assign n10475 = ~n8434 & ~n10474;
  assign n10476 = Ng1768 & ~n10475;
  assign n10477 = Pg35 & ~n6364;
  assign n10478 = ~Pg35 & Ng1748;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = n10475 & ~n10479;
  assign n4818_1 = n10476 | n10480;
  assign n10482 = ~Pg35 & Ng4849;
  assign n10483 = Ng4849 & n4604;
  assign n10484 = Ng4854 & n10483;
  assign n10485 = ~Ng4854 & ~n10483;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = n10259 & n10486;
  assign n4823_1 = n10482 | n10487;
  assign n10489 = n7216 & n8079;
  assign n10490 = n5018 & n10489;
  assign n10491 = ~Pg35 & ~Ng3901;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = Pg35 & ~n10489;
  assign n10494 = ~Ng3925 & n10493;
  assign n4828 = n10492 & ~n10494;
  assign n10496 = ~Ng6509 & n7840;
  assign n10497 = Pg35 & Ng6505;
  assign n10498 = ~Ng6500 & n10497;
  assign n10499 = Ng6500 & ~n10497;
  assign n10500 = ~n10498 & ~n10499;
  assign n10501 = ~n7840 & n10500;
  assign n4833_1 = ~n10496 & ~n10501;
  assign n10503 = Ng732 & ~n5120;
  assign n10504 = ~n5694 & ~n5702;
  assign n10505 = ~n5692 & ~n5701;
  assign n10506 = n10504 & ~n10505;
  assign n10507 = ~n10504 & n10505;
  assign n10508 = ~n10506 & ~n10507;
  assign n10509 = ~n5695 & ~n5700;
  assign n10510 = Ng255 & ~n10509;
  assign n10511 = ~Ng255 & n10509;
  assign n10512 = ~n10510 & ~n10511;
  assign n10513 = ~n10508 & ~n10512;
  assign n10514 = n10508 & n10512;
  assign n10515 = ~n10513 & ~n10514;
  assign n10516 = ~n10503 & ~n10515;
  assign n10517 = n10503 & n10515;
  assign n10518 = Pg35 & ~n10517;
  assign n4838_1 = ~n10516 & n10518;
  assign n10520 = ~Ng2476 & Ng2453;
  assign n10521 = Ng2445 & n10520;
  assign n10522 = Ng2485 & ~Ng2476;
  assign n10523 = Ng2437 & n10522;
  assign n10524 = ~Ng2485 & Ng2441;
  assign n10525 = ~Ng2453 & n10524;
  assign n10526 = ~n10523 & ~n10525;
  assign n10527 = Ng2449 & n4649_1;
  assign n10528 = Ng2429 & n9338;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = n10526 & n10529;
  assign n10531 = ~n10521 & n10530;
  assign n10532 = n6154 & ~n10531;
  assign n10533 = Ng2504 & n6149;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = Pg35 & Ng2453;
  assign n10536 = Ng2433 & n10535;
  assign n10537 = n5008_1 & n10536;
  assign n10538 = ~Pg35 & Ng2485;
  assign n10539 = ~n10537 & ~n10538;
  assign n4843 = ~n10534 | ~n10539;
  assign n10541 = Ng2185 & n5259;
  assign n10542 = n7159 & n8499;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = ~Pg35 & Ng2193;
  assign n10545 = ~n10039 & ~n10544;
  assign n4860_1 = ~n10543 | ~n10545;
  assign n10547 = Pg35 & Ng37;
  assign n10548 = ~Pg35 & Ng2894;
  assign n4865 = n10547 | n10548;
  assign n10550 = Pg35 & n8945;
  assign n10551 = Ng2040 & ~n5661;
  assign n10552 = ~n10550 & n10551;
  assign n10553 = Ng2070 & n5661;
  assign n4874 = n10552 | n10553;
  assign n10555 = ~Ng4176 & n6209;
  assign n10556 = ~Pg35 & ~Ng4172;
  assign n4883_1 = ~n10555 & ~n10556;
  assign n10558 = ~Pg16775 & ~Pg13966;
  assign n10559 = ~n4993_1 & ~n10558;
  assign n10560 = Pg35 & ~Pg14518;
  assign n10561 = ~Pg16659 & ~Pg16693;
  assign n10562 = n10560 & n10561;
  assign n4888_1 = ~n10559 & n10562;
  assign n10564 = ~Ng6181 & n5387;
  assign n10565 = ~Pg35 & Ng6177;
  assign n10566 = ~n7091 & ~n10565;
  assign n10567 = ~n5387 & n10566;
  assign n4900_1 = ~n10564 & ~n10567;
  assign n10569 = ~Pg35 & Ng6377;
  assign n10570 = ~Ng6381 & ~n6875;
  assign n10571 = n6877 & ~n10570;
  assign n4905 = n10569 | n10571;
  assign n10573 = ~Ng4765 & ~n9794;
  assign n10574 = ~n5669 & ~n10573;
  assign n10575 = n6519 & ~n10574;
  assign n10576 = ~n6513_1 & n9794;
  assign n10577 = Pg35 & ~n10576;
  assign n10578 = ~Ng4771 & ~n10577;
  assign n4910_1 = ~n10575 & ~n10578;
  assign n10580 = n4726 & n6174;
  assign n10581 = Pg35 & ~n10580;
  assign n10582 = ~Pg35 & ~Ng5567;
  assign n10583 = ~n5018 & ~n10582;
  assign n10584 = ~n10581 & ~n10583;
  assign n10585 = ~Ng5563 & n10581;
  assign n4915_1 = ~n10584 & ~n10585;
  assign n10587 = ~Ng1395 & ~n9409;
  assign n10588 = ~n9410 & ~n10587;
  assign n4920 = n9408 & n10588;
  assign n10590 = ~Pg35 & Ng1862;
  assign n10591 = ~Ng112 & ~n4580;
  assign n10592 = Ng112 & n4580;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = n4579_1 & n4942;
  assign n10595 = n10593 & n10594;
  assign n10596 = n5842 & n10595;
  assign n10597 = ~n10590 & ~n10596;
  assign n10598 = n4928 & n10594;
  assign n10599 = Ng1913 & ~n10598;
  assign n10600 = Pg35 & n10599;
  assign n4925 = ~n10597 | n10600;
  assign n10602 = n6532_1 & n7965;
  assign n10603 = ~Pg35 & Ng2338;
  assign n10604 = Ng2331 & n6528;
  assign n10605 = ~n10603 & ~n10604;
  assign n4930_1 = n10602 | ~n10605;
  assign n10607 = n6386 & n7336;
  assign n10608 = n5018 & n10607;
  assign n10609 = ~Pg35 & ~Ng6235;
  assign n10610 = ~n10608 & ~n10609;
  assign n10611 = Pg35 & ~n10607;
  assign n10612 = ~Ng6263 & n10611;
  assign n4935_1 = n10610 & ~n10612;
  assign n10614 = n4733 & n6918;
  assign n10615 = Pg35 & ~n10614;
  assign n10616 = Ng3945 & n10615;
  assign n10617 = ~Pg35 & Ng3929;
  assign n10618 = ~n5083 & ~n10617;
  assign n10619 = ~n10615 & ~n10618;
  assign n4945_1 = n10616 | n10619;
  assign n10621 = ~Pg35 & ~Ng4369;
  assign n10622 = ~Ng4462 & Ng4473;
  assign n10623 = ~Ng4459 & ~n10622;
  assign n10624 = n8410 & n10623;
  assign n4954_1 = ~n10621 & ~n10624;
  assign n10626 = Pg35 & ~Pg12923;
  assign n10627 = Pg35 & Ng1266;
  assign n10628 = Ng1249 & ~n10627;
  assign n10629 = ~Ng1249 & n10627;
  assign n10630 = ~n10628 & ~n10629;
  assign n4959_1 = ~n10626 & ~n10630;
  assign n10632 = Pg17604 & n4549;
  assign n10633 = Ng5689 & n10632;
  assign n10634 = n6893 & n10633;
  assign n10635 = Pg35 & ~n10634;
  assign n10636 = ~Ng5489 & n10635;
  assign n10637 = ~Pg35 & Ng5485;
  assign n10638 = ~n7207 & ~n10637;
  assign n10639 = ~n10635 & n10638;
  assign n4964_1 = ~n10636 & ~n10639;
  assign n10641 = ~Ng714 & n5897;
  assign n10642 = Pg35 & ~n10641;
  assign n10643 = Ng676 & ~n10642;
  assign n10644 = ~Ng676 & n5899_1;
  assign n10645 = ~n5900 & ~n10644;
  assign n10646 = Ng714 & ~n10645;
  assign n4969_1 = n10643 | n10646;
  assign n10648 = ~Pg35 & Ng2741;
  assign n10649 = ~Ng2748 & ~n7801;
  assign n10650 = n7718 & ~n7801;
  assign n10651 = Ng2841 & ~Ng2748;
  assign n10652 = ~n10650 & ~n10651;
  assign n10653 = ~n10649 & ~n10652;
  assign n4974 = n10648 | n10653;
  assign n10655 = Pg35 & Ng5467;
  assign n10656 = ~Ng5462 & n10655;
  assign n10657 = n10634 & n10656;
  assign n10658 = Ng5462 & ~n10655;
  assign n10659 = ~n10635 & n10658;
  assign n10660 = n4793 & ~n10634;
  assign n10661 = ~n10659 & ~n10660;
  assign n4979 = n10657 | ~n10661;
  assign n10663 = ~Pg35 & Ng4423;
  assign n10664 = ~n5409 & ~n8747;
  assign n4984_1 = n10663 | ~n10664;
  assign n10666 = Ng6561 & n7557;
  assign n10667 = n5083 & n10666;
  assign n10668 = ~Pg35 & Ng6649;
  assign n10669 = ~n10667 & ~n10668;
  assign n10670 = Pg35 & Ng6605;
  assign n10671 = ~n10666 & n10670;
  assign n4993 = ~n10669 | n10671;
  assign n10673 = ~n6959 & n7790;
  assign n10674 = n7004 & n10673;
  assign n10675 = ~Pg35 & Ng2449;
  assign n10676 = Pg35 & Ng2445;
  assign n10677 = ~n10673 & n10676;
  assign n10678 = ~n10675 & ~n10677;
  assign n4998_1 = n10674 | ~n10678;
  assign n10680 = Ng2153 & ~n6498_1;
  assign n10681 = Ng2227 & n10680;
  assign n10682 = Pg35 & ~n10681;
  assign n10683 = Ng2173 & n10682;
  assign n10684 = ~Pg35 & Ng2177;
  assign n10685 = ~n6505 & ~n10684;
  assign n10686 = ~n10682 & ~n10685;
  assign n5003 = n10683 | n10686;
  assign n10688 = Pg35 & Ng4291;
  assign n10689 = ~Pg35 & ~Ng4284;
  assign n5008 = ~n10688 & ~n10689;
  assign n10691 = n4928 & n6152;
  assign n10692 = Ng2491 & ~n10691;
  assign n10693 = Pg35 & n10692;
  assign n10694 = Ng110 & n10522;
  assign n10695 = ~Ng110 & ~n10522;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = n5842 & n10696;
  assign n10698 = n6152 & n10697;
  assign n10699 = ~Pg35 & Ng2476;
  assign n10700 = ~n10698 & ~n10699;
  assign n5012_1 = n10693 | ~n10700;
  assign n10702 = ~Pg35 & Ng4843;
  assign n10703 = Ng4849 & n10259;
  assign n10704 = n4604 & ~n5817;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n10483 & ~n10705;
  assign n5017 = n10702 | n10706;
  assign n10708 = ~Pg35 & Ng2161;
  assign n10709 = Ng2197 & ~n6498_1;
  assign n10710 = ~Ng2227 & n10709;
  assign n10711 = n6505 & n10710;
  assign n10712 = Pg35 & Ng2169;
  assign n10713 = ~n10710 & n10712;
  assign n10714 = ~n10711 & ~n10713;
  assign n5022 = n10708 | ~n10714;
  assign n10716 = Ng2279 & n9778;
  assign n10717 = ~Ng2279 & ~n9778;
  assign n10718 = ~n10716 & ~n10717;
  assign n10719 = ~n6707 & ~n10718;
  assign n10720 = ~Ng2283 & n6707;
  assign n5027 = ~n10719 & ~n10720;
  assign n10722 = n7380 & n8691;
  assign n10723 = Pg35 & ~Ng6585;
  assign n10724 = ~n10722 & n10723;
  assign n10725 = n5018 & n10722;
  assign n10726 = ~Pg35 & ~Ng6589;
  assign n10727 = ~n10725 & ~n10726;
  assign n5032 = ~n10724 & n10727;
  assign n10729 = ~Pg35 & Ng2831;
  assign n5037 = n9928 | n10729;
  assign n10731 = Ng2407 & n4981;
  assign n10732 = ~Pg35 & Ng2403;
  assign n10733 = n4980 & n8161;
  assign n10734 = ~n10732 & ~n10733;
  assign n5042 = n10731 | ~n10734;
  assign n10736 = Pg35 & Ng2868;
  assign n10737 = ~Pg35 & Ng2988;
  assign n5047_1 = n10736 | n10737;
  assign n10739 = ~Ng1632 & n8039;
  assign n10740 = ~Pg35 & Ng2763;
  assign n10741 = Ng2767 & n8036;
  assign n10742 = ~n10740 & ~n10741;
  assign n5052_1 = n10739 | ~n10742;
  assign n10744 = Ng1783 & n8434;
  assign n10745 = Ng1760 & ~n8434;
  assign n10746 = ~n8433 & ~n10745;
  assign n5057_1 = n10744 | ~n10746;
  assign n10748 = Pg35 & ~n5510;
  assign n10749 = Ng1312 & n10748;
  assign n10750 = Ng1389 & n5509;
  assign n10751 = n7243 & ~n10750;
  assign n10752 = ~Ng1351 & n8712;
  assign n10753 = ~n10751 & ~n10752;
  assign n10754 = Pg35 & ~n5506;
  assign n10755 = ~n10753 & n10754;
  assign n5065 = n10749 | n10755;
  assign n10757 = Ng5176 & n10319;
  assign n10758 = Ng5212 & ~n10757;
  assign n10759 = Pg35 & n10758;
  assign n10760 = n5083 & n10757;
  assign n10761 = ~Pg35 & Ng5260;
  assign n10762 = ~n10760 & ~n10761;
  assign n5070_1 = n10759 | ~n10762;
  assign n10764 = Pg35 & Ng4245;
  assign n10765 = ~Pg35 & Ng4249;
  assign n5075_1 = n10764 | n10765;
  assign n10767 = Pg35 & n6094;
  assign n10768 = Ng446 & n10767;
  assign n10769 = Ng645 & n6095;
  assign n5080 = n10768 | n10769;
  assign n10771 = ~Ng661 & n5884;
  assign n10772 = Pg35 & ~n10771;
  assign n10773 = ~Ng728 & ~n10772;
  assign n10774 = Pg35 & ~n5884;
  assign n10775 = ~\[4435]  & n10774;
  assign n5089_1 = ~n10773 & ~n10775;
  assign n10777 = Ng182 & n5027_1;
  assign n10778 = ~Pg35 & Ng405;
  assign n10779 = Ng446 & n8865;
  assign n10780 = ~n10778 & ~n10779;
  assign n5094_1 = n10777 | ~n10780;
  assign n10782 = ~Pg35 & Ng1124;
  assign n10783 = Ng1124 & n10175;
  assign n10784 = n6104 & n10783;
  assign n10785 = Ng1129 & n10784;
  assign n10786 = Pg35 & Ng1129;
  assign n10787 = ~n10784 & ~n10786;
  assign n10788 = ~n10785 & ~n10787;
  assign n5099 = n10782 | n10788;
  assign n10790 = Pg35 & n9515;
  assign n10791 = Ng2197 & ~n9513;
  assign n10792 = ~n10790 & n10791;
  assign n10793 = Ng2227 & n9513;
  assign n5104 = n10792 | n10793;
  assign n10795 = Ng2241 & n9781;
  assign n10796 = Ng2246 & ~n9781;
  assign n5112 = n10795 | n10796;
  assign n10798 = ~Ng1830 & ~n10445;
  assign n10799 = Pg35 & Ng1821;
  assign n10800 = Ng1825 & n10799;
  assign n10801 = ~Ng1825 & ~n10799;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = n10445 & ~n10802;
  assign n5117 = ~n10798 & ~n10803;
  assign n10805 = n5201 & n5828;
  assign n10806 = n5018 & n10805;
  assign n10807 = ~Pg35 & ~Ng3574;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = Pg35 & ~n10805;
  assign n10810 = ~Ng3590 & n10809;
  assign n5122_1 = n10808 & ~n10810;
  assign n10812 = Ng392 & n5151;
  assign n10813 = ~Pg35 & Ng401;
  assign n10814 = n5150 & n8921;
  assign n10815 = Ng854 & n10814;
  assign n10816 = ~n10813 & ~n10815;
  assign n5127 = n10812 | ~n10816;
  assign n10818 = Ng1592 & n5244;
  assign n10819 = ~Ng1592 & ~n5228;
  assign n10820 = Pg35 & ~n8835;
  assign n10821 = ~Ng1668 & n10820;
  assign n10822 = ~n10819 & n10821;
  assign n5132_1 = n10818 | n10822;
  assign n10824 = Ng6505 & n7313;
  assign n10825 = Ng6541 & ~n7313;
  assign n5137_1 = n10824 | n10825;
  assign n10827 = ~Pg35 & Ng1205;
  assign n10828 = Pg35 & Ng1221;
  assign n10829 = ~n7499 & ~n10828;
  assign n10830 = ~n7500 & ~n10829;
  assign n5142_1 = n10827 | n10830;
  assign n10832 = n7650 & n9706;
  assign n10833 = n5083 & n10832;
  assign n10834 = ~Pg35 & Ng5893;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = Pg35 & Ng5921;
  assign n10837 = ~n10832 & n10836;
  assign n5147_1 = ~n10835 | n10837;
  assign n10839 = ~Pg35 & \[4436] ;
  assign n10840 = ~Ng341 & n8272;
  assign n10841 = n8276 & n10840;
  assign n5152_1 = n10839 | n10841;
  assign n10843 = ~Pg35 & Ng142;
  assign n10844 = ~Ng146 & ~n6880;
  assign n10845 = ~n7264 & ~n10844;
  assign n10846 = n7270 & n10845;
  assign n5157 = n10843 | n10846;
  assign n10848 = n4928 & n5841;
  assign n10849 = Ng1932 & ~n10848;
  assign n10850 = Pg35 & n10849;
  assign n10851 = Ng110 & n9536;
  assign n10852 = ~Ng110 & ~n9536;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = n5841 & n10853;
  assign n10855 = n5842 & n10854;
  assign n10856 = ~Pg35 & Ng1917;
  assign n10857 = ~n10855 & ~n10856;
  assign n5166 = n10850 | ~n10857;
  assign n10859 = ~Pg35 & Ng1632;
  assign n10860 = n6250 & n8572;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = Ng1624 & n8570;
  assign n10863 = ~n9632 & ~n10862;
  assign n5171 = ~n10861 | ~n10863;
  assign n10865 = ~Ng5109 & Pg9497;
  assign n10866 = ~Ng5062 & ~n10865;
  assign n10867 = Pg35 & ~Pg9553;
  assign n10868 = ~n10866 & n10867;
  assign n10869 = ~Pg35 & Ng5109;
  assign n5176_1 = n10868 | n10869;
  assign n10871 = ~Ng5703 & ~Ng5644;
  assign n10872 = Ng5583 & Pg14694;
  assign n10873 = n10871 & n10872;
  assign n10874 = Pg12300 & ~Ng5689;
  assign n10875 = ~Pg12300 & Ng5689;
  assign n10876 = ~n10874 & ~n10875;
  assign n10877 = ~Ng5703 & Ng5644;
  assign n10878 = Ng5615 & Pg17580;
  assign n10879 = n10877 & n10878;
  assign n10880 = ~n10876 & ~n10879;
  assign n10881 = Ng5703 & ~Ng5644;
  assign n10882 = Ng5599 & n10881;
  assign n10883 = Pg17711 & n10882;
  assign n10884 = n10880 & ~n10883;
  assign n10885 = ~n10873 & n10884;
  assign n10886 = Ng5575 & Pg14694;
  assign n10887 = n10877 & n10886;
  assign n10888 = Pg17711 & n4549;
  assign n10889 = Ng5591 & n10888;
  assign n10890 = Ng5607 & Pg17580;
  assign n10891 = n10871 & n10890;
  assign n10892 = n10876 & ~n10891;
  assign n10893 = ~n10889 & n10892;
  assign n10894 = ~n10887 & n10893;
  assign n10895 = ~n10885 & ~n10894;
  assign n10896 = Ng5611 & Pg17678;
  assign n10897 = Ng5559 & Pg17604;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = n10881 & ~n10898;
  assign n10900 = Ng5595 & n10871;
  assign n10901 = Pg14635 & n10900;
  assign n10902 = ~n10899 & ~n10901;
  assign n10903 = Ng5579 & Pg17813;
  assign n10904 = Pg12300 & Ng5563;
  assign n10905 = ~n10903 & ~n10904;
  assign n10906 = n4549 & ~n10905;
  assign n10907 = Ng5555 & Pg13049;
  assign n10908 = Ng5567 & Ng5685;
  assign n10909 = ~n10907 & ~n10908;
  assign n10910 = n10877 & ~n10909;
  assign n10911 = ~Ng5689 & ~n10910;
  assign n10912 = ~n10906 & n10911;
  assign n10913 = n10902 & n10912;
  assign n10914 = Ng5543 & Pg13049;
  assign n10915 = Ng5551 & Ng5685;
  assign n10916 = ~n10914 & ~n10915;
  assign n10917 = n10871 & ~n10916;
  assign n10918 = Ng5571 & Pg17813;
  assign n10919 = Pg12300 & Ng5547;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = n10881 & ~n10920;
  assign n10922 = Ng5689 & ~n10921;
  assign n10923 = Ng5587 & n10877;
  assign n10924 = Pg14635 & n10923;
  assign n10925 = Ng5603 & n4549;
  assign n10926 = Pg17678 & n10925;
  assign n10927 = ~n10924 & ~n10926;
  assign n10928 = n10922 & n10927;
  assign n10929 = ~n10917 & n10928;
  assign n10930 = ~n10913 & ~n10929;
  assign n10931 = ~n10895 & ~n10930;
  assign n10932 = ~Ng5619 & n10931;
  assign n10933 = ~n10633 & n10931;
  assign n10934 = n6904 & ~n10933;
  assign n10935 = ~n10932 & n10934;
  assign n10936 = ~Ng5462 & n10935;
  assign n10937 = Pg35 & Ng5462;
  assign n10938 = n10633 & ~n10932;
  assign n10939 = n6893 & ~n10933;
  assign n10940 = ~n10938 & n10939;
  assign n10941 = n10937 & ~n10940;
  assign n10942 = ~Pg35 & Ng5467;
  assign n10943 = ~n10941 & ~n10942;
  assign n5181_1 = n10936 | ~n10943;
  assign n5186_1 = Pg35 & Ng2689;
  assign n10946 = ~Pg35 & Ng6565;
  assign n10947 = Ng6565 & Ng6561;
  assign n10948 = ~n4288_1 & ~n10947;
  assign n10949 = ~n7713 & ~n10948;
  assign n10950 = ~n4714 & n10949;
  assign n5191 = n10946 | n10950;
  assign n10952 = Ng1604 & n7902;
  assign n10953 = Pg35 & n10952;
  assign n10954 = ~Pg35 & Ng1657;
  assign n10955 = Ng1624 & ~Ng1648;
  assign n10956 = Ng1616 & n10955;
  assign n10957 = Ng1620 & Pg31863;
  assign n10958 = Ng1608 & n7369;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = Ng1600 & n8571;
  assign n10961 = ~Ng1624 & Ng1612;
  assign n10962 = ~Ng1657 & n10961;
  assign n10963 = ~n10960 & ~n10962;
  assign n10964 = n10959 & n10963;
  assign n10965 = ~n10956 & n10964;
  assign n10966 = n9628 & ~n10965;
  assign n10967 = Ng1677 & n8570;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = ~n10954 & n10968;
  assign n5196_1 = n10953 | ~n10969;
  assign n10971 = Pg35 & n6947;
  assign n10972 = ~Ng2060 & n10971;
  assign n10973 = ~Ng2051 & n10972;
  assign n10974 = n4638 & n6947;
  assign n10975 = n5843 & n10974;
  assign n10976 = ~Pg35 & Ng2036;
  assign n10977 = Pg35 & Ng2028;
  assign n10978 = ~n6948 & n10977;
  assign n10979 = ~n10976 & ~n10978;
  assign n10980 = ~n10975 & n10979;
  assign n5201_1 = n10973 | ~n10980;
  assign n10982 = Ng2671 & ~n8993;
  assign n10983 = Pg35 & ~Ng2661;
  assign n10984 = ~Ng2667 & n10983;
  assign n10985 = Ng2667 & ~n10983;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = n8993 & ~n10986;
  assign n5206_1 = n10982 | n10987;
  assign n10989 = ~Pg35 & Ng1589;
  assign n10990 = Pg17423 & ~Pg12923;
  assign n10991 = ~Pg10527 & ~Pg17423;
  assign n10992 = Pg35 & ~n10991;
  assign n10993 = ~n10990 & n10992;
  assign n5211_1 = n10989 | n10993;
  assign n10995 = ~Pg35 & Ng4411;
  assign n10996 = ~n6865 & ~n6867;
  assign n5215_1 = n10995 | ~n10996;
  assign n10998 = ~Pg35 & Ng1844;
  assign n10999 = Pg35 & ~Ng1848;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = n8858 & n11000;
  assign n11002 = ~Ng1848 & ~n8858;
  assign n5219_1 = ~n11001 & ~n11002;
  assign n11004 = Pg35 & \[4434] ;
  assign n11005 = Ng5097 & ~n6786;
  assign n11006 = ~n11004 & n11005;
  assign n11007 = n11004 & ~n11005;
  assign n5224_1 = n11006 | n11007;
  assign n11009 = Ng5485 & n10635;
  assign n11010 = Ng5481 & ~n9968;
  assign n11011 = ~Ng5481 & n9968;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = ~n10635 & ~n11012;
  assign n5229_1 = n11009 | n11013;
  assign n11015 = ~Ng2741 & ~n7800;
  assign n11016 = n10650 & ~n11015;
  assign n11017 = ~Pg35 & Ng2735;
  assign n5234_1 = n11016 | n11017;
  assign n11019 = Ng2619 & n5329;
  assign n11020 = Ng2587 & n11019;
  assign n11021 = Ng2567 & n11020;
  assign n11022 = Pg35 & n11021;
  assign n11023 = ~Pg35 & Ng2619;
  assign n11024 = ~Ng2587 & Ng2575;
  assign n11025 = ~Ng2619 & n11024;
  assign n11026 = Ng2571 & n8556;
  assign n11027 = Ng2563 & n5331;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = Ng2583 & n4634;
  assign n11030 = Ng2587 & Ng2579;
  assign n11031 = ~Ng2610 & n11030;
  assign n11032 = ~n11029 & ~n11031;
  assign n11033 = n11028 & n11032;
  assign n11034 = ~n11025 & n11033;
  assign n11035 = n8463 & ~n11034;
  assign n11036 = Ng2638 & n5330;
  assign n11037 = ~n11035 & ~n11036;
  assign n11038 = ~n11023 & n11037;
  assign n5242_1 = n11022 | ~n11038;
  assign n11040 = n6200 & n9023;
  assign n11041 = Pg35 & ~n11040;
  assign n11042 = Ng4122 & n11041;
  assign n11043 = ~Pg35 & Ng4119;
  assign n11044 = ~n9029 & ~n11043;
  assign n11045 = ~n11041 & ~n11044;
  assign n5247_1 = n11042 | n11045;
  assign n11047 = n5912 & ~n5914_1;
  assign n11048 = Ng4322 & n11047;
  assign n11049 = ~Pg35 & Ng4311;
  assign n11050 = ~Ng4322 & n5915;
  assign n11051 = ~n11049 & ~n11050;
  assign n5252_1 = n11048 | ~n11051;
  assign n11053 = n6426 & n6754;
  assign n11054 = Pg35 & ~n11053;
  assign n11055 = Ng5941 & n11054;
  assign n11056 = ~Pg35 & Ng5925;
  assign n11057 = ~n5083 & ~n11056;
  assign n11058 = ~n11054 & ~n11057;
  assign n5257_1 = n11055 | n11058;
  assign n11060 = Ng2102 & n5664;
  assign n11061 = Ng2108 & ~n5664;
  assign n5262_1 = n11060 | n11061;
  assign n11063 = ~Pg35 & Ng1592;
  assign n11064 = n4575_1 & Pg33533;
  assign n11065 = Ng112 & Pg31862;
  assign n11066 = ~Ng112 & ~Pg31862;
  assign n11067 = ~n11065 & ~n11066;
  assign n11068 = n11064 & n11067;
  assign n11069 = n5842 & n11068;
  assign n11070 = ~n11063 & ~n11069;
  assign n11071 = n4928 & n11064;
  assign n11072 = Ng1644 & ~n11071;
  assign n11073 = Pg35 & n11072;
  assign n5274_1 = ~n11070 | n11073;
  assign n11075 = ~Pg35 & Ng590;
  assign n11076 = Ng595 & n5737;
  assign n11077 = ~n5753 & ~n11076;
  assign n11078 = ~n5754 & ~n11077;
  assign n5279 = n11075 | n11078;
  assign n11080 = Ng2208 & n5261;
  assign n11081 = Ng2217 & n5259;
  assign n11082 = ~n11080 & ~n11081;
  assign n11083 = ~Pg35 & Ng2223;
  assign n11084 = ~n10039 & ~n11083;
  assign n5284_1 = ~n11082 | ~n11084;
  assign n11086 = ~Ng1404 & n10626;
  assign n11087 = Pg35 & Ng1395;
  assign n11088 = ~Ng1404 & ~n11087;
  assign n11089 = ~n10626 & ~n11088;
  assign n11090 = Pg35 & ~Pg19357;
  assign n11091 = ~n11089 & ~n11090;
  assign n5289 = n11086 | ~n11091;
  assign n11093 = n4928 & n10974;
  assign n11094 = Ng2066 & ~n11093;
  assign n11095 = Pg35 & n11094;
  assign n11096 = ~Ng2051 & Ng2060;
  assign n11097 = Ng110 & n11096;
  assign n11098 = ~Ng110 & ~n11096;
  assign n11099 = ~n11097 & ~n11098;
  assign n11100 = n5842 & n11099;
  assign n11101 = n10974 & n11100;
  assign n11102 = ~Pg35 & Ng2051;
  assign n11103 = ~n11101 & ~n11102;
  assign n5294 = n11095 | ~n11103;
  assign n11105 = Ng1152 & n5813;
  assign n11106 = Ng1146 & ~n5813;
  assign n5299_1 = n11105 | n11106;
  assign n11108 = ~Pg35 & ~Ng5236;
  assign n11109 = n4708_1 & n9551;
  assign n11110 = n5018 & n11109;
  assign n11111 = Pg35 & ~Ng5252;
  assign n11112 = ~n11109 & n11111;
  assign n11113 = ~n11110 & ~n11112;
  assign n5304_1 = ~n11108 & n11113;
  assign n11115 = ~Pg35 & Ng2246;
  assign n11116 = ~n6505 & ~n11115;
  assign n11117 = n9781 & n11116;
  assign n11118 = ~Ng2165 & ~n9781;
  assign n5309_1 = ~n11117 & ~n11118;
  assign n11120 = ~Pg35 & Ng2563;
  assign n11121 = Ng2599 & ~n5533;
  assign n11122 = ~Ng2629 & n11121;
  assign n11123 = n5543 & n11122;
  assign n11124 = Pg35 & Ng2571;
  assign n11125 = ~n11122 & n11124;
  assign n11126 = ~n11123 & ~n11125;
  assign n5314 = n11120 | ~n11126;
  assign n11128 = ~Pg35 & Ng5170;
  assign n11129 = n5599 & n6412;
  assign n5319_1 = n11128 | n11129;
  assign n11131 = ~Ng1211 & ~n7501;
  assign n11132 = n7503 & ~n11131;
  assign n11133 = ~Pg35 & Ng1216;
  assign n5327_1 = n11132 | n11133;
  assign n11135 = ~Ng2595 & n8039;
  assign n11136 = ~Pg35 & Ng2823;
  assign n11137 = ~n8036 & ~n11136;
  assign n11138 = ~n6715 & ~n11137;
  assign n5332_1 = n11135 | n11138;
  assign n11140 = Ng4859 & n10259;
  assign n11141 = n10258 & n10484;
  assign n11142 = ~Pg35 & Ng4854;
  assign n11143 = ~n11141 & ~n11142;
  assign n5340_1 = n11140 | ~n11143;
  assign n11145 = Ng424 & n5151;
  assign n11146 = Ng411 & ~n5151;
  assign n5345_1 = n11145 | n11146;
  assign n11148 = ~Ng1274 & n7939;
  assign n11149 = Pg35 & ~n11148;
  assign n11150 = Ng1270 & ~n11149;
  assign n11151 = n5591 & ~n9468;
  assign n11152 = Ng1274 & n11151;
  assign n5350_1 = n11150 | n11152;
  assign n11154 = Ng2799 & ~n4928;
  assign n11155 = n4931 & ~n6719;
  assign n11156 = ~n11154 & n11155;
  assign n11157 = Ng2803 & ~n4931;
  assign n11158 = Pg35 & ~n11157;
  assign n11159 = ~n11156 & n11158;
  assign n11160 = ~Pg35 & ~Ng2807;
  assign n5362_1 = ~n11159 & ~n11160;
  assign n11162 = Ng1816 & n8858;
  assign n11163 = Ng1821 & ~n8858;
  assign n5367_1 = n11162 | n11163;
  assign n11165 = ~Pg35 & Ng2495;
  assign n11166 = ~Ng2509 & n6959;
  assign n11167 = Ng1589 & ~n6956;
  assign n11168 = ~n7002 & ~n11167;
  assign n11169 = Ng2509 & ~n7007;
  assign n11170 = n11168 & n11169;
  assign n11171 = ~n11168 & ~n11169;
  assign n11172 = ~n11170 & ~n11171;
  assign n11173 = ~n6959 & n11172;
  assign n11174 = Pg35 & ~n11173;
  assign n11175 = ~n11166 & n11174;
  assign n5372_1 = n11165 | n11175;
  assign n11177 = ~Pg35 & Ng5069;
  assign n5377_1 = n7590 | n11177;
  assign n11179 = ~Pg35 & Ng1266;
  assign n11180 = Ng1280 & n5591;
  assign n11181 = ~n7816 & ~n11180;
  assign n11182 = ~n7817 & ~n11181;
  assign n5382_1 = n11179 | n11182;
  assign n11184 = ~Pg35 & ~Ng6617;
  assign n11185 = n7103 & n7557;
  assign n11186 = Pg35 & ~Ng6633;
  assign n11187 = ~n11185 & n11186;
  assign n11188 = n5018 & n11185;
  assign n11189 = ~n11187 & ~n11188;
  assign n5394_1 = ~n11184 & n11189;
  assign n11191 = Ng5124 & n6143_1;
  assign n11192 = Pg35 & Ng5120;
  assign n11193 = ~Ng5115 & n11192;
  assign n11194 = Ng5115 & ~n11192;
  assign n11195 = ~n11193 & ~n11194;
  assign n11196 = ~n6143_1 & ~n11195;
  assign n5399_1 = n11191 | n11196;
  assign n11198 = n5498 & n5849;
  assign n11199 = Pg35 & ~n11198;
  assign n11200 = ~Pg35 & ~Ng6287;
  assign n11201 = ~n5018 & ~n11200;
  assign n11202 = ~n11199 & ~n11201;
  assign n11203 = ~Ng6303 & n11199;
  assign n5407_1 = ~n11202 & ~n11203;
  assign n11205 = ~Pg35 & Ng5057;
  assign n5412 = n4921 | n11205;
  assign n11207 = Pg35 & Ng2994;
  assign n11208 = ~Pg35 & Ng2999;
  assign n5417_1 = n11207 | n11208;
  assign n11210 = Ng650 & n6095;
  assign n11211 = ~Pg35 & Ng699;
  assign n11212 = Ng681 & n10767;
  assign n11213 = ~n11211 & ~n11212;
  assign n5422_1 = n11210 | ~n11213;
  assign n11215 = Ng1636 & n5244;
  assign n11216 = ~Pg35 & Ng1644;
  assign n11217 = Ng1592 & ~n5227;
  assign n11218 = n10820 & n11217;
  assign n11219 = ~n11216 & ~n11218;
  assign n5427_1 = n11215 | ~n11219;
  assign n11221 = ~Pg35 & ~Ng3893;
  assign n11222 = n8079 & n9940;
  assign n11223 = n5018 & n11222;
  assign n11224 = Pg35 & ~Ng3921;
  assign n11225 = ~n11222 & n11224;
  assign n11226 = ~n11223 & ~n11225;
  assign n5432 = ~n11221 & n11226;
  assign n11228 = Pg35 & Ng2093;
  assign n11229 = ~Ng2079 & ~n10395;
  assign n11230 = n6947 & ~n11229;
  assign n11231 = n11228 & ~n11230;
  assign n11232 = ~n10395 & n11228;
  assign n11233 = Pg35 & ~n6947;
  assign n11234 = Ng2079 & ~n11233;
  assign n11235 = ~n11232 & n11234;
  assign n5437_1 = n11231 | n11235;
  assign n11237 = ~Pg35 & Ng6727;
  assign n11238 = ~Ng6736 & n6466;
  assign n5442_1 = n11237 | n11238;
  assign n11240 = ~Pg35 & Ng1521;
  assign n11241 = Ng1526 & n9267;
  assign n11242 = ~Ng1306 & ~n11241;
  assign n11243 = ~Ng1339 & n11241;
  assign n11244 = Pg35 & ~n11243;
  assign n11245 = ~n11242 & n11244;
  assign n5447 = n11240 | n11245;
  assign n11247 = ~Pg35 & Ng1052;
  assign n11248 = Ng1061 & n6941;
  assign n11249 = Pg35 & Ng1061;
  assign n11250 = ~n6941 & ~n11249;
  assign n11251 = ~Ng979 & ~n11250;
  assign n11252 = ~n11248 & n11251;
  assign n5452_1 = n11247 | n11252;
  assign n11254 = Ng3462 & n5213;
  assign n11255 = Ng3498 & ~n5213;
  assign n5457 = n11254 | n11255;
  assign n11257 = ~Pg35 & Ng2169;
  assign n11258 = n4590 & ~n6498_1;
  assign n11259 = Pg35 & ~n11258;
  assign n11260 = ~n6505 & ~n11259;
  assign n11261 = ~n11257 & n11260;
  assign n11262 = ~Ng2181 & n11259;
  assign n5462_1 = ~n11261 & ~n11262;
  assign n11264 = ~Pg35 & Ng1141;
  assign n11265 = Ng1141 & n5812;
  assign n11266 = n6104 & n11265;
  assign n11267 = Ng956 & n11266;
  assign n11268 = Pg35 & Ng956;
  assign n11269 = ~n11266 & ~n11268;
  assign n11270 = ~n11267 & ~n11269;
  assign n5467_1 = n11264 | n11270;
  assign n11272 = n4593 & ~n5063;
  assign n11273 = n5070 & n11272;
  assign n11274 = ~Pg35 & Ng1744;
  assign n11275 = Pg35 & Ng1756;
  assign n11276 = ~n11272 & n11275;
  assign n11277 = ~n11274 & ~n11276;
  assign n5472_1 = n11273 | ~n11277;
  assign n11279 = Ng5849 & ~n4718_1;
  assign n11280 = n5018 & n11279;
  assign n11281 = n5083 & ~n11279;
  assign n5477_1 = n11280 | n11281;
  assign n11283 = n9007 & n9022;
  assign n11284 = Pg35 & ~n11283;
  assign n11285 = Ng4112 & n11284;
  assign n11286 = Ng4145 & ~n11284;
  assign n5482_1 = n11285 | n11286;
  assign n11288 = Pg35 & ~n11020;
  assign n11289 = Ng2681 & n10244;
  assign n11290 = ~Ng2681 & ~n10244;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = ~n11288 & ~n11291;
  assign n11293 = ~Ng2685 & n11288;
  assign n5487_1 = ~n11292 & ~n11293;
  assign n11295 = n9516 & n10680;
  assign n11296 = ~Pg35 & Ng2204;
  assign n11297 = Ng2197 & n9513;
  assign n11298 = ~n11296 & ~n11297;
  assign n5492_1 = n11295 | ~n11298;
  assign n11300 = Ng2421 & n6965;
  assign n11301 = ~Ng2421 & ~n10222;
  assign n11302 = ~Ng2495 & n6962;
  assign n11303 = ~n11301 & n11302;
  assign n5497_1 = n11300 | n11303;
  assign n11305 = ~Pg35 & ~Ng1041;
  assign n11306 = Ng1046 & ~n8104;
  assign n11307 = n5610 & n8104;
  assign n11308 = Pg35 & ~n11307;
  assign n11309 = ~n11306 & n11308;
  assign n5502_1 = ~n11305 & ~n11309;
  assign n11311 = ~Pg35 & Ng528;
  assign n11312 = ~Ng482 & ~n5356;
  assign n11313 = n5358 & ~n11312;
  assign n11314 = ~n5349 & ~n11313;
  assign n5507_1 = n11311 | ~n11314;
  assign n11316 = Ng4388 & n6865;
  assign n5512_1 = Ng4405 | n11316;
  assign n11318 = ~Pg7946 & ~Ng1514;
  assign n11319 = ~n9267 & ~n11318;
  assign n11320 = ~n8717 & ~n11319;
  assign n5517_1 = Pg35 & ~n11320;
  assign n11322 = ~Ng6565 & ~n7713;
  assign n11323 = Pg35 & ~n11322;
  assign n11324 = Ng6561 & ~n11323;
  assign n11325 = Ng6565 & n7715;
  assign n5527_1 = n11324 | n11325;
  assign n11327 = Pg35 & Ng2950;
  assign n11328 = ~Pg35 & Ng2936;
  assign n5532_1 = n11327 | n11328;
  assign n11330 = ~Ng1345 & n5506;
  assign n11331 = Pg35 & ~n11330;
  assign n11332 = ~n7248 & n11331;
  assign n11333 = ~Pg35 & Ng1351;
  assign n5537_1 = n11332 | n11333;
  assign n11335 = Ng6533 & n7313;
  assign n11336 = Ng6527 & ~n7313;
  assign n5542 = n11335 | n11336;
  assign n5550_1 = Pg35 & Ng4727;
  assign n11339 = ~Pg14828 & ~Pg17778;
  assign n11340 = ~n6461 & ~n11339;
  assign n11341 = Pg35 & ~Pg17722;
  assign n11342 = ~Pg13099 & ~Pg17688;
  assign n11343 = n11341 & n11342;
  assign n5555_1 = ~n11340 & n11343;
  assign n11345 = Ng1536 & ~n8718;
  assign n11346 = Pg35 & ~n8715;
  assign n11347 = ~n11345 & n11346;
  assign n11348 = ~Pg35 & ~Ng1532;
  assign n5559_1 = ~n11347 & ~n11348;
  assign n11350 = n6918 & n7216;
  assign n11351 = Pg35 & ~n11350;
  assign n11352 = ~Pg35 & ~Ng3925;
  assign n11353 = ~n5018 & ~n11352;
  assign n11354 = ~n11351 & ~n11353;
  assign n11355 = ~Ng3941 & n11351;
  assign n5564_1 = ~n11354 & ~n11355;
  assign n11357 = ~Pg35 & ~Ng358;
  assign n11358 = Ng370 & ~n5808;
  assign n11359 = ~Ng370 & n5808;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = Pg35 & n11360;
  assign n5569_1 = ~n11357 & ~n11361;
  assign n11363 = ~Pg35 & Ng5689;
  assign n11364 = ~Ng5698 & n8653;
  assign n5574 = n11363 | n11364;
  assign n11366 = Ng1854 & n10999;
  assign n11367 = ~Ng1854 & ~n10999;
  assign n11368 = ~n11366 & ~n11367;
  assign n11369 = ~n10001 & ~n11368;
  assign n11370 = ~Ng1858 & n10001;
  assign n5579_1 = ~n11369 & ~n11370;
  assign n11372 = Ng446 & n7393;
  assign n11373 = Ng872 & n7390;
  assign n11374 = ~Pg35 & Ng246;
  assign n11375 = ~n11373 & ~n11374;
  assign n5584_1 = n11372 | ~n11375;
  assign n11377 = n6658 & n8807;
  assign n11378 = Pg35 & ~n11377;
  assign n11379 = ~Pg35 & ~Ng3191;
  assign n11380 = ~n5018 & ~n11379;
  assign n11381 = ~n11378 & ~n11380;
  assign n11382 = ~Ng3219 & n11378;
  assign n5589_1 = ~n11381 & ~n11382;
  assign n11384 = ~Pg35 & Ng1792;
  assign n11385 = Ng1740 & n10000;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = Pg35 & n6185;
  assign n11388 = Ng1748 & ~Ng1792;
  assign n11389 = ~Ng1760 & n11388;
  assign n11390 = Ng1744 & n6188;
  assign n11391 = Ng1756 & n4659;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = Ng1736 & n8428;
  assign n11394 = Ng1760 & ~Ng1783;
  assign n11395 = Ng1752 & n11394;
  assign n11396 = ~n11393 & ~n11395;
  assign n11397 = n11392 & n11396;
  assign n11398 = ~n11389 & n11397;
  assign n11399 = n11387 & ~n11398;
  assign n11400 = Ng1811 & n8434;
  assign n11401 = ~n11399 & ~n11400;
  assign n5594 = ~n11386 | ~n11401;
  assign n11403 = ~Pg35 & ~Ng6605;
  assign n11404 = n4713 & n8691;
  assign n11405 = ~n5018 & n11404;
  assign n11406 = Pg35 & ~Ng6601;
  assign n11407 = ~n11404 & ~n11406;
  assign n11408 = ~n11405 & ~n11407;
  assign n5599_1 = ~n11403 & ~n11408;
  assign n11410 = Ng2495 & n6960;
  assign n11411 = Pg35 & ~n11410;
  assign n11412 = Ng2441 & n11411;
  assign n11413 = ~Pg35 & Ng2445;
  assign n11414 = ~n7004 & ~n11413;
  assign n11415 = ~n11411 & ~n11414;
  assign n5604_1 = n11412 | n11415;
  assign n11417 = ~Pg35 & Ng1955;
  assign n11418 = ~n4960 & ~n11417;
  assign n11419 = n9768 & n11418;
  assign n11420 = ~Ng1874 & ~n9768;
  assign n5609_1 = ~n11419 & ~n11420;
  assign n11422 = ~Pg35 & Ng4340;
  assign n11423 = ~Ng4349 & ~n5561;
  assign n11424 = ~n5309 & ~n11423;
  assign n11425 = Pg35 & n11424;
  assign n11426 = ~n5562 & n11425;
  assign n5614_1 = n11422 | n11426;
  assign n11428 = n7753 & n8691;
  assign n11429 = n5083 & n11428;
  assign n11430 = ~Pg35 & Ng6573;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = Pg35 & Ng6581;
  assign n11433 = ~n11428 & n11432;
  assign n5619_1 = ~n11431 | n11433;
  assign n11435 = ~Ng6573 & n10947;
  assign n11436 = n5083 & n11435;
  assign n11437 = ~Pg35 & Ng6645;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = Pg35 & Ng6597;
  assign n11440 = ~n11435 & n11439;
  assign n5624 = ~n11438 | n11440;
  assign n11442 = n4705 & n5634;
  assign n11443 = n5018 & n11442;
  assign n11444 = ~Pg35 & ~Ng3594;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = Pg35 & ~n11442;
  assign n11447 = ~Ng3610 & n11446;
  assign n5629 = n11445 & ~n11447;
  assign n11449 = ~Ng2890 & n9852;
  assign n11450 = ~Pg35 & ~Ng2873;
  assign n5634_1 = ~n11449 & ~n11450;
  assign n11452 = ~Ng1978 & ~n9768;
  assign n11453 = Ng1974 & n5302;
  assign n11454 = ~Ng1974 & ~n5302;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = n9768 & ~n11455;
  assign n5639 = ~n11452 & ~n11456;
  assign n11458 = Ng1668 & n11217;
  assign n11459 = Pg35 & ~n11458;
  assign n11460 = Ng1612 & n11459;
  assign n11461 = ~Pg35 & Ng1616;
  assign n11462 = ~n5237 & ~n11461;
  assign n11463 = ~n11459 & ~n11462;
  assign n5644_1 = n11460 | n11463;
  assign n11465 = Pg35 & ~Ng2856;
  assign n11466 = n5799 & n11465;
  assign n11467 = ~Pg35 & ~Ng2848;
  assign n5654_1 = ~n11466 & ~n11467;
  assign n11469 = ~Pg35 & Ng1978;
  assign n11470 = ~n8230 & ~n11469;
  assign n11471 = n9768 & n11470;
  assign n11472 = ~Ng1982 & ~n9768;
  assign n5659 = ~n11471 & ~n11472;
  assign n11474 = n5042_1 & n10319;
  assign n11475 = Pg35 & ~n11474;
  assign n11476 = Ng5228 & n11475;
  assign n11477 = ~Pg35 & Ng5200;
  assign n11478 = ~n5083 & ~n11477;
  assign n11479 = ~n11475 & ~n11478;
  assign n5667 = n11476 | n11479;
  assign n11481 = ~Ng4064 & Ng4057;
  assign n11482 = n9023 & n11481;
  assign n11483 = Pg35 & ~n11482;
  assign n11484 = Ng4119 & n11483;
  assign n11485 = ~Pg35 & Ng4116;
  assign n11486 = ~n9029 & ~n11485;
  assign n11487 = ~n11483 & ~n11486;
  assign n5672 = n11484 | n11487;
  assign n11489 = Pg35 & n6876;
  assign n5677_1 = Ng6386 & ~n11489;
  assign n11491 = ~n8707 & ~n8717;
  assign n11492 = ~Ng1542 & ~n8706;
  assign n11493 = Pg35 & ~n11492;
  assign n11494 = n11491 & n11493;
  assign n11495 = ~Pg35 & Ng1536;
  assign n5682_1 = n11494 | n11495;
  assign n11497 = ~n4901 & ~n4908;
  assign n11498 = n7591 & n11497;
  assign n11499 = Ng5033 & n11498;
  assign n11500 = ~n4901 & ~n7832;
  assign n11501 = ~Ng5033 & ~n11500;
  assign n11502 = ~Pg35 & Ng5029;
  assign n11503 = ~n11501 & ~n11502;
  assign n5696 = n11499 | ~n11503;
  assign n11505 = Pg35 & Ng4717;
  assign n11506 = ~Pg35 & Ng4732;
  assign n5701_1 = n11505 | n11506;
  assign n11508 = Ng1559 & n7548;
  assign n11509 = ~Ng1554 & ~n11508;
  assign n11510 = Pg35 & ~n7766;
  assign n11511 = ~n11509 & n11510;
  assign n11512 = ~Pg35 & Ng1559;
  assign n5706_1 = n11511 | n11512;
  assign n11514 = Ng3849 & ~n4734;
  assign n11515 = n5018 & n11514;
  assign n11516 = n5083 & ~n11514;
  assign n5711 = n11515 | n11516;
  assign n11518 = ~Ng3155 & ~Ng3161;
  assign n11519 = ~Ng3167 & n11518;
  assign n11520 = n6081 & n11519;
  assign n11521 = Pg35 & ~n11520;
  assign n11522 = ~Pg35 & ~Ng3203;
  assign n11523 = ~n5018 & ~n11522;
  assign n11524 = ~n11521 & ~n11523;
  assign n11525 = ~Ng3199 & n11521;
  assign n5719_1 = ~n11524 & ~n11525;
  assign n11527 = Ng5841 & n6562;
  assign n11528 = ~Ng5841 & ~n6562;
  assign n11529 = ~n11527 & ~n11528;
  assign n11530 = ~n5050 & ~n11529;
  assign n11531 = ~Ng5845 & n5050;
  assign n5724_1 = ~n11530 & ~n11531;
  assign n11533 = ~n5817 & n6593;
  assign n11534 = ~Ng4975 & n11533;
  assign n11535 = Ng4975 & n6595;
  assign n11536 = ~Pg35 & Ng4966;
  assign n11537 = ~n11535 & ~n11536;
  assign n5729 = n11534 | ~n11537;
  assign n11539 = ~Pg35 & Ng785;
  assign n11540 = Ng790 & n5145;
  assign n11541 = ~n5141 & ~n11540;
  assign n11542 = ~n5142 & ~n11541;
  assign n5734_1 = n11539 | n11542;
  assign n11544 = Ng5869 & n6754;
  assign n11545 = Pg35 & ~Ng5913;
  assign n11546 = ~n11544 & n11545;
  assign n11547 = n5018 & n11544;
  assign n11548 = ~Pg35 & ~Ng5957;
  assign n11549 = ~n11547 & ~n11548;
  assign n5739 = ~n11546 & n11549;
  assign n11551 = Pg35 & ~n4654;
  assign n11552 = ~n5838 & ~n11551;
  assign n11553 = Ng1902 & ~n11552;
  assign n11554 = ~Pg35 & Ng1882;
  assign n11555 = Pg35 & ~n10424;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = n11552 & ~n11556;
  assign n5744_1 = n11553 | n11557;
  assign n11559 = Ng6163 & n5387;
  assign n11560 = Pg35 & Ng6159;
  assign n11561 = ~Ng6154 & n11560;
  assign n11562 = Ng6154 & ~n11560;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = ~n5387 & ~n11563;
  assign n5749_1 = n11559 | n11564;
  assign n11566 = ~Ng4125 & n9816;
  assign n5754_1 = n9818 | n11566;
  assign n11568 = Ng4821 & n6894;
  assign n11569 = ~Pg35 & Ng5619;
  assign n11570 = ~n11568 & ~n11569;
  assign n5759 = n10935 | ~n11570;
  assign n11572 = Ng4939 & n9130;
  assign n11573 = ~Ng3343 & ~Ng3352;
  assign n11574 = ~Ng3347 & Ng3352;
  assign n11575 = ~n11573 & ~n11574;
  assign n11576 = ~Ng3288 & ~n11575;
  assign n11577 = Ng3288 & n11575;
  assign n11578 = ~Ng4939 & ~n11577;
  assign n11579 = ~n11576 & n11578;
  assign n11580 = n5671 & n9195;
  assign n11581 = ~n11579 & n11580;
  assign n5764 = n11572 | n11581;
  assign n11583 = Ng990 & ~n8966;
  assign n11584 = ~Ng990 & n8966;
  assign n5769 = n11583 | n11584;
  assign n11586 = n4730 & n11519;
  assign n11587 = Pg35 & ~n11586;
  assign n11588 = Ng3207 & n11587;
  assign n11589 = ~Pg35 & Ng3211;
  assign n11590 = ~n5083 & ~n11589;
  assign n11591 = ~n11587 & ~n11590;
  assign n5773 = n11588 | n11591;
  assign n11593 = n4730 & n5396;
  assign n11594 = n5083 & n11593;
  assign n11595 = ~Pg35 & Ng3243;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = Pg35 & Ng3259;
  assign n11598 = ~n11593 & n11597;
  assign n5782 = ~n11596 | n11598;
  assign n11600 = ~Ng5142 & n6143_1;
  assign n11601 = Pg35 & ~Ng5142;
  assign n11602 = ~Pg35 & Ng5138;
  assign n11603 = ~n11601 & ~n11602;
  assign n11604 = ~n6143_1 & n11603;
  assign n5787 = ~n11600 & ~n11604;
  assign n11606 = n5041 & n9551;
  assign n11607 = n5018 & n11606;
  assign n11608 = Pg35 & ~Ng5248;
  assign n11609 = ~n11606 & n11608;
  assign n11610 = ~Pg35 & ~Ng5232;
  assign n11611 = ~n11609 & ~n11610;
  assign n5792 = ~n11607 & n11611;
  assign n11613 = Ng2126 & n6950;
  assign n11614 = Pg35 & ~Ng2116;
  assign n11615 = ~Ng2122 & n11614;
  assign n11616 = Ng2122 & ~n11614;
  assign n11617 = ~n11615 & ~n11616;
  assign n11618 = ~n6950 & ~n11617;
  assign n5797 = n11613 | n11618;
  assign n11620 = ~Pg35 & Ng3689;
  assign n11621 = ~Ng3698 & n8918;
  assign n5802 = n11620 | n11621;
  assign n11623 = Ng5481 & n10635;
  assign n11624 = Ng5475 & ~n10635;
  assign n5807 = n11623 | n11624;
  assign n11626 = ~Ng1964 & ~n9572;
  assign n11627 = Pg35 & Ng1955;
  assign n11628 = Ng1959 & n11627;
  assign n11629 = ~Ng1959 & ~n11627;
  assign n11630 = ~n11628 & ~n11629;
  assign n11631 = n9572 & ~n11630;
  assign n5812_1 = ~n11626 & ~n11631;
  assign n11633 = ~Pg35 & Ng5092;
  assign n11634 = ~Ng5097 & ~n6785;
  assign n11635 = ~n11005 & ~n11634;
  assign n5817_1 = n11633 | n11635;
  assign n11637 = ~Pg35 & ~Ng3187;
  assign n11638 = n7522 & n8807;
  assign n11639 = n5018 & n11638;
  assign n11640 = Pg35 & ~Ng3215;
  assign n11641 = ~n11638 & n11640;
  assign n11642 = ~n11639 & ~n11641;
  assign n5822 = ~n11637 & n11642;
  assign n11644 = Pg35 & Ng4388;
  assign n11645 = Ng4430 & ~n11644;
  assign n11646 = ~Ng4430 & n11644;
  assign n11647 = ~n11645 & ~n11646;
  assign n11648 = Ng4434 & ~Ng4401;
  assign n11649 = ~Ng4434 & Ng4401;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = Pg35 & ~n11650;
  assign n5834 = ~n11647 | n11651;
  assign n11653 = ~Ng1768 & n8039;
  assign n11654 = Ng2779 & n8036;
  assign n11655 = ~Pg35 & Ng2767;
  assign n11656 = ~n11654 & ~n11655;
  assign n5839 = n11653 | ~n11656;
  assign n11658 = ~Pg35 & Ng4443;
  assign n11659 = Ng4438 & n6732;
  assign n11660 = ~n9041 & ~n11659;
  assign n5847_1 = n11658 | ~n11660;
  assign n11662 = Ng1720 & n7903;
  assign n11663 = Ng1714 & ~n7903;
  assign n5851 = n11662 | n11663;
  assign n11665 = ~Pg35 & Ng1361;
  assign n11666 = ~Ng1367 & ~n7250;
  assign n11667 = n7253 & ~n11666;
  assign n5856 = n11665 | n11667;
  assign n11669 = ~Pg35 & ~Ng4104;
  assign n11670 = Pg120 & ~Ng4146;
  assign n11671 = Pg124 & Ng4146;
  assign n11672 = Pg35 & ~n11671;
  assign n11673 = ~n11670 & n11672;
  assign n5865_1 = ~n11669 & ~n11673;
  assign n11675 = ~Ng2197 & n10680;
  assign n11676 = Pg35 & ~n11675;
  assign n11677 = Ng2161 & n11676;
  assign n11678 = ~Pg35 & Ng2165;
  assign n11679 = ~n6505 & ~n11678;
  assign n11680 = ~n11676 & ~n11679;
  assign n5870_1 = n11677 | n11680;
  assign n11682 = ~Pg35 & Ng370;
  assign n11683 = ~Ng358 & ~Ng376;
  assign n11684 = ~n5024 & ~n11683;
  assign n11685 = Pg35 & n11684;
  assign n5875_1 = n11682 | n11685;
  assign n11687 = Ng2361 & n6528;
  assign n11688 = Pg35 & n6531;
  assign n11689 = Ng2331 & ~n11688;
  assign n11690 = ~n6528 & n11689;
  assign n5880_1 = n11687 | n11690;
  assign n11692 = ~Pg35 & ~Ng2946;
  assign n11693 = Pg8786 & ~Ng4180;
  assign n11694 = ~Pg8784 & ~Pg8787;
  assign n11695 = ~Pg8783 & ~Pg8785;
  assign n11696 = ~Pg8789 & ~Pg11447;
  assign n11697 = ~Pg8788 & n11696;
  assign n11698 = n11695 & n11697;
  assign n11699 = n11694 & n11698;
  assign n11700 = ~Ng4180 & ~n11699;
  assign n11701 = ~Pg8786 & ~n11700;
  assign n11702 = Pg35 & ~n11701;
  assign n11703 = ~n11693 & n11702;
  assign n5885_1 = ~n11692 & ~n11703;
  assign n11705 = ~Pg35 & Ng577;
  assign n11706 = Ng582 & n5737;
  assign n11707 = ~n5751 & ~n11706;
  assign n11708 = ~n5752 & ~n11707;
  assign n5889 = n11705 | n11708;
  assign n11710 = Ng2028 & ~n11233;
  assign n11711 = Ng2051 & n11233;
  assign n11712 = ~n10975 & ~n11711;
  assign n5894_1 = n11710 | ~n11712;
  assign n11714 = Ng1193 & ~n7034;
  assign n11715 = Pg35 & ~n6574;
  assign n11716 = ~n11714 & n11715;
  assign n11717 = ~Pg35 & ~Ng1189;
  assign n5899 = ~n11716 & ~n11717;
  assign n11719 = Pg35 & ~n4667;
  assign n11720 = ~n7142 & ~n11719;
  assign n11721 = Ng2327 & ~n11720;
  assign n11722 = ~Pg35 & Ng2307;
  assign n11723 = Pg35 & ~n8751;
  assign n11724 = ~n11722 & ~n11723;
  assign n11725 = n11720 & ~n11724;
  assign n5904 = n11721 | n11725;
  assign n11727 = ~Pg35 & Ng936;
  assign n11728 = Ng907 & n6167;
  assign n11729 = ~n6161_1 & ~n11728;
  assign n11730 = ~n6162 & ~n11729;
  assign n5909 = n11727 | n11730;
  assign n5914 = Pg35 & Ng947;
  assign n11733 = ~Ng1834 & n10001;
  assign n11734 = ~Pg35 & Ng1830;
  assign n11735 = ~n9699 & ~n11734;
  assign n11736 = ~n10001 & n11735;
  assign n5919_1 = ~n11733 & ~n11736;
  assign n11738 = n4705 & n5201;
  assign n11739 = Pg35 & ~n11738;
  assign n11740 = Ng3594 & n11739;
  assign n11741 = ~Pg35 & Ng3578;
  assign n11742 = ~n5083 & ~n11741;
  assign n11743 = ~n11739 & ~n11742;
  assign n5924_1 = n11740 | n11743;
  assign n11745 = ~Ng2932 & ~Ng2999;
  assign n5929 = Pg35 & ~n11745;
  assign n11747 = ~Pg35 & Ng2295;
  assign n11748 = Ng2331 & ~Ng2361;
  assign n11749 = ~n4978 & n11748;
  assign n11750 = Pg35 & ~n11749;
  assign n11751 = ~n11747 & ~n11750;
  assign n11752 = ~n4986 & n11751;
  assign n11753 = ~Ng2303 & n11750;
  assign n5934 = ~n11752 & ~n11753;
  assign n11755 = Ng699 & n5151;
  assign n11756 = ~Pg35 & Ng681;
  assign n11757 = ~n10767 & ~n11756;
  assign n5942 = n11755 | ~n11757;
  assign n11759 = Ng822 & n9235;
  assign n11760 = ~Ng723 & n11759;
  assign n11761 = Pg35 & ~n11760;
  assign n11762 = Ng827 & ~n11761;
  assign n11763 = ~Ng827 & n7045;
  assign n11764 = ~n7046 & ~n11763;
  assign n11765 = Ng723 & ~n11764;
  assign n5947_1 = n11762 | n11765;
  assign n11767 = Ng5703 & n6894;
  assign n11768 = ~Pg35 & Ng5698;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = n4531 & n6893;
  assign n11771 = n5933 & n11770;
  assign n11772 = n6904 & ~n11771;
  assign n11773 = ~Ng5703 & n11772;
  assign n5952_1 = ~n11769 | n11773;
  assign n11775 = ~Ng546 & Ng691;
  assign n11776 = Pg35 & n11775;
  assign n11777 = ~Pg35 & ~Ng538;
  assign n5957_1 = ~n11776 & ~n11777;
  assign n11779 = ~Pg35 & Ng2421;
  assign n11780 = ~Ng112 & ~n4571;
  assign n11781 = Ng112 & n4571;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = n4570 & n6955;
  assign n11784 = n11782 & n11783;
  assign n11785 = n5842 & n11784;
  assign n11786 = ~n11779 & ~n11785;
  assign n11787 = n4928 & n11783;
  assign n11788 = Ng2472 & ~n11787;
  assign n11789 = Pg35 & n11788;
  assign n5962_1 = ~n11786 | n11789;
  assign n11791 = n7328 & n9706;
  assign n11792 = n5083 & n11791;
  assign n11793 = ~Pg35 & Ng5937;
  assign n11794 = ~n11792 & ~n11793;
  assign n11795 = Pg35 & Ng5953;
  assign n11796 = ~n11791 & n11795;
  assign n5967 = ~n11794 | n11796;
  assign n11798 = Pg35 & Ng3338;
  assign n11799 = ~Pg35 & Ng3050;
  assign n5972 = n11798 | n11799;
  assign n11801 = ~Pg35 & Ng1821;
  assign n11802 = ~n5070 & ~n11801;
  assign n11803 = n8858 & n11802;
  assign n11804 = ~Ng1740 & ~n8858;
  assign n5976 = ~n11803 & ~n11804;
  assign n11806 = ~Pg35 & ~Ng3554;
  assign n11807 = n5034 & n5828;
  assign n11808 = ~n5018 & n11807;
  assign n11809 = Pg35 & ~Ng3550;
  assign n11810 = ~n11807 & ~n11809;
  assign n11811 = ~n11808 & ~n11810;
  assign n5981 = ~n11806 & ~n11811;
  assign n11813 = Ng3841 & n7019;
  assign n11814 = ~Ng3841 & ~n7019;
  assign n11815 = ~n11813 & ~n11814;
  assign n11816 = ~n5730 & ~n11815;
  assign n11817 = ~Ng3845 & n5730;
  assign n5986_1 = ~n11816 & ~n11817;
  assign n11819 = ~Pg35 & Ng2112;
  assign n11820 = ~n11614 & ~n11819;
  assign n11821 = n5664 & n11820;
  assign n11822 = ~Ng2116 & ~n5664;
  assign n5991 = ~n11821 & ~n11822;
  assign n11824 = Ng3167 & n7522;
  assign n11825 = Pg35 & ~n11824;
  assign n11826 = Ng3195 & n11825;
  assign n11827 = ~Pg35 & Ng3247;
  assign n11828 = ~n5083 & ~n11827;
  assign n11829 = ~n11825 & ~n11828;
  assign n5999_1 = n11826 | n11829;
  assign n11831 = Ng3869 & n7216;
  assign n11832 = Pg35 & ~n11831;
  assign n11833 = Ng3913 & n11832;
  assign n11834 = ~Pg35 & Ng3957;
  assign n11835 = ~n5083 & ~n11834;
  assign n11836 = ~n11832 & ~n11835;
  assign n6004_1 = n11833 | n11836;
  assign n11838 = n6677 & ~n9692;
  assign n11839 = ~Ng4581 & ~Ng4512;
  assign n11840 = ~n5182 & n11839;
  assign n11841 = Pg35 & ~n11840;
  assign n11842 = ~n11838 & n11841;
  assign n11843 = ~Pg35 & Ng4492;
  assign n6009 = n11842 | n11843;
  assign n11845 = Ng1682 & n5247;
  assign n11846 = Ng1687 & ~n5247;
  assign n6013_1 = n11845 | n11846;
  assign n11848 = Ng2681 & n11288;
  assign n11849 = Ng2675 & ~n11288;
  assign n6018 = n11848 | n11849;
  assign n11851 = Ng2527 & n7009;
  assign n11852 = Ng2533 & ~n7009;
  assign n6023_1 = n11851 | n11852;
  assign n11854 = ~Pg35 & ~Ng336;
  assign n11855 = ~Ng311 & Ng324;
  assign n11856 = n8268 & ~n11855;
  assign n6028 = ~n11854 & ~n11856;
  assign n11858 = Pg35 & Ng2697;
  assign n11859 = ~Pg35 & Ng2689;
  assign n6033_1 = n11858 | n11859;
  assign n11861 = ~Pg35 & Ng4382;
  assign n6038 = n5842 | n11861;
  assign n11863 = ~Pg35 & Ng6555;
  assign n11864 = n7556 & n7715;
  assign n6043_1 = n11863 | n11864;
  assign n11866 = ~Pg35 & Ng1129;
  assign n11867 = ~Ng1141 & ~n10181;
  assign n11868 = Ng1141 & n5813;
  assign n11869 = ~Ng956 & n10176;
  assign n11870 = Ng956 & ~n10176;
  assign n11871 = ~n11869 & ~n11870;
  assign n11872 = n8547 & ~n11871;
  assign n11873 = ~n11868 & ~n11872;
  assign n11874 = ~n11867 & ~n11873;
  assign n6048_1 = n11866 | n11874;
  assign n11876 = Pg35 & Ng496;
  assign n11877 = ~Pg35 & Ng1554;
  assign n6053 = n11876 | n11877;
  assign n11879 = Ng2413 & n8160;
  assign n11880 = Ng2407 & ~n8160;
  assign n6057_1 = n11879 | n11880;
  assign n11882 = Ng1706 & n7905;
  assign n11883 = ~Ng1706 & ~n7905;
  assign n11884 = ~n11882 & ~n11883;
  assign n11885 = n5247 & n11884;
  assign n11886 = Ng1710 & ~n5247;
  assign n6062_1 = n11885 | n11886;
  assign n11888 = ~Pg35 & Ng6523;
  assign n11889 = ~Ng6527 & ~n7839;
  assign n11890 = ~n7314 & ~n7840;
  assign n11891 = ~n11889 & ~n11890;
  assign n6067 = n11888 | n11891;
  assign n11893 = n5396 & n6081;
  assign n11894 = n5018 & n11893;
  assign n11895 = ~Pg35 & ~Ng3239;
  assign n11896 = ~n11894 & ~n11895;
  assign n11897 = Pg35 & ~n11893;
  assign n11898 = ~Ng3255 & n11897;
  assign n6072_1 = n11896 & ~n11898;
  assign n11900 = Ng1677 & ~n8570;
  assign n11901 = Ng1691 & ~n8573;
  assign n11902 = ~n11900 & n11901;
  assign n11903 = n11900 & ~n11901;
  assign n6077_1 = n11902 | n11903;
  assign n11905 = Pg35 & Ng2936;
  assign n11906 = ~Pg35 & Ng2922;
  assign n6082_1 = n11905 | n11906;
  assign n11908 = ~Pg35 & Ng5703;
  assign n11909 = Ng5644 & n6894;
  assign n11910 = ~n4549 & n6904;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n10871 & ~n11771;
  assign n11913 = ~n11911 & n11912;
  assign n6087 = n11908 | n11913;
  assign n11915 = Ng5148 & n11601;
  assign n11916 = ~Ng5148 & ~n11601;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = ~n10211 & ~n11917;
  assign n11919 = ~Ng5152 & n10211;
  assign n6092_1 = ~n11918 & ~n11919;
  assign n11921 = Pg35 & n6123;
  assign n6097_1 = Ng5348 & ~n11921;
  assign n11923 = Ng2779 & ~n4928;
  assign n11924 = ~n4932 & n7075;
  assign n11925 = ~n11923 & n11924;
  assign n11926 = Ng2775 & ~n7075;
  assign n11927 = Pg35 & ~n11926;
  assign n11928 = ~n11925 & n11927;
  assign n11929 = ~Pg35 & ~Ng2783;
  assign n6105_1 = ~n11928 & ~n11929;
  assign n11931 = Pg35 & Ng2922;
  assign n11932 = ~Pg35 & Ng2912;
  assign n6110 = n11931 | n11932;
  assign n11934 = ~Ng1105 & n10176;
  assign n11935 = Ng1105 & ~n10176;
  assign n11936 = ~n11934 & ~n11935;
  assign n11937 = n7132 & n11936;
  assign n11938 = n7132 & n10181;
  assign n11939 = ~Ng1111 & ~n11938;
  assign n11940 = Pg35 & ~n11939;
  assign n11941 = ~n11937 & n11940;
  assign n11942 = ~Pg35 & Ng1135;
  assign n6115_1 = n11941 | n11942;
  assign n11944 = n5078 & n9706;
  assign n11945 = n5083 & n11944;
  assign n11946 = ~Pg35 & Ng5897;
  assign n11947 = ~n11945 & ~n11946;
  assign n11948 = Pg35 & Ng5893;
  assign n11949 = ~n11944 & n11948;
  assign n6120_1 = ~n11947 | n11949;
  assign n11951 = ~Pg35 & ~Ng6593;
  assign n11952 = n7557 & n8582;
  assign n11953 = Pg35 & ~Ng6617;
  assign n11954 = ~n11952 & n11953;
  assign n11955 = n5018 & n11952;
  assign n11956 = ~n11954 & ~n11955;
  assign n6128_1 = ~n11951 & n11956;
  assign n11958 = ~Pg35 & Ng2066;
  assign n11959 = Ng2051 & n10971;
  assign n11960 = ~n11958 & ~n11959;
  assign n11961 = Ng2060 & n11233;
  assign n11962 = ~n10975 & ~n11961;
  assign n6133_1 = ~n11960 | ~n11962;
  assign n11964 = ~n5182 & n5406;
  assign n11965 = Ng4504 & ~n5406;
  assign n11966 = ~n6976 & ~n11965;
  assign n6138 = n11964 | ~n11966;
  assign n11968 = n4726 & n5373;
  assign n11969 = n5083 & n11968;
  assign n11970 = ~Pg35 & Ng5583;
  assign n11971 = ~n11969 & ~n11970;
  assign n11972 = Pg35 & Ng5599;
  assign n11973 = ~n11968 & n11972;
  assign n6143 = ~n11971 | n11973;
  assign n11975 = ~Ng3451 & Pg8279;
  assign n11976 = ~Ng3401 & ~n11975;
  assign n11977 = Pg35 & ~Pg8342;
  assign n11978 = ~n11976 & n11977;
  assign n11979 = ~Pg35 & Ng3451;
  assign n6148 = n11978 | n11979;
  assign n11981 = Ng4633 & n4534;
  assign n11982 = n5180 & n5560;
  assign n11983 = n11981 & n11982;
  assign n6153 = Pg35 & ~n11983;
  assign n11985 = Pg35 & \[4433] ;
  assign n11986 = ~Pg35 & Ng37;
  assign n6161 = n11985 | n11986;
  assign n11988 = Ng3129 & n9124;
  assign n11989 = Pg35 & ~Ng3119;
  assign n11990 = ~Ng3125 & n11989;
  assign n11991 = n9123 & n11990;
  assign n11992 = ~n11988 & ~n11991;
  assign n11993 = Ng3125 & ~n11989;
  assign n11994 = ~n9124 & n11993;
  assign n6166 = ~n11992 | n11994;
  assign n11996 = ~Pg35 & Ng5164;
  assign n11997 = ~n5042_1 & ~n9551;
  assign n11998 = n5598 & ~n11997;
  assign n6175 = n11996 | n11998;
  assign n6180 = ~Pg35 & Ng4392;
  assign n12001 = ~Ng5821 & n5050;
  assign n12002 = ~Pg35 & Ng5817;
  assign n12003 = ~n7487 & ~n12002;
  assign n12004 = ~n5050 & n12003;
  assign n6184 = ~n12001 & ~n12004;
  assign n12006 = n5849 & n6385;
  assign n12007 = Pg35 & ~n12006;
  assign n12008 = ~Pg35 & ~Ng6283;
  assign n12009 = ~n5018 & ~n12008;
  assign n12010 = ~n12007 & ~n12009;
  assign n12011 = ~Ng6299 & n12007;
  assign n6189 = ~n12010 & ~n12011;
  assign n12013 = n6948 & n10977;
  assign n12014 = Ng2008 & n12013;
  assign n12015 = Ng2079 & n11233;
  assign n12016 = ~Pg35 & Ng2060;
  assign n12017 = Ng2024 & n4639;
  assign n12018 = Ng2016 & ~Ng2060;
  assign n12019 = ~Ng2028 & n12018;
  assign n12020 = Ng2004 & n10395;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = Ng2020 & Ng2028;
  assign n12023 = ~Ng2051 & n12022;
  assign n12024 = Ng2012 & n11096;
  assign n12025 = ~n12023 & ~n12024;
  assign n12026 = n12021 & n12025;
  assign n12027 = ~n12017 & n12026;
  assign n12028 = n10971 & ~n12027;
  assign n12029 = ~n12016 & ~n12028;
  assign n12030 = ~n12015 & n12029;
  assign n6197 = n12014 | ~n12030;
  assign n12032 = ~Ng4698 & ~n4616;
  assign n12033 = ~n5669 & ~n12032;
  assign n12034 = n6519 & ~n12033;
  assign n12035 = n4616 & ~n6513_1;
  assign n12036 = Pg35 & ~n12035;
  assign n12037 = ~Ng4704 & ~n12036;
  assign n6202 = ~n12034 & ~n12037;
  assign n12039 = ~Pg35 & Ng3698;
  assign n12040 = Ng3703 & n8292;
  assign n12041 = ~n12039 & ~n12040;
  assign n12042 = n5484 & ~n8301;
  assign n12043 = ~Ng3703 & n12042;
  assign n6207_1 = ~n12041 | n12043;
  assign n12045 = ~Pg35 & Ng1564;
  assign n12046 = ~Ng1559 & ~n7548;
  assign n12047 = ~n11508 & ~n12046;
  assign n12048 = n11510 & n12047;
  assign n6212 = n12045 | n12048;
  assign n12050 = ~Pg35 & ~Ng939;
  assign n12051 = ~Ng943 & n9487;
  assign n6217 = ~n12050 & ~n12051;
  assign n12053 = ~Pg35 & Ng417;
  assign n12054 = Ng411 & n5151;
  assign n12055 = n6741 & n9287;
  assign n12056 = ~n12054 & ~n12055;
  assign n6222 = n12053 | ~n12056;
  assign n12058 = n7736 & n9940;
  assign n12059 = n5083 & n12058;
  assign n12060 = ~Pg35 & Ng3937;
  assign n12061 = ~n12059 & ~n12060;
  assign n12062 = Pg35 & Ng3953;
  assign n12063 = ~n12058 & n12062;
  assign n6231 = ~n12061 | n12063;
  assign n12065 = Pg35 & Ng2704;
  assign n12066 = ~Pg35 & Ng2697;
  assign n6236 = n12065 | n12066;
  assign n12068 = ~Pg35 & Ng6031;
  assign n12069 = ~Ng6035 & ~n8326;
  assign n12070 = n8328 & ~n12069;
  assign n6241 = n12068 | n12070;
  assign n12072 = ~Pg35 & Ng1484;
  assign n12073 = Ng1484 & n6265;
  assign n12074 = n7677 & n12073;
  assign n12075 = Ng1300 & n12074;
  assign n12076 = Pg35 & Ng1300;
  assign n12077 = ~n12074 & ~n12076;
  assign n12078 = ~n12075 & ~n12077;
  assign n6246 = n12072 | n12078;
  assign n12080 = ~Pg35 & Ng4064;
  assign n12081 = ~n9024 & ~n11481;
  assign n12082 = n7718 & ~n12081;
  assign n6251_1 = n12080 | n12082;
  assign n12084 = n7616 & n10319;
  assign n12085 = Pg35 & ~n12084;
  assign n12086 = Ng5200 & n12085;
  assign n12087 = ~Pg35 & Ng5204;
  assign n12088 = ~n5083 & ~n12087;
  assign n12089 = ~n12085 & ~n12088;
  assign n6256_1 = n12086 | n12089;
  assign n12091 = Pg35 & Ng4843;
  assign n12092 = ~Ng4878 & ~n12091;
  assign n12093 = Ng4878 & n12091;
  assign n12094 = ~n12092 & ~n12093;
  assign n6261_1 = ~n5818 & n12094;
  assign n12096 = ~Pg35 & Ng5041;
  assign n12097 = Ng5046 & ~n4911;
  assign n12098 = ~n4904 & ~n12097;
  assign n12099 = ~n4912 & n12098;
  assign n12100 = n7590 & ~n12099;
  assign n12101 = ~n4905_1 & n12100;
  assign n6266 = n12096 | n12101;
  assign n12103 = Ng2236 & ~n5259;
  assign n12104 = Ng2250 & ~n7160;
  assign n12105 = ~n12103 & n12104;
  assign n12106 = n12103 & ~n12104;
  assign n6271 = n12105 | n12106;
  assign n12108 = ~Pg35 & ~Ng316;
  assign n6276 = ~n8269 & ~n12108;
  assign n12110 = Ng4546 & ~n5406;
  assign n12111 = ~n5409 & ~n12110;
  assign n6280 = n7572 | ~n12111;
  assign n12113 = ~Ng2476 & n6154;
  assign n12114 = ~Ng2485 & n12113;
  assign n12115 = ~n5008_1 & n10535;
  assign n12116 = ~Pg35 & Ng2461;
  assign n12117 = ~n12115 & ~n12116;
  assign n12118 = ~n6153_1 & n12117;
  assign n6285 = n12114 | ~n12118;
  assign n12120 = Ng5841 & n5050;
  assign n12121 = Ng5835 & ~n5050;
  assign n6290_1 = n12120 | n12121;
  assign n12123 = Pg35 & Ng2912;
  assign n12124 = ~Pg35 & Ng2907;
  assign n6298 = n12123 | n12124;
  assign n12126 = n4928 & n7145;
  assign n12127 = Ng2357 & ~n12126;
  assign n12128 = Pg35 & n12127;
  assign n12129 = Ng110 & n7696;
  assign n12130 = ~Ng110 & ~n7696;
  assign n12131 = ~n12129 & ~n12130;
  assign n12132 = n5842 & n12131;
  assign n12133 = n7145 & n12132;
  assign n12134 = ~Pg35 & Ng2342;
  assign n12135 = ~n12133 & ~n12134;
  assign n6303 = n12128 | ~n12135;
  assign n12137 = ~Pg35 & Ng146;
  assign n12138 = Ng164 & n7270;
  assign n12139 = ~n7265 & ~n12138;
  assign n12140 = ~n7266 & ~n12139;
  assign n6311 = n12137 | n12140;
  assign n12142 = Pg35 & Ng4253;
  assign n12143 = ~Pg35 & Ng4300;
  assign n6316 = n12142 | n12143;
  assign n12145 = ~Ng5022 & ~Ng5062;
  assign n12146 = n7829 & ~n12145;
  assign n12147 = ~Pg35 & Ng5022;
  assign n12148 = Ng5016 & n12145;
  assign n12149 = Pg35 & n12148;
  assign n12150 = ~n12147 & ~n12149;
  assign n6321 = n12146 | ~n12150;
  assign n12152 = ~Ng3119 & n5955;
  assign n12153 = ~Pg35 & Ng3115;
  assign n12154 = ~n11989 & ~n12153;
  assign n12155 = ~n5955 & n12154;
  assign n6326 = ~n12152 & ~n12155;
  assign n12157 = Ng1312 & ~n10748;
  assign n12158 = ~n7242 & ~n10750;
  assign n12159 = ~n5506 & ~n12158;
  assign n12160 = n6547_1 & ~n12159;
  assign n6331 = n12157 | n12160;
  assign n12162 = Ng1624 & ~n8570;
  assign n12163 = Ng1648 & n8570;
  assign n12164 = ~n9632 & ~n12163;
  assign n6336 = n12162 | ~n12164;
  assign n12166 = Ng4581 & ~\[4437] ;
  assign n12167 = n5182 & n12166;
  assign n12168 = Pg35 & ~n11839;
  assign n12169 = ~n12167 & n12168;
  assign n12170 = ~Pg35 & Ng4515;
  assign n6341_1 = n12169 | n12170;
  assign n12172 = ~Pg35 & Ng5120;
  assign n12173 = ~n6062 & n6064;
  assign n12174 = n6066 & ~n12173;
  assign n12175 = Pg35 & ~n12174;
  assign n12176 = Ng5115 & n12175;
  assign n12177 = ~Ng5115 & n6068;
  assign n12178 = ~n12176 & ~n12177;
  assign n6345 = n12172 | ~n12178;
  assign n12180 = Ng3352 & n9130;
  assign n12181 = ~Pg35 & Ng3347;
  assign n12182 = ~n12180 & ~n12181;
  assign n12183 = ~n7882 & n9195;
  assign n12184 = ~Ng3352 & n12183;
  assign n6350 = ~n12182 | n12184;
  assign n12186 = Ng6657 & n7313;
  assign n12187 = ~Pg35 & Ng6653;
  assign n12188 = ~n5083 & ~n12187;
  assign n12189 = ~n7313 & ~n12188;
  assign n6355 = n12186 | n12189;
  assign n12191 = Ng4549 & ~n5406;
  assign n12192 = ~n6666_1 & ~n12191;
  assign n6360 = n11964 | ~n12192;
  assign n12194 = n5767 & n9940;
  assign n12195 = Pg35 & ~n12194;
  assign n12196 = Ng3893 & n12195;
  assign n12197 = ~Pg35 & Ng3897;
  assign n12198 = ~n5083 & ~n12197;
  assign n12199 = ~n12195 & ~n12198;
  assign n6365 = n12196 | n12199;
  assign n12201 = Ng3167 & n6081;
  assign n12202 = Pg35 & ~n12201;
  assign n12203 = Ng3211 & n12202;
  assign n12204 = ~Pg35 & Ng3255;
  assign n12205 = ~n5083 & ~n12204;
  assign n12206 = ~n12202 & ~n12205;
  assign n6370 = n12203 | n12206;
  assign n12208 = n5373 & n6172;
  assign n12209 = n5083 & n12208;
  assign n12210 = ~Pg35 & Ng5579;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = Pg35 & Ng5595;
  assign n12213 = ~n12208 & n12212;
  assign n6381 = ~n12211 | n12213;
  assign n12215 = Ng3614 & n5213;
  assign n12216 = ~Pg35 & Ng3610;
  assign n12217 = ~n5083 & ~n12216;
  assign n12218 = ~n5213 & ~n12217;
  assign n6386_1 = n12215 | n12218;
  assign n12220 = Pg35 & Ng2894;
  assign n12221 = ~Pg35 & Ng2860;
  assign n6391 = n12220 | n12221;
  assign n12223 = Ng3125 & n9124;
  assign n12224 = Ng3119 & ~n9124;
  assign n6396 = n12223 | n12224;
  assign n12226 = ~Ng3821 & n5730;
  assign n12227 = ~Pg35 & Ng3817;
  assign n12228 = ~n7870 & ~n12227;
  assign n12229 = ~n5730 & n12228;
  assign n6404 = ~n12226 & ~n12229;
  assign n12231 = ~Pg35 & Ng4057;
  assign n12232 = Pg35 & Ng4141;
  assign n12233 = ~n6200 & ~n12232;
  assign n12234 = Ng2841 & ~n12233;
  assign n12235 = ~n6201 & n12234;
  assign n6409 = n12231 | n12235;
  assign n12237 = Ng4552 & ~n5406;
  assign n12238 = ~n5409 & ~n12237;
  assign n6414 = n11964 | ~n12238;
  assign n12240 = Ng5272 & n10211;
  assign n12241 = ~Pg35 & Ng5268;
  assign n12242 = ~n5083 & ~n12241;
  assign n12243 = ~n10211 & ~n12242;
  assign n6418 = n12240 | n12243;
  assign n12245 = ~Pg35 & Ng2729;
  assign n12246 = ~n6197_1 & ~n12245;
  assign n12247 = Pg35 & Ng2735;
  assign n12248 = ~n7798 & ~n12247;
  assign n12249 = ~n7800 & ~n12248;
  assign n6423 = ~n12246 | n12249;
  assign n12251 = Ng728 & n6095;
  assign n12252 = Ng661 & ~n6095;
  assign n6428 = n12251 | n12252;
  assign n12254 = n5849 & n7336;
  assign n12255 = Pg35 & ~n12254;
  assign n12256 = Ng6295 & n12255;
  assign n12257 = ~Pg35 & Ng6279;
  assign n12258 = ~n5083 & ~n12257;
  assign n12259 = ~n12255 & ~n12258;
  assign n6433 = n12256 | n12259;
  assign n12261 = ~Ng2661 & n11288;
  assign n12262 = ~Pg35 & Ng2657;
  assign n12263 = ~n10983 & ~n12262;
  assign n12264 = ~n11288 & n12263;
  assign n6438 = ~n12261 & ~n12264;
  assign n12266 = Ng1988 & n5300;
  assign n12267 = Ng1982 & ~n5300;
  assign n6443 = n12266 | n12267;
  assign n12269 = ~Ng5128 & n10211;
  assign n12270 = ~Pg35 & Ng5124;
  assign n12271 = ~n7958 & ~n12270;
  assign n12272 = ~n10211 & n12271;
  assign n6448 = ~n12269 & ~n12272;
  assign n12274 = Pg35 & Ng1548;
  assign n12275 = ~Ng1430 & n12274;
  assign n12276 = Ng1430 & ~n12274;
  assign n6453 = n12275 | n12276;
  assign n12278 = ~Ng3106 & n9197;
  assign n12279 = Pg35 & Ng3106;
  assign n12280 = n9122 & ~n9193;
  assign n12281 = n7880 & ~n9194;
  assign n12282 = ~n12280 & n12281;
  assign n12283 = n12279 & ~n12282;
  assign n12284 = ~Pg35 & Ng3111;
  assign n12285 = ~n12283 & ~n12284;
  assign n6458 = n12278 | ~n12285;
  assign n12287 = ~Pg35 & Ng4653;
  assign n12288 = Ng4659 & n7978;
  assign n12289 = n4617 & ~n5548;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n4618_1 & ~n12290;
  assign n6463 = n12287 | n12291;
  assign n12293 = ~Pg35 & Ng4349;
  assign n12294 = ~Ng4358 & ~n5562;
  assign n12295 = ~n10249 & ~n12294;
  assign n12296 = ~n5309 & ~n5563;
  assign n12297 = n12295 & n12296;
  assign n6468 = n12293 | n12297;
  assign n12299 = ~Pg35 & Ng1798;
  assign n12300 = Ng1783 & n11387;
  assign n12301 = ~n12299 & ~n12300;
  assign n12302 = Ng1792 & n8434;
  assign n12303 = ~n8433 & ~n12302;
  assign n6473 = ~n12301 | ~n12303;
  assign n12305 = ~Pg35 & Ng2070;
  assign n12306 = ~Ng2084 & n5660;
  assign n12307 = ~Ng1246 & ~n5657;
  assign n12308 = ~n6910 & ~n12307;
  assign n12309 = Ng2084 & ~n5662;
  assign n12310 = n12308 & n12309;
  assign n12311 = ~n12308 & ~n12309;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = ~n5660 & n12312;
  assign n12314 = Pg35 & ~n12313;
  assign n12315 = ~n12306 & n12314;
  assign n6478 = n12305 | n12315;
  assign n12317 = ~Pg35 & ~Ng3179;
  assign n12318 = n7522 & n11519;
  assign n12319 = ~n5018 & n12318;
  assign n12320 = Pg35 & ~Ng3187;
  assign n12321 = ~n12318 & ~n12320;
  assign n12322 = ~n12319 & ~n12321;
  assign n6483 = ~n12317 & ~n12322;
  assign n12324 = ~Ng4311 & ~n5563;
  assign n6488 = n11047 & ~n12324;
  assign n12326 = ~Pg35 & Ng2571;
  assign n12327 = n4568 & ~n5533;
  assign n12328 = Pg35 & ~n12327;
  assign n12329 = ~n5543 & ~n12328;
  assign n12330 = ~n12326 & n12329;
  assign n12331 = ~Ng2583 & n12328;
  assign n6493 = ~n12330 & ~n12331;
  assign n6498 = ~Pg35 & Ng2975;
  assign n12334 = ~Ng1135 & n10176;
  assign n12335 = Ng1135 & ~n10176;
  assign n12336 = ~n12334 & ~n12335;
  assign n12337 = n6105 & n12336;
  assign n12338 = n6105 & n10181;
  assign n12339 = ~Ng1094 & ~n12338;
  assign n12340 = Pg35 & ~n12339;
  assign n12341 = ~n12337 & n12340;
  assign n12342 = ~Pg35 & Ng1099;
  assign n6503 = n12341 | n12342;
  assign n12344 = Ng3841 & n5730;
  assign n12345 = Ng3835 & ~n5730;
  assign n6508 = n12344 | n12345;
  assign n12347 = Pg35 & Pg8839;
  assign n12348 = ~Ng4281 & ~n12347;
  assign n12349 = Pg8839 & n9764;
  assign n6513 = ~n12348 & ~n12349;
  assign n12351 = n6658 & n11519;
  assign n12352 = Pg35 & ~n12351;
  assign n12353 = Ng3191 & n12352;
  assign n12354 = ~Pg35 & Ng3195;
  assign n12355 = ~n5083 & ~n12354;
  assign n12356 = ~n12352 & ~n12355;
  assign n6518 = n12353 | n12356;
  assign n12358 = Pg35 & Ng4239;
  assign n12359 = ~Pg35 & ~Ng4273;
  assign n6523 = ~n12358 & ~n12359;
  assign n12361 = Ng703 & ~Ng714;
  assign n12362 = n5351 & ~n12361;
  assign n12363 = Ng691 & ~n12362;
  assign n12364 = n10094 & ~n12363;
  assign n12365 = ~Pg35 & ~\[4435] ;
  assign n6532 = ~n12364 & ~n12365;
  assign n12367 = ~Ng534 & n8264;
  assign n12368 = ~Pg35 & ~Ng542;
  assign n6537 = ~n12367 & ~n12368;
  assign n12370 = Ng376 & ~n6980;
  assign n12371 = ~n6739 & ~n12370;
  assign n6542 = ~n6740 & ~n12371;
  assign n12373 = ~Ng2040 & n8013;
  assign n12374 = Pg35 & ~n12373;
  assign n12375 = Ng2004 & n12374;
  assign n12376 = ~Pg35 & Ng2008;
  assign n12377 = ~n6912 & ~n12376;
  assign n12378 = ~n12374 & ~n12377;
  assign n6547 = n12375 | n12378;
  assign n12380 = ~Ng2527 & n5010;
  assign n12381 = ~Pg35 & Ng2523;
  assign n12382 = ~n8120 & ~n12381;
  assign n12383 = ~n5010 & n12382;
  assign n6552 = ~n12380 & ~n12383;
  assign n12385 = Pg35 & Pg10306;
  assign n12386 = ~Ng4534 & n12385;
  assign n12387 = Ng4534 & ~n12385;
  assign n6561 = n12386 | n12387;
  assign n12389 = Ng5148 & n10211;
  assign n12390 = Ng5142 & ~n10211;
  assign n6566 = n12389 | n12390;
  assign n12392 = ~Ng4459 & Ng4473;
  assign n12393 = Ng4507 & ~n12392;
  assign n12394 = Pg113 & n12392;
  assign n12395 = Pg35 & ~n12394;
  assign n6571 = n12393 | ~n12395;
  assign n12397 = ~Pg35 & \[4415] ;
  assign n12398 = ~Ng5352 & n6124;
  assign n6576 = n12397 | n12398;
  assign n12400 = n6081 & n8807;
  assign n12401 = n5083 & n12400;
  assign n12402 = ~Pg35 & Ng3199;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = Pg35 & Ng3223;
  assign n12405 = ~n12400 & n12404;
  assign n6581 = ~n12403 | n12405;
  assign n12407 = Pg35 & Ng2970;
  assign n12408 = ~Pg35 & Ng2960;
  assign n6586 = n12407 | n12408;
  assign n12410 = Pg35 & n8652;
  assign n6591 = Ng5694 & ~n12410;
  assign n12412 = n6412 & n10319;
  assign n12413 = n5018 & n12412;
  assign n12414 = ~Pg35 & ~Ng5244;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416 = Pg35 & ~n12412;
  assign n12417 = ~Ng5260 & n12416;
  assign n6596 = n12415 & ~n12417;
  assign n12419 = ~Pg35 & Ng1526;
  assign n12420 = Pg7946 & ~Ng1339;
  assign n12421 = ~Pg7946 & ~Ng1521;
  assign n12422 = Pg35 & ~n12421;
  assign n12423 = ~n12420 & n12422;
  assign n6601 = n12419 | n12423;
  assign n12425 = ~Ng3522 & ~n5204;
  assign n12426 = Pg35 & ~n12425;
  assign n12427 = Ng3518 & ~n12426;
  assign n12428 = Ng3522 & n5950;
  assign n6606 = n12427 | n12428;
  assign n12430 = Pg35 & Ng3111;
  assign n12431 = Ng3106 & n12430;
  assign n12432 = ~Ng3106 & ~n12430;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~n9124 & ~n12433;
  assign n12435 = ~Ng3115 & n9124;
  assign n6611 = ~n12434 & ~n12435;
  assign n12437 = n5396 & n6658;
  assign n12438 = n5018 & n12437;
  assign n12439 = ~Pg35 & ~Ng3235;
  assign n12440 = ~n12438 & ~n12439;
  assign n12441 = Pg35 & ~n12437;
  assign n12442 = ~Ng3251 & n12441;
  assign n6616 = n12440 & ~n12442;
  assign n12444 = ~Pg35 & Ng4455;
  assign n6621 = ~n10457 | n12444;
  assign n12446 = ~Pg35 & Ng4621;
  assign n12447 = ~Ng4628 & ~n8953;
  assign n12448 = ~n8957 & ~n12447;
  assign n6625 = n12446 | n12448;
  assign n12450 = ~Ng1996 & n5660;
  assign n12451 = ~Ng2070 & ~n8816;
  assign n12452 = n8946 & n12451;
  assign n12453 = ~n5661 & ~n12452;
  assign n6630 = ~n12450 & ~n12453;
  assign n12455 = Pg35 & Ng3689;
  assign n12456 = ~Pg35 & Ng3401;
  assign n6635 = n12455 | n12456;
  assign n12458 = Pg35 & Ng4521;
  assign n12459 = Ng4515 & n12458;
  assign n12460 = ~Pg35 & ~Ng4527;
  assign n12461 = ~n12458 & ~n12460;
  assign n12462 = ~n9696 & n12461;
  assign n6639 = n12459 | n12462;
  assign n12464 = ~Ng4242 & ~Ng4300;
  assign n12465 = Pg35 & n12464;
  assign n12466 = ~Pg35 & ~Ng4297;
  assign n6647 = ~n12465 & ~n12466;
  assign n12468 = Ng1720 & n5242;
  assign n12469 = ~Ng1720 & ~n5242;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = ~n7903 & ~n12470;
  assign n12472 = ~Ng1724 & n7903;
  assign n6652 = ~n12471 & ~n12472;
  assign n12474 = Ng1379 & ~n7256;
  assign n12475 = ~Ng1379 & n7246;
  assign n12476 = Pg35 & ~n12475;
  assign n12477 = Ng1373 & ~n7253;
  assign n12478 = ~n12476 & n12477;
  assign n6657 = n12474 | n12478;
  assign n12480 = ~Pg13926 & ~Pg16744;
  assign n12481 = ~n5282 & ~n12480;
  assign n12482 = Pg35 & ~Pg16656;
  assign n12483 = ~Pg14451 & ~Pg16627;
  assign n12484 = n12482 & n12483;
  assign n6662 = ~n12481 & n12484;
  assign n12486 = ~Pg35 & Ng1870;
  assign n12487 = Ng1906 & ~n4950;
  assign n12488 = ~Ng1936 & n12487;
  assign n12489 = n4960 & n12488;
  assign n12490 = Pg35 & Ng1878;
  assign n12491 = ~n12488 & n12490;
  assign n12492 = ~n12489 & ~n12491;
  assign n6666 = n12486 | ~n12492;
  assign n12494 = Ng5619 & n7205;
  assign n12495 = ~Pg35 & Ng5615;
  assign n12496 = ~n5083 & ~n12495;
  assign n12497 = ~n7205 & ~n12496;
  assign n6671 = n12494 | n12497;
  assign Pg34597 = 1'b0;
  assign Pg34240 = 1'b0;
  assign Pg34239 = 1'b0;
  assign Pg34238 = 1'b0;
  assign Pg34237 = 1'b0;
  assign Pg34236 = 1'b0;
  assign Pg34235 = 1'b0;
  assign Pg34234 = 1'b0;
  assign Pg34233 = 1'b0;
  assign Pg34232 = 1'b0;
  assign Pg33950 = 1'b0;
  assign Pg33949 = 1'b0;
  assign Pg33948 = 1'b0;
  assign Pg33947 = 1'b0;
  assign Pg33946 = 1'b0;
  assign Pg33945 = 1'b0;
  assign Pg32454 = 1'b0;
  assign Pg32429 = 1'b0;
  assign Pg25590 = 1'b0;
  assign Pg25589 = 1'b0;
  assign Pg25588 = 1'b0;
  assign Pg25587 = 1'b0;
  assign Pg25586 = 1'b0;
  assign Pg25585 = 1'b0;
  assign Pg25584 = 1'b0;
  assign Pg25583 = 1'b0;
  assign Pg25582 = 1'b0;
  assign Pg24151 = 1'b0;
  assign Pg30331 = ~Ng2831;
  assign Pg30330 = ~Ng2834;
  assign Pg30329 = ~\[4426] ;
  assign Pg30327 = ~Ng37;
  assign Pg12833 = ~Pg5;
  assign Pg34839 = Pg34956;
  assign Pg33894 = Pg34788;
  assign Pg31861 = \[4415] ;
  assign Pg31665 = Pg34437;
  assign Pg31656 = Pg34436;
  assign Pg31521 = Pg34435;
  assign Pg30332 = \[4421] ;
  assign Pg29221 = \[4426] ;
  assign Pg29220 = \[4427] ;
  assign Pg29219 = \[4428] ;
  assign Pg29218 = \[4507] ;
  assign Pg29217 = \[4430] ;
  assign Pg29216 = \[4431] ;
  assign Pg29215 = \[4432] ;
  assign Pg29214 = \[4433] ;
  assign Pg29213 = \[4434] ;
  assign Pg29212 = \[4435] ;
  assign Pg29211 = \[4436] ;
  assign Pg29210 = \[4437] ;
  assign Pg28753 = Pg33959;
  assign Pg27831 = Pg33533;
  assign Pg26801 = Pg32975;
  assign Pg25259 = Pg31862;
  assign Pg25219 = \[4415] ;
  assign Pg25167 = Pg31863;
  assign Pg25114 = Pg31860;
  assign Pg24185 = Pg44;
  assign Pg24184 = Pg135;
  assign Pg24183 = Pg134;
  assign Pg24182 = Pg127;
  assign Pg24181 = Pg126;
  assign Pg24180 = Pg125;
  assign Pg24179 = Pg124;
  assign Pg24178 = Pg120;
  assign Pg24177 = Pg116;
  assign Pg24176 = Pg115;
  assign Pg24175 = Pg114;
  assign Pg24174 = Pg113;
  assign Pg24173 = Pg100;
  assign Pg24172 = Pg99;
  assign Pg24171 = Pg92;
  assign Pg24170 = Pg91;
  assign Pg24169 = Pg90;
  assign Pg24168 = Pg84;
  assign Pg24167 = Pg73;
  assign Pg24166 = Pg72;
  assign Pg24165 = Pg64;
  assign Pg24164 = Pg57;
  assign Pg24163 = Pg56;
  assign Pg24162 = Pg54;
  assign Pg24161 = Pg53;
  assign Pg23759 = Pg30331;
  assign Pg23683 = \[4421] ;
  assign Pg23652 = Pg30330;
  assign Pg23612 = Pg30329;
  assign Pg23002 = Pg30327;
  assign Pg21698 = Pg36;
  assign Pg21292 = \[4426] ;
  assign Pg21270 = \[4430] ;
  assign Pg21245 = \[4427] ;
  assign Pg21176 = \[4431] ;
  assign Pg20901 = \[4432] ;
  assign Pg20899 = \[4435] ;
  assign Pg20763 = \[4436] ;
  assign Pg20654 = \[4428] ;
  assign Pg20652 = \[4433] ;
  assign Pg20557 = \[4434] ;
  assign Pg20049 = \[4437] ;
  assign Pg18881 = \[4507] ;
  assign Pg18101 = Pg6746;
  assign Pg18100 = Pg6751;
  assign Pg18099 = Pg6745;
  assign Pg18098 = Pg6744;
  assign Pg18097 = Pg6747;
  assign Pg18096 = Pg6750;
  assign Pg18095 = Pg6749;
  assign Pg18094 = Pg6748;
  assign Pg18092 = Pg6753;
  assign Pg8403 = \[4651] ;
  assign Pg8353 = \[4651] ;
  assign Pg8283 = \[4658] ;
  assign Pg8235 = \[4658] ;
  assign Pg8178 = \[4661] ;
  assign Pg8132 = \[4661] ;
  assign n717_1 = Pg9048;
  assign n781 = Pg17715;
  assign n824 = Pg8920;
  assign n838_1 = Pg16656;
  assign n852_1 = Ng4571;
  assign n915_1 = Pg17743;
  assign n1023_1 = Pg16874;
  assign n1046_1 = Pg16627;
  assign n1137 = Pg17580;
  assign n1175_1 = Pg12368;
  assign n1178_1 = Pg17739;
  assign n1206 = Pg14694;
  assign n1229_1 = Pg17649;
  assign n1332 = Pg17320;
  assign n1359_1 = Pg14217;
  assign n1412_1 = Pg17722;
  assign n1424 = Pg8215;
  assign n1443 = Pg10527;
  assign n1482 = Pg16775;
  assign n1496 = Ng26960;
  assign n1514_1 = Pg12422;
  assign n1651_1 = Pg16744;
  assign n1718_1 = Pg9617;
  assign n1817 = Pg11678;
  assign n1841_1 = Pg17711;
  assign n1913_1 = Pg14673;
  assign n1921_1 = Pg17639;
  assign n1960_1 = Pg16722;
  assign n1984_1 = Pg17400;
  assign n2003_1 = Pg8344;
  assign n2032 = Pg13966;
  assign n2075_1 = Pg17760;
  assign n2097_1 = Pg8839;
  assign n2121_1 = Pg10122;
  assign n2125 = Pg12350;
  assign n2128_1 = Pg19357;
  assign n2151_1 = Pg7946;
  assign n2262 = Pg14597;
  assign n2290_1 = Pg14518;
  assign n2298 = Pg16924;
  assign n2310_1 = Pg17423;
  assign n2314 = Pg7245;
  assign n2332_1 = Pg9682;
  assign n2346_1 = Pg14125;
  assign n2433_1 = Pg11418;
  assign n2446_1 = Pg14096;
  assign n2459_1 = Pg8475;
  assign n2503_1 = Pg8870;
  assign n2620_1 = Ng26936;
  assign n2664_1 = Pg9497;
  assign n2702_1 = Pg11388;
  assign n2730_1 = Pg14779;
  assign n2753_1 = Pg11447;
  assign n2756_1 = Pg12923;
  assign n2775_1 = Pg8915;
  assign n2877_1 = Pg9251;
  assign n2886_1 = Pg8416;
  assign n2935_1 = Ng6974;
  assign n2938_1 = Pg11349;
  assign n2942_1 = Ng26959;
  assign n2976_1 = Pg17787;
  assign n3062_1 = Pg14189;
  assign n3080_1 = Pg8784;
  assign n3083_1 = Pg17519;
  assign n3220_1 = Pg19334;
  assign n3233_1 = Pg9743;
  assign n3271 = Pg7257;
  assign n3280 = Ng10384;
  assign n3283_1 = Pg17577;
  assign n3380_1 = Pg16693;
  assign n3383_1 = Pg17291;
  assign n3436_1 = Pg12238;
  assign n3469 = Pg16955;
  assign n3472 = Pg10306;
  assign n3481_1 = Pg17678;
  assign n3562 = Pg7260;
  assign n3596 = Pg13049;
  assign n3609_1 = Pg13259;
  assign n3628_1 = Pg8788;
  assign n3780_1 = Pg17607;
  assign n3901_1 = Pg14147;
  assign n3904_1 = Pg13039;
  assign n3972 = Pg14749;
  assign n3985_1 = Pg14635;
  assign n3993_1 = Pg16659;
  assign n4011 = Pg10500;
  assign n4040 = Pg14738;
  assign n4043 = Pg8719;
  assign n4067_1 = Pg12470;
  assign n4085_1 = Pg8279;
  assign n4152_1 = Pg12919;
  assign n4179 = Pg17871;
  assign n4207 = Pg8358;
  assign n4236_1 = Pg13068;
  assign n4264 = Pg14421;
  assign n4341_1 = Pg14451;
  assign n4394_1 = Pg8917;
  assign n4457 = Pg14705;
  assign n4490_1 = Pg17845;
  assign n4493 = Pg17674;
  assign n4496 = Pg8783;
  assign n4579 = Pg14662;
  assign n4641_1 = Pg13926;
  assign n4649 = Pg8918;
  assign n4732 = \[4507] ;
  assign n4771_1 = Pg13085;
  assign n4774_1 = Pg13099;
  assign n4847 = Pg13272;
  assign n4852_1 = Ng6972;
  assign n4856_1 = Pg8916;
  assign n4869 = Pg16748;
  assign n4878_1 = \[4661] ;
  assign n4891 = Pg7243;
  assign n4895_1 = Pg14167;
  assign n4949_1 = Pg7540;
  assign n4988 = Pg17764;
  assign n5061 = Pg13895;
  assign n5084_1 = Pg9019;
  assign n5108 = Pg8787;
  assign n5161 = Pg8291;
  assign n5238_1 = Pg12184;
  assign n5266_1 = Pg17646;
  assign n5270 = Ng25;
  assign n5323_1 = Pg17819;
  assign n5336_1 = Pg14201;
  assign n5354_1 = Pg17404;
  assign n5357_1 = Pg33435;
  assign n5386_1 = \[4658] ;
  assign n5390_1 = Pg17685;
  assign n5403_1 = Pg17316;
  assign n5522_1 = Ng26885;
  assign n5546_1 = Pg16624;
  assign n5663_1 = Pg17688;
  assign n5691 = \[4651] ;
  assign n5715_1 = Pg14828;
  assign n5777_1 = Ng4520;
  assign n5826 = Pg13906;
  assign n5829_1 = Pg33079;
  assign n5843_1 = Pg8785;
  assign n5860_1 = Pg9553;
  assign n5938_1 = Pg17778;
  assign n5995_1 = Pg17813;
  assign n6101 = Pg11770;
  assign n6124_1 = Pg16718;
  assign n6157 = Pg13881;
  assign n6170 = Pg16686;
  assign n6193 = Pg7916;
  assign n6294 = Pg12300;
  assign n6307 = Pg8919;
  assign n6374 = Pg17604;
  assign n6377 = Pg16603;
  assign n6400 = Pg13865;
  assign n6527 = Pg8789;
  assign n6556 = Pg9555;
  assign n6643 = Pg8786;
  always @ (posedge clock) begin
    Ng5057 <= n688;
    Ng2771 <= n693;
    Ng1882 <= n698_1;
    Ng2299 <= n703_1;
    Ng4040 <= n708_1;
    Ng2547 <= n713_1;
    Ng559 <= n717_1;
    Ng3243 <= n722_1;
    Ng452 <= n727_1;
    Ng3542 <= n732_1;
    Ng5232 <= n737_1;
    Ng5813 <= n742_1;
    Ng2907 <= n747_1;
    Ng1744 <= n752_1;
    Ng5909 <= n757_1;
    Ng1802 <= n762_1;
    Ng3554 <= n767_1;
    Ng6219 <= n772_1;
    Ng807 <= n777_1;
    Ng6031 <= n781;
    Ng847 <= n786_1;
    Ng976 <= n791_1;
    Ng4172 <= n796_1;
    Ng4372 <= n801_1;
    Ng3512 <= n806_1;
    Ng749 <= n811_1;
    Ng3490 <= n816_1;
    Pg12350 <= n821_1;
    Ng4235 <= n824;
    Ng1600 <= n829_1;
    Ng1714 <= n834_1;
    Pg14451 <= n838_1;
    Ng3155 <= n842_1;
    Ng2236 <= n847_1;
    Ng4555 <= n852_1;
    Ng3698 <= n857_1;
    Ng1736 <= n862_1;
    Ng1968 <= n867_1;
    Ng4621 <= n872_1;
    Ng5607 <= n877_1;
    Ng2657 <= n882_1;
    Pg12300 <= n887_1;
    Ng490 <= n891_1;
    Ng311 <= n896_1;
    Ng772 <= n901_1;
    Ng5587 <= n906_1;
    Ng6177 <= n911_1;
    Ng6377 <= n915_1;
    Ng3167 <= n920_1;
    Ng5615 <= n925_1;
    Ng4567 <= n930;
    Ng3457 <= n935_1;
    Ng6287 <= n940_1;
    Pg7946 <= n945_1;
    Ng2563 <= n949_1;
    Ng4776 <= n954_1;
    Ng4593 <= n959_1;
    Ng6199 <= n964_1;
    Ng2295 <= n969_1;
    Ng1384 <= n974_1;
    Ng1339 <= n979_1;
    Ng5180 <= n984_1;
    Ng2844 <= n989_1;
    Ng1024 <= n994_1;
    Ng5591 <= n999_1;
    Ng3598 <= n1004_1;
    Ng4264 <= n1009_1;
    Ng767 <= n1014_1;
    Ng5853 <= n1019_1;
    Pg13865 <= n1023_1;
    Ng2089 <= n1027_1;
    Ng4933 <= n1032_1;
    Ng4521 <= n1037_1;
    Ng5507 <= n1042_1;
    Pg16656 <= n1046_1;
    Ng6291 <= n1050_1;
    Ng294 <= n1055_1;
    Ng5559 <= n1060;
    Pg9617 <= n1065_1;
    Pg9741 <= n1069_1;
    Ng3813 <= n1073_1;
    Ng562 <= n1078_1;
    Ng608 <= n1083_1;
    Ng1205 <= n1088_1;
    Ng3909 <= n1093_1;
    Ng6259 <= n1098;
    Ng5905 <= n1103;
    Ng921 <= n1108_1;
    Ng2955 <= n1113_1;
    Ng203 <= n1118_1;
    Ng1099 <= n1123;
    Ng4878 <= n1128;
    Ng5204 <= n1133_1;
    Pg17604 <= n1137;
    Ng3606 <= n1141_1;
    Ng1926 <= n1146_1;
    Ng6215 <= n1151_1;
    Ng3586 <= n1156_1;
    Ng291 <= n1161;
    Ng4674 <= n1166_1;
    Ng3570 <= n1171;
    Pg9048 <= n1175_1;
    Pg17607 <= n1178_1;
    Ng1862 <= n1182_1;
    Ng676 <= n1187_1;
    Ng843 <= n1192_1;
    Ng4332 <= n1197_1;
    Ng4153 <= n1202;
    Pg17711 <= n1206;
    Ng6336 <= n1210;
    Ng622 <= n1215_1;
    Ng3506 <= n1220_1;
    Ng4558 <= n1225;
    Pg17685 <= n1229_1;
    Ng3111 <= n1233_1;
    \[4430]  <= n1238_1;
    Ng26936 <= n1243_1;
    Ng939 <= n1248_1;
    Ng278 <= n1253_1;
    Ng4492 <= n1258_1;
    Ng4864 <= n1263_1;
    Ng1036 <= n1268_1;
    \[4427]  <= n1273_1;
    Ng1178 <= n1278_1;
    Ng3239 <= n1283_1;
    Ng718 <= n1288_1;
    Ng6195 <= n1293_1;
    Ng1135 <= n1298_1;
    Ng6395 <= n1303_1;
    \[4415]  <= n1308_1;
    Ng554 <= n1313_1;
    Ng496 <= n1318_1;
    Ng3853 <= n1323_1;
    Ng5134 <= n1328_1;
    Pg17404 <= n1332;
    Pg8344 <= n1336_1;
    Ng2485 <= n1340;
    Ng925 <= n1345_1;
    Ng48 <= n1350_1;
    Ng5555 <= n1355_1;
    Pg14096 <= n1359_1;
    Ng1798 <= n1363_1;
    Ng4076 <= n1368_1;
    Ng2941 <= n1373_1;
    Ng3905 <= n1378_1;
    Ng763 <= n1383_1;
    Ng6255 <= n1388_1;
    Ng4375 <= n1393_1;
    Ng4871 <= n1398_1;
    Ng4722 <= n1403_1;
    Ng590 <= n1408_1;
    Pg13099 <= n1412_1;
    Ng1632 <= n1416_1;
    Pg12238 <= n1421_1;
    Ng3100 <= n1424;
    Ng1495 <= n1429_1;
    Ng1437 <= n1434;
    Ng6154 <= n1439_1;
    Ng1579 <= n1443;
    Ng5567 <= n1448;
    Ng1752 <= n1453;
    Ng1917 <= n1458_1;
    Ng744 <= n1463;
    Ng4737 <= n1468_1;
    \[4661]  <= n1473;
    Ng6267 <= n1478_1;
    Pg16659 <= n1482;
    Ng1442 <= n1486;
    Ng5965 <= n1491_1;
    Ng4477 <= n1496;
    Pg10500 <= n1501_1;
    Ng4643 <= n1505_1;
    Ng5264 <= n1510_1;
    Pg14779 <= n1514_1;
    Ng2610 <= n1518_1;
    Ng5160 <= n1523_1;
    Ng5933 <= n1528;
    Ng1454 <= n1533_1;
    Ng753 <= n1538;
    Ng1296 <= n1543_1;
    Ng3151 <= n1548_1;
    Ng2980 <= n1553;
    Ng6727 <= n1558_1;
    Ng3530 <= n1563_1;
    Ng4104 <= n1568;
    Ng1532 <= n1573;
    Pg9251 <= n1578_1;
    Ng2177 <= n1582_1;
    Ng52 <= n1587_1;
    Ng4754 <= n1592_1;
    Ng1189 <= n1597_1;
    Ng2287 <= n1602_1;
    Ng4273 <= n1607_1;
    Ng1389 <= n1612_1;
    Ng1706 <= n1617_1;
    Ng5835 <= n1622_1;
    Ng1171 <= n1627_1;
    Ng4269 <= n1632_1;
    Ng2399 <= n1637;
    Ng4983 <= n1642_1;
    Ng5611 <= n1647_1;
    Pg16627 <= n1651_1;
    Ng4572 <= n1655_1;
    Ng3143 <= n1660_1;
    Ng2898 <= n1665;
    Ng3343 <= n1670_1;
    Ng3235 <= n1675_1;
    Ng4543 <= n1680;
    Ng3566 <= n1685_1;
    Ng4534 <= n1690_1;
    Ng4961 <= n1695_1;
    Ng4927 <= n1700_1;
    Ng2259 <= n1705;
    Ng2819 <= n1710_1;
    Pg7257 <= n1715_1;
    Ng5802 <= n1718_1;
    Ng2852 <= n1723;
    Ng417 <= n1728;
    Ng681 <= n1733_1;
    Ng437 <= n1738;
    Ng351 <= n1743_1;
    Ng5901 <= n1748;
    Ng2886 <= n1753_1;
    Ng3494 <= n1758_1;
    Ng5511 <= n1763_1;
    Ng3518 <= n1768_1;
    Ng1604 <= n1773_1;
    Ng5092 <= n1778;
    Ng4831 <= n1783_1;
    Ng4382 <= n1788_1;
    Ng6386 <= n1793_1;
    Ng479 <= n1798_1;
    Ng3965 <= n1803;
    Ng4749 <= n1808_1;
    Ng2008 <= n1813_1;
    Ng736 <= n1817;
    Ng3933 <= n1822;
    Ng222 <= n1827_1;
    Ng3050 <= n1832_1;
    Ng1052 <= n1837_1;
    Pg17580 <= n1841_1;
    Ng2122 <= n1845_1;
    Ng2465 <= n1850;
    Ng5889 <= n1855_1;
    Ng4495 <= n1860_1;
    Pg8719 <= n1865_1;
    Ng4653 <= n1869_1;
    Ng3179 <= n1874;
    Ng1728 <= n1879_1;
    Ng2433 <= n1884_1;
    Ng3835 <= n1889_1;
    Ng6187 <= n1894;
    Ng4917 <= n1899;
    Ng1070 <= n1904;
    Ng822 <= n1909_1;
    Pg17715 <= n1913_1;
    Ng914 <= n1917;
    Ng5339 <= n1921_1;
    Ng4164 <= n1926;
    Ng969 <= n1931_1;
    Ng2807 <= n1936_1;
    Ng4054 <= n1941_1;
    Ng6191 <= n1946;
    Ng5077 <= n1951;
    Ng5523 <= n1956_1;
    Ng3680 <= n1960_1;
    Ng6637 <= n1965_1;
    Ng174 <= n1970_1;
    Ng1682 <= n1975_1;
    Ng355 <= n1980_1;
    Ng1087 <= n1984_1;
    Ng1105 <= n1989;
    Ng2342 <= n1994_1;
    Ng6307 <= n1999_1;
    Ng3802 <= n2003_1;
    Ng6159 <= n2008_1;
    Ng2255 <= n2013_1;
    Ng2815 <= n2018;
    Ng911 <= n2023_1;
    Ng43 <= n2028;
    Pg16775 <= n2032;
    Ng1748 <= n2036_1;
    Ng5551 <= n2041;
    Ng3558 <= n2046_1;
    Ng5499 <= n2051_1;
    Ng2960 <= n2056;
    Ng3901 <= n2061;
    Ng4888 <= n2066;
    Ng6251 <= n2071;
    Pg17649 <= n2075_1;
    Ng1373 <= n2079_1;
    Pg8215 <= n2084_1;
    Ng157 <= n2088_1;
    Ng2783 <= n2093_1;
    Ng4281 <= n2097_1;
    Ng3574 <= n2102;
    Ng2112 <= n2107_1;
    Ng1283 <= n2112;
    Ng433 <= n2117_1;
    Ng4297 <= n2121_1;
    Pg14738 <= n2125;
    Pg13272 <= n2128_1;
    Ng758 <= n2132;
    Ng4639 <= n2137;
    Ng6537 <= n2142_1;
    Ng5543 <= n2147_1;
    Pg8475 <= n2151_1;
    Ng5961 <= n2155;
    Ng6243 <= n2160_1;
    Ng632 <= n2165;
    Pg12919 <= n2170_1;
    Ng3889 <= n2174;
    Ng3476 <= n2179;
    Ng1664 <= n2184;
    Ng1246 <= n2189;
    Ng6629 <= n2194_1;
    Ng246 <= n2199;
    Ng4049 <= n2204_1;
    Pg7260 <= n2209_1;
    Ng2932 <= n2213;
    Ng4575 <= n2218_1;
    Ng4098 <= n2223_1;
    Ng4498 <= n2228_1;
    Ng528 <= n2233_1;
    Ng16 <= n2238_1;
    Ng3139 <= n2243_1;
    \[4432]  <= n2248_1;
    Ng4584 <= n2253_1;
    Ng142 <= n2258_1;
    Pg17639 <= n2262;
    Ng5831 <= n2266_1;
    Ng239 <= n2271_1;
    Ng1216 <= n2276_1;
    Ng2848 <= n2281_1;
    Ng5022 <= n2286;
    Pg16955 <= n2290_1;
    Ng1030 <= n2294_1;
    Pg13881 <= n2298;
    Ng3231 <= n2302_1;
    Pg9817 <= n2307;
    Ng1430 <= n2310_1;
    Ng4452 <= n2314;
    Ng2241 <= n2319_1;
    Ng1564 <= n2324;
    Pg9680 <= n2329_1;
    Ng6148 <= n2332_1;
    Ng6649 <= n2337;
    Ng110 <= n2342_1;
    Pg14147 <= n2346_1;
    Ng225 <= n2350;
    Ng4486 <= n2355_1;
    Ng4504 <= n2360;
    Ng5873 <= n2365;
    Ng5037 <= n2370_1;
    Ng2319 <= n2375;
    Ng5495 <= n2380_1;
    Pg11770 <= n2385_1;
    Ng5208 <= n2389;
    Ng5579 <= n2394_1;
    Ng5869 <= n2399_1;
    Ng1589 <= n2404_1;
    Ng5752 <= n2409_1;
    Ng6279 <= n2414_1;
    Ng5917 <= n2419_1;
    Ng2975 <= n2424_1;
    Ng6167 <= n2429;
    Pg13966 <= n2433_1;
    Ng2599 <= n2437_1;
    Ng1448 <= n2442;
    Pg14125 <= n2446_1;
    Ng2370 <= n2450_1;
    Ng5164 <= n2455;
    Ng1333 <= n2459_1;
    Ng153 <= n2464_1;
    Ng6549 <= n2469_1;
    Ng4087 <= n2474_1;
    Ng4801 <= n2479_1;
    Ng2984 <= n2484_1;
    Ng3961 <= n2489_1;
    Ng962 <= n2494;
    Ng101 <= n2499;
    Pg8918 <= n2503_1;
    Ng6625 <= n2507_1;
    Ng51 <= n2512;
    Ng1018 <= n2517_1;
    Pg17320 <= n2522_1;
    Ng4045 <= n2526_1;
    Ng1467 <= n2531;
    Ng2461 <= n2536_1;
    Ng2756 <= n2541_1;
    Ng5990 <= n2546_1;
    Ng1256 <= n2551_1;
    Ng5029 <= n2556;
    Ng6519 <= n2561_1;
    Ng1816 <= n2566;
    Ng4369 <= n2571_1;
    Ng4578 <= n2576_1;
    Ng4459 <= n2581;
    Ng3831 <= n2586_1;
    Ng2514 <= n2591_1;
    Ng3288 <= n2596;
    Ng2403 <= n2601_1;
    Ng2145 <= n2606_1;
    Ng1700 <= n2611_1;
    Ng513 <= n2616_1;
    Ng2841 <= n2620_1;
    Ng5297 <= n2625_1;
    Ng2763 <= n2630_1;
    Ng4793 <= n2635_1;
    Ng952 <= n2640_1;
    Ng1263 <= n2645_1;
    Ng1950 <= n2650_1;
    Ng5138 <= n2655_1;
    Ng2307 <= n2660_1;
    Ng5109 <= n2664_1;
    Pg8398 <= n2669_1;
    Ng4664 <= n2673_1;
    Ng2223 <= n2678_1;
    Ng5808 <= n2683_1;
    Ng6645 <= n2688_1;
    Ng2016 <= n2693_1;
    Ng3873 <= n2698_1;
    Pg13926 <= n2702_1;
    Ng2315 <= n2706_1;
    Ng2811 <= n2711_1;
    Ng5957 <= n2716_1;
    Ng2047 <= n2721_1;
    Ng3869 <= n2726_1;
    Pg17760 <= n2730_1;
    Ng5575 <= n2734_1;
    Ng46 <= n2739_1;
    Ng3752 <= n2744_1;
    Ng3917 <= n2749;
    Pg8783 <= n2753_1;
    Ng1585 <= n2756_1;
    Ng4388 <= n2761_1;
    Ng6275 <= n2766_1;
    Ng6311 <= n2771_1;
    Pg8916 <= n2775_1;
    Ng1041 <= n2779_1;
    Ng2595 <= n2784_1;
    Ng2537 <= n2789_1;
    \[4426]  <= n2794_1;
    Ng4430 <= n2799_1;
    Ng4564 <= n2804_1;
    Ng4826 <= n2809_1;
    Ng6239 <= n2814_1;
    Ng232 <= n2819;
    Ng5268 <= n2824_1;
    Ng6545 <= n2829_1;
    Ng2417 <= n2834_1;
    Ng1772 <= n2839_1;
    Ng5052 <= n2844_1;
    Pg9615 <= n2849_1;
    Ng1890 <= n2853_1;
    Ng2629 <= n2858_1;
    Ng572 <= n2863_1;
    Ng2130 <= n2868_1;
    Ng4108 <= n2873_1;
    Ng4308 <= n2877_1;
    Ng475 <= n2882_1;
    Ng990 <= n2886_1;
    Ng45 <= n2891_1;
    Pg12184 <= n2896;
    Ng3990 <= n2900_1;
    Ng5881 <= n2905_1;
    Ng1992 <= n2910_1;
    Ng3171 <= n2915_1;
    Ng812 <= n2920_1;
    Ng832 <= n2925_1;
    Ng5897 <= n2930_1;
    Ng4571 <= n2935_1;
    Pg13895 <= n2938_1;
    Ng4455 <= n2942_1;
    Ng2902 <= n2947_1;
    Ng333 <= n2952_1;
    Ng168 <= n2957_1;
    Ng2823 <= n2962_1;
    Ng3684 <= n2967_1;
    Ng3639 <= n2972_1;
    Pg14597 <= n2976_1;
    Ng3338 <= n2980_1;
    Ng5406 <= n2985;
    Ng269 <= n2990_1;
    Ng401 <= n2995_1;
    Ng6040 <= n3000_1;
    Ng441 <= n3005_1;
    Pg9553 <= n3010_1;
    Ng3808 <= n3014_1;
    Ng10384 <= n3019_1;
    Ng3957 <= n3024_1;
    Ng4093 <= n3029_1;
    Ng1760 <= n3034_1;
    Pg12422 <= n3039_1;
    Ng160 <= n3043_1;
    Ng2279 <= n3048_1;
    Ng3498 <= n3053_1;
    Ng586 <= n3058;
    Pg14201 <= n3062_1;
    Ng2619 <= n3066;
    Ng1183 <= n3071_1;
    Ng1608 <= n3076;
    Pg8785 <= n3080_1;
    Pg17577 <= n3083_1;
    Ng1779 <= n3087;
    Ng2652 <= n3092_1;
    Ng2193 <= n3097;
    Ng2393 <= n3102;
    Ng661 <= n3107_1;
    Ng4950 <= n3112;
    Ng5535 <= n3117;
    Ng2834 <= n3122_1;
    Ng1361 <= n3127;
    Ng6235 <= n3132_1;
    Ng1146 <= n3137_1;
    Ng2625 <= n3142;
    Ng150 <= n3147;
    Ng1696 <= n3152_1;
    Ng6555 <= n3157_1;
    Pg14189 <= n3162;
    Ng3881 <= n3166;
    Ng6621 <= n3171_1;
    Ng3470 <= n3176_1;
    Ng3897 <= n3181_1;
    Ng518 <= n3186;
    Ng538 <= n3191;
    Ng2606 <= n3196;
    Ng1472 <= n3201;
    Ng542 <= n3206;
    Ng5188 <= n3211_1;
    Ng5689 <= n3216;
    Pg13259 <= n3220_1;
    Ng405 <= n3224;
    Ng5216 <= n3229_1;
    Ng6494 <= n3233_1;
    Ng4669 <= n3238_1;
    Ng996 <= n3243_1;
    Ng4531 <= n3248;
    Ng2860 <= n3253_1;
    Ng4743 <= n3258;
    Ng6593 <= n3263_1;
    Pg8291 <= n3268;
    Ng4411 <= n3271;
    Ng1413 <= n3276_1;
    Ng26960 <= n3280;
    Pg13039 <= n3283_1;
    Ng6641 <= n3287_1;
    Ng1936 <= n3292_1;
    Ng55 <= n3297;
    Ng504 <= n3302_1;
    Ng2587 <= n3307;
    Ng4480 <= n3312;
    Ng2311 <= n3317_1;
    Ng3602 <= n3322_1;
    Ng5571 <= n3327_1;
    Ng3578 <= n3332;
    Pg9555 <= n3337_1;
    Ng5827 <= n3341_1;
    Ng3582 <= n3346_1;
    Ng6271 <= n3351_1;
    Ng4688 <= n3356;
    Ng2380 <= n3361_1;
    Ng5196 <= n3366;
    Ng3227 <= n3371_1;
    Ng2020 <= n3376;
    Pg14518 <= n3380_1;
    Pg17316 <= n3383_1;
    Ng6541 <= n3387;
    Ng3203 <= n3392_1;
    Ng1668 <= n3397_1;
    Ng4760 <= n3402_1;
    Ng262 <= n3407;
    Ng1840 <= n3412_1;
    Ng5467 <= n3417_1;
    Ng460 <= n3422;
    Ng6209 <= n3427_1;
    \[4436]  <= n3432;
    Pg14662 <= n3436_1;
    Ng655 <= n3440_1;
    Ng3502 <= n3445;
    Ng2204 <= n3450_1;
    Ng5256 <= n3455_1;
    Ng4608 <= n3460;
    Ng794 <= n3465_1;
    Pg13906 <= n3469;
    Ng4423 <= n3472;
    Ng3689 <= n3477_1;
    Ng5685 <= n3481_1;
    Ng703 <= n3486;
    Ng862 <= n3491_1;
    Ng3247 <= n3496;
    Ng2040 <= n3501_1;
    Ng4146 <= n3506;
    Ng4633 <= n3511_1;
    Pg7916 <= n3516_1;
    Ng4732 <= n3520_1;
    Pg9497 <= n3525_1;
    Ng5817 <= n3529_1;
    Ng2351 <= n3534_1;
    Ng2648 <= n3539_1;
    Ng6736 <= n3544;
    Ng4944 <= n3549;
    Ng4072 <= n3554_1;
    Pg7540 <= n3559;
    Ng4443 <= n3562;
    Ng3466 <= n3567_1;
    Ng4116 <= n3572_1;
    Ng5041 <= n3577_1;
    Ng4434 <= n3582;
    Ng3827 <= n3587_1;
    Ng6500 <= n3592;
    Pg17813 <= n3596;
    Ng3133 <= n3600;
    Ng3333 <= n3605;
    Ng979 <= n3609_1;
    Ng4681 <= n3614;
    Ng298 <= n3619_1;
    Ng2667 <= n3624_1;
    Pg8789 <= n3628_1;
    Ng1894 <= n3632;
    Ng2988 <= n3637;
    Ng3538 <= n3642_1;
    Ng301 <= n3647_1;
    Ng341 <= n3652_1;
    Ng827 <= n3657_1;
    Pg17291 <= n3662;
    Ng2555 <= n3666;
    Ng5011 <= n3671;
    Ng199 <= n3676_1;
    Ng6523 <= n3681_1;
    Ng1526 <= n3686_1;
    Ng4601 <= n3691;
    Ng854 <= n3696;
    Ng1484 <= n3701;
    Ng4922 <= n3706_1;
    Ng5080 <= n3711;
    Ng5863 <= n3716_1;
    Ng4581 <= n3721_1;
    Ng2518 <= n3726;
    Ng2567 <= n3731_1;
    Ng568 <= n3736_1;
    Ng3263 <= n3741_1;
    Ng6613 <= n3746;
    Ng6044 <= n3751;
    Ng6444 <= n3756;
    Ng2965 <= n3761_1;
    Ng5857 <= n3766_1;
    Ng1616 <= n3771_1;
    Ng890 <= n3776_1;
    Pg17646 <= n3780_1;
    Ng3562 <= n3784_1;
    Pg10122 <= n3789_1;
    Ng1404 <= n3793_1;
    Ng3817 <= n3798_1;
    Ng93 <= n3803_1;
    Ng4501 <= n3808;
    Ng287 <= n3813_1;
    Ng2724 <= n3818_1;
    Ng4704 <= n3823_1;
    Ng22 <= n3828_1;
    Ng2878 <= n3833_1;
    Ng5220 <= n3838_1;
    Ng617 <= n3843_1;
    Pg12368 <= n3848;
    Ng316 <= n3852_1;
    Ng1277 <= n3857;
    Ng6513 <= n3862_1;
    Ng336 <= n3867_1;
    Ng2882 <= n3872_1;
    Ng933 <= n3877_1;
    Ng1906 <= n3882_1;
    Ng305 <= n3887_1;
    Ng8 <= n3892;
    Ng2799 <= n3897;
    Pg14167 <= n3901_1;
    Pg17787 <= n3904_1;
    Ng4912 <= n3908;
    Ng4157 <= n3913;
    Ng2541 <= n3918_1;
    Ng2153 <= n3923_1;
    Ng550 <= n3928;
    Ng255 <= n3933_1;
    Ng1945 <= n3938;
    Ng5240 <= n3943_1;
    Ng1478 <= n3948_1;
    Ng3863 <= n3953_1;
    Ng1959 <= n3958;
    Ng3480 <= n3963_1;
    Ng6653 <= n3968;
    Pg17764 <= n3972;
    Ng2864 <= n3976_1;
    Ng4894 <= n3981;
    Pg17678 <= n3985_1;
    Ng3857 <= n3989;
    Pg16693 <= n3993_1;
    Ng499 <= n3997_1;
    Ng1002 <= n4002;
    Ng776 <= n4007;
    Ng1236 <= n4011;
    Ng4646 <= n4016;
    Ng2476 <= n4021_1;
    Ng1657 <= n4026;
    Ng2375 <= n4031_1;
    Ng63 <= n4036_1;
    Pg17739 <= n4040;
    Ng358 <= n4043;
    Ng896 <= n4048_1;
    Ng283 <= n4053;
    Ng3161 <= n4058_1;
    Ng2384 <= n4063_1;
    Pg14828 <= n4067_1;
    Ng4616 <= n4071_1;
    Ng4561 <= n4076_1;
    Ng2024 <= n4081;
    Ng3451 <= n4085_1;
    Ng2795 <= n4090;
    Ng613 <= n4095_1;
    Ng4527 <= n4100_1;
    Ng1844 <= n4105;
    Ng5937 <= n4110_1;
    Ng4546 <= n4115_1;
    Ng2523 <= n4120_1;
    Pg11349 <= n4125;
    Ng2643 <= n4129_1;
    Ng1489 <= n4134_1;
    Pg8358 <= n4139_1;
    Ng2551 <= n4143;
    Ng5156 <= n4148;
    \[4421]  <= n4152_1;
    Pg8279 <= n4157_1;
    Pg8839 <= n4161;
    Ng1955 <= n4165_1;
    Ng6049 <= n4170_1;
    Ng2273 <= n4175;
    Pg14749 <= n4179;
    Ng4771 <= n4183_1;
    Ng6098 <= n4188;
    Ng3147 <= n4193;
    Ng3347 <= n4198_1;
    Ng2269 <= n4203_1;
    Ng191 <= n4207;
    Ng2712 <= n4212_1;
    Ng626 <= n4217_1;
    Ng2729 <= n4222_1;
    Ng5357 <= n4227_1;
    Ng4991 <= n4232;
    Pg17819 <= n4236_1;
    Ng4709 <= n4240;
    Ng2927 <= n4245_1;
    Ng4340 <= n4250;
    Ng5929 <= n4255;
    Ng4907 <= n4260;
    Pg16874 <= n4264;
    Ng4035 <= n4268_1;
    Ng2946 <= n4273;
    Ng918 <= n4278;
    Ng4082 <= n4283_1;
    Pg9743 <= n4288_1;
    Ng2036 <= n4292_1;
    Ng577 <= n4297_1;
    Ng1620 <= n4302_1;
    Ng2831 <= n4307_1;
    Ng667 <= n4312_1;
    Ng930 <= n4317_1;
    Ng3937 <= n4322_1;
    Ng817 <= n4327_1;
    Ng1249 <= n4332_1;
    Ng837 <= n4337_1;
    Pg16924 <= n4341_1;
    Ng599 <= n4345_1;
    Ng5475 <= n4350_1;
    Ng739 <= n4355_1;
    Ng5949 <= n4360_1;
    Ng6682 <= n4365_1;
    Ng904 <= n4370;
    Ng2873 <= n4375;
    Ng1854 <= n4380_1;
    Ng5084 <= n4385_1;
    Ng5603 <= n4390;
    Pg8870 <= n4394_1;
    Ng2495 <= n4398_1;
    Ng2437 <= n4403_1;
    Ng2102 <= n4408;
    Ng2208 <= n4413;
    Ng2579 <= n4418_1;
    Ng4064 <= n4423;
    Ng4899 <= n4428_1;
    Ng2719 <= n4433_1;
    Ng4785 <= n4438;
    Ng5583 <= n4443_1;
    Ng781 <= n4448;
    Ng6173 <= n4453;
    Pg17743 <= n4457;
    Ng2917 <= n4461;
    Ng686 <= n4466;
    Ng1252 <= n4471;
    Ng671 <= n4476;
    Ng2265 <= n4481;
    Ng6283 <= n4486_1;
    Pg14705 <= n4490_1;
    Pg17519 <= n4493;
    Pg8784 <= n4496;
    Ng5527 <= n4500;
    Ng4489 <= n4505;
    Ng1974 <= n4510_1;
    Ng1270 <= n4515_1;
    Ng4966 <= n4520;
    Ng6227 <= n4525;
    Ng3929 <= n4530_1;
    Ng5503 <= n4535_1;
    Ng4242 <= n4540_1;
    Ng5925 <= n4545;
    Ng1124 <= n4550_1;
    Ng4955 <= n4555;
    Ng5224 <= n4560;
    Ng2012 <= n4565;
    Ng6203 <= n4570_1;
    Ng5120 <= n4575;
    Pg17674 <= n4579;
    Ng2389 <= n4583;
    Ng4438 <= n4588_1;
    Ng2429 <= n4593_1;
    Ng2787 <= n4598;
    Ng1287 <= n4603;
    Ng2675 <= n4608;
    \[4507]  <= n4613;
    Ng4836 <= n4618;
    Ng1199 <= n4623;
    Pg19357 <= n4628;
    Ng5547 <= n4632_1;
    Ng2138 <= n4637_1;
    Pg16744 <= n4641_1;
    Ng2338 <= n4645;
    Pg8919 <= n4649;
    Ng6247 <= n4653_1;
    Ng2791 <= n4658;
    Ng3949 <= n4663_1;
    Ng1291 <= n4668;
    Ng5945 <= n4673_1;
    Ng5244 <= n4678;
    Ng2759 <= n4683;
    Ng6741 <= n4688;
    Ng785 <= n4693;
    Ng1259 <= n4698;
    Ng3484 <= n4703_1;
    Ng209 <= n4708;
    Ng6609 <= n4713_1;
    Ng5517 <= n4718;
    Ng2449 <= n4723_1;
    Ng2575 <= n4728;
    Ng65 <= n4732;
    Ng2715 <= n4737_1;
    Ng936 <= n4742_1;
    Ng2098 <= n4747_1;
    Ng4462 <= n4752_1;
    Ng604 <= n4757_1;
    Ng6589 <= n4762;
    Ng1886 <= n4767_1;
    Pg17845 <= n4771_1;
    Pg17871 <= n4774_1;
    Ng429 <= n4778_1;
    Ng1870 <= n4783_1;
    Ng4249 <= n4788;
    Ng1825 <= n4793_1;
    Ng1008 <= n4798;
    Ng4392 <= n4803;
    Ng3546 <= n4808_1;
    Ng5236 <= n4813_1;
    Ng1768 <= n4818_1;
    Ng4854 <= n4823_1;
    Ng3925 <= n4828;
    Ng6509 <= n4833_1;
    Ng732 <= n4838_1;
    Ng2504 <= n4843;
    Ng1322 <= n4847;
    Ng4520 <= n4852_1;
    Pg8917 <= n4856_1;
    Ng2185 <= n4860_1;
    Ng37 <= n4865;
    Ng4031 <= n4869;
    Ng2070 <= n4874;
    \[4658]  <= n4878_1;
    Ng4176 <= n4883_1;
    Pg11418 <= n4888_1;
    Ng4405 <= n4891;
    Ng872 <= n4895_1;
    Ng6181 <= n4900_1;
    Ng6381 <= n4905;
    Ng4765 <= n4910_1;
    Ng5563 <= n4915_1;
    Ng1395 <= n4920;
    Ng1913 <= n4925;
    Ng2331 <= n4930_1;
    Ng6263 <= n4935_1;
    Ng50 <= n4940_1;
    Ng3945 <= n4945_1;
    Ng347 <= n4949_1;
    Ng4473 <= n4954_1;
    Ng1266 <= n4959_1;
    Ng5489 <= n4964_1;
    Ng714 <= n4969_1;
    Ng2748 <= n4974;
    Ng5471 <= n4979;
    Ng4540 <= n4984_1;
    Ng6723 <= n4988;
    Ng6605 <= n4993;
    Ng2445 <= n4998_1;
    Ng2173 <= n5003;
    Pg9019 <= n5008;
    Ng2491 <= n5012_1;
    Ng4849 <= n5017;
    Ng2169 <= n5022;
    Ng2283 <= n5027;
    Ng6585 <= n5032;
    \[4428]  <= n5037;
    Ng2407 <= n5042;
    Ng2868 <= n5047_1;
    Ng2767 <= n5052_1;
    Ng1783 <= n5057_1;
    Pg16718 <= n5061;
    Ng1312 <= n5065;
    Ng5212 <= n5070_1;
    Ng4245 <= n5075_1;
    Ng645 <= n5080;
    Ng4291 <= n5084_1;
    \[4435]  <= n5089_1;
    Ng182 <= n5094_1;
    Ng1129 <= n5099;
    Ng2227 <= n5104;
    Pg8788 <= n5108;
    Ng2246 <= n5112;
    Ng1830 <= n5117;
    Ng3590 <= n5122_1;
    Ng392 <= n5127;
    Ng1592 <= n5132_1;
    Ng6505 <= n5137_1;
    Ng1221 <= n5142_1;
    Ng5921 <= n5147_1;
    \[4431]  <= n5152_1;
    Ng146 <= n5157;
    Ng218 <= n5161;
    Ng1932 <= n5166;
    Ng1624 <= n5171;
    Ng5062 <= n5176_1;
    Ng5462 <= n5181_1;
    Ng2689 <= n5186_1;
    Ng6573 <= n5191;
    Ng1677 <= n5196_1;
    Ng2028 <= n5201_1;
    Ng2671 <= n5206_1;
    Pg10527 <= n5211_1;
    Pg7243 <= n5215_1;
    Ng1848 <= n5219_1;
    \[4434]  <= n5224_1;
    Ng5485 <= n5229_1;
    Ng2741 <= n5234_1;
    Pg11678 <= n5238_1;
    Ng2638 <= n5242_1;
    Ng4122 <= n5247_1;
    Ng4322 <= n5252_1;
    Ng5941 <= n5257_1;
    Ng2108 <= n5262_1;
    Pg13068 <= n5266_1;
    Ng25 <= n5270;
    Ng1644 <= n5274_1;
    Ng595 <= n5279;
    Ng2217 <= n5284_1;
    Ng1319 <= n5289;
    Ng2066 <= n5294;
    Ng1152 <= n5299_1;
    Ng5252 <= n5304_1;
    Ng2165 <= n5309_1;
    Ng2571 <= n5314;
    Ng5176 <= n5319_1;
    Pg14673 <= n5323_1;
    Ng1211 <= n5327_1;
    Ng2827 <= n5332_1;
    Pg14217 <= n5336_1;
    Ng4859 <= n5340_1;
    Ng424 <= n5345_1;
    Ng1274 <= n5350_1;
    Pg17423 <= n5354_1;
    Ng85 <= n5357_1;
    Ng2803 <= n5362_1;
    Ng1821 <= n5367_1;
    Ng2509 <= n5372_1;
    Ng5073 <= n5377_1;
    Ng1280 <= n5382_1;
    \[4651]  <= n5386_1;
    Pg13085 <= n5390_1;
    Ng6633 <= n5394_1;
    Ng5124 <= n5399_1;
    Pg17400 <= n5403_1;
    Ng6303 <= n5407_1;
    Ng5069 <= n5412;
    Ng2994 <= n5417_1;
    Ng650 <= n5422_1;
    Ng1636 <= n5427_1;
    Ng3921 <= n5432;
    Ng2093 <= n5437_1;
    Ng6732 <= n5442_1;
    Ng1306 <= n5447;
    Ng1061 <= n5452_1;
    Ng3462 <= n5457;
    Ng2181 <= n5462_1;
    Ng956 <= n5467_1;
    Ng1756 <= n5472_1;
    Ng5849 <= n5477_1;
    Ng4112 <= n5482_1;
    Ng2685 <= n5487_1;
    Ng2197 <= n5492_1;
    Ng2421 <= n5497_1;
    Ng1046 <= n5502_1;
    Ng482 <= n5507_1;
    Ng4401 <= n5512_1;
    Ng1514 <= n5517_1;
    Ng329 <= n5522_1;
    Ng6565 <= n5527_1;
    Ng2950 <= n5532_1;
    Ng1345 <= n5537_1;
    Ng6533 <= n5542;
    Pg14421 <= n5546_1;
    Ng4727 <= n5550_1;
    Pg12470 <= n5555_1;
    Ng1536 <= n5559_1;
    Ng3941 <= n5564_1;
    Ng370 <= n5569_1;
    Ng5694 <= n5574;
    Ng1858 <= n5579_1;
    Ng446 <= n5584_1;
    Ng3219 <= n5589_1;
    Ng1811 <= n5594;
    Ng6601 <= n5599_1;
    Ng2441 <= n5604_1;
    Ng1874 <= n5609_1;
    Ng4349 <= n5614_1;
    Ng6581 <= n5619_1;
    Ng6597 <= n5624;
    Ng3610 <= n5629;
    Ng2890 <= n5634_1;
    Ng1978 <= n5639;
    Ng1612 <= n5644_1;
    Ng112 <= n5649_1;
    Ng2856 <= n5654_1;
    Ng1982 <= n5659;
    Pg17722 <= n5663_1;
    Ng5228 <= n5667;
    Ng4119 <= n5672;
    Ng6390 <= n5677_1;
    Ng1542 <= n5682_1;
    Ng4258 <= n5687_1;
    Ng4818 <= n5691;
    Ng5033 <= n5696;
    Ng4717 <= n5701_1;
    Ng1554 <= n5706_1;
    Ng3849 <= n5711;
    Pg17778 <= n5715_1;
    Ng3199 <= n5719_1;
    Ng5845 <= n5724_1;
    Ng4975 <= n5729;
    Ng790 <= n5734_1;
    Ng5913 <= n5739;
    Ng1902 <= n5744_1;
    Ng6163 <= n5749_1;
    Ng4125 <= n5754_1;
    Ng4821 <= n5759;
    Ng4939 <= n5764;
    Pg19334 <= n5769;
    Ng3207 <= n5773;
    Ng4483 <= n5777_1;
    Ng3259 <= n5782;
    Ng5142 <= n5787;
    Ng5248 <= n5792;
    Ng2126 <= n5797;
    Ng3694 <= n5802;
    Ng5481 <= n5807;
    Ng1964 <= n5812_1;
    Ng5097 <= n5817_1;
    Ng3215 <= n5822;
    Pg16748 <= n5826;
    Ng111 <= n5829_1;
    Ng4427 <= n5834;
    Ng2779 <= n5839;
    Pg8786 <= n5843_1;
    Pg7245 <= n5847_1;
    Ng1720 <= n5851;
    Ng1367 <= n5856;
    Ng5112 <= n5860_1;
    Ng4145 <= n5865_1;
    Ng2161 <= n5870_1;
    Ng376 <= n5875_1;
    Ng2361 <= n5880_1;
    Pg11447 <= n5885_1;
    Ng582 <= n5889;
    Ng2051 <= n5894_1;
    Ng1193 <= n5899;
    Ng2327 <= n5904;
    Ng907 <= n5909;
    Ng947 <= n5914;
    Ng1834 <= n5919_1;
    Ng3594 <= n5924_1;
    Ng2999 <= n5929;
    Ng2303 <= n5934;
    Pg17688 <= n5938_1;
    Ng699 <= n5942;
    Ng723 <= n5947_1;
    Ng5703 <= n5952_1;
    Ng546 <= n5957_1;
    Ng2472 <= n5962_1;
    Ng5953 <= n5967;
    Pg8277 <= n5972;
    Ng1740 <= n5976;
    Ng3550 <= n5981;
    Ng3845 <= n5986_1;
    Ng2116 <= n5991;
    Pg14635 <= n5995_1;
    Ng3195 <= n5999_1;
    Ng3913 <= n6004_1;
    Pg10306 <= n6009;
    Ng1687 <= n6013_1;
    Ng2681 <= n6018;
    Ng2533 <= n6023_1;
    Ng324 <= n6028;
    Ng2697 <= n6033_1;
    Ng4417 <= n6038;
    Ng6561 <= n6043_1;
    Ng1141 <= n6048_1;
    Pg12923 <= n6053;
    Ng2413 <= n6057_1;
    Ng1710 <= n6062_1;
    Ng6527 <= n6067;
    Ng3255 <= n6072_1;
    Ng1691 <= n6077_1;
    Ng2936 <= n6082_1;
    Ng5644 <= n6087;
    Ng5152 <= n6092_1;
    Ng5352 <= n6097_1;
    Pg8915 <= n6101;
    Ng2775 <= n6105_1;
    Ng2922 <= n6110;
    Ng1111 <= n6115_1;
    Ng5893 <= n6120_1;
    Pg16603 <= n6124_1;
    Ng6617 <= n6128_1;
    Ng2060 <= n6133_1;
    Ng4512 <= n6138;
    Ng5599 <= n6143;
    Ng3401 <= n6148;
    Ng4366 <= n6153;
    Pg16722 <= n6157;
    \[4433]  <= n6161;
    Ng3129 <= n6166;
    Ng3329 <= n6170;
    Ng5170 <= n6175;
    Ng26959 <= n6180;
    Ng5821 <= n6184;
    Ng6299 <= n6189;
    Pg8416 <= n6193;
    Ng2079 <= n6197;
    Ng4698 <= n6202;
    Ng3703 <= n6207_1;
    Ng1559 <= n6212;
    Ng943 <= n6217;
    Ng411 <= n6222;
    Pg9682 <= n6227;
    Ng3953 <= n6231;
    Ng2704 <= n6236;
    Ng6035 <= n6241;
    Ng1300 <= n6246;
    Ng4057 <= n6251_1;
    Ng5200 <= n6256_1;
    Ng4843 <= n6261_1;
    Ng5046 <= n6266;
    Ng2250 <= n6271;
    Ng26885 <= n6276;
    Ng4549 <= n6280;
    Ng2453 <= n6285;
    Ng5841 <= n6290_1;
    Pg14694 <= n6294;
    Ng2912 <= n6298;
    Ng2357 <= n6303;
    Pg8920 <= n6307;
    Ng164 <= n6311;
    Ng4253 <= n6316;
    Ng5016 <= n6321;
    Ng3119 <= n6326;
    Ng1351 <= n6331;
    Ng1648 <= n6336;
    Ng6972 <= n6341_1;
    Ng5115 <= n6345;
    Ng3352 <= n6350;
    Ng6657 <= n6355;
    Ng4552 <= n6360;
    Ng3893 <= n6365;
    Ng3211 <= n6370;
    Pg13049 <= n6374;
    Pg16624 <= n6377;
    Ng5595 <= n6381;
    Ng3614 <= n6386_1;
    Ng2894 <= n6391;
    Ng3125 <= n6396;
    Pg16686 <= n6400;
    Ng3821 <= n6404;
    Ng4141 <= n6409;
    Ng6974 <= n6414;
    Ng5272 <= n6418;
    Ng2735 <= n6423;
    Ng728 <= n6428;
    Ng6295 <= n6433;
    Ng2661 <= n6438;
    Ng1988 <= n6443;
    Ng5128 <= n6448;
    Ng1548 <= n6453;
    Ng3106 <= n6458;
    Ng4659 <= n6463;
    Ng4358 <= n6468;
    Ng1792 <= n6473;
    Ng2084 <= n6478;
    Ng3187 <= n6483;
    Ng4311 <= n6488;
    Ng2583 <= n6493;
    Ng3003 <= n6498;
    Ng1094 <= n6503;
    Ng3841 <= n6508;
    Ng4284 <= n6513;
    Ng3191 <= n6518;
    Ng4239 <= n6523;
    Ng4180 <= n6527;
    Ng691 <= n6532;
    Ng534 <= n6537;
    Ng385 <= n6542;
    Ng2004 <= n6547;
    Ng2527 <= n6552;
    Ng5456 <= n6556;
    Ng4420 <= n6561;
    Ng5148 <= n6566;
    Ng4507 <= n6571;
    Ng5348 <= n6576;
    Ng3223 <= n6581;
    Ng2970 <= n6586;
    Ng5698 <= n6591;
    Ng5260 <= n6596;
    Ng1521 <= n6601;
    Ng3522 <= n6606;
    Ng3115 <= n6611;
    Ng3251 <= n6616;
    Pg12832 <= n6621;
    Ng4628 <= n6625;
    Ng1996 <= n6630;
    Pg8342 <= n6635;
    Ng4515 <= n6639;
    Pg8787 <= n6643;
    Ng4300 <= n6647;
    Ng1724 <= n6652;
    Ng1379 <= n6657;
    Pg11388 <= n6662;
    Ng1878 <= n6666;
    Ng5619 <= n6671;
    Ng71 <= n6676;
    \[4437]  <= n6681;
  end
endmodule


