// Benchmark "mul9" written by ABC on Sat Apr 23 20:18:07 2016

module mul9 ( 
    a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7, b8, a8,
    z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15,
    z16, z17  );
  input  a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7,
    b8, a8;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15,
    z16, z17;
  wire n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n53,
    n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
    n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n634, n635, n636;
  assign z0 = a0 & b0;
  assign n38 = a0 & b1;
  assign n39 = b0 & a1;
  assign n40 = n38 & n39;
  assign n41 = ~n38 & ~n39;
  assign z1 = ~n40 & ~n41;
  assign n43 = a0 & b2;
  assign n44 = b0 & a2;
  assign n45 = b1 & a1;
  assign n46 = ~z0 & n45;
  assign n47 = n44 & ~n46;
  assign n48 = ~n44 & n46;
  assign n49 = ~n47 & ~n48;
  assign n50 = n43 & ~n49;
  assign n51 = ~n43 & n49;
  assign z2 = ~n50 & ~n51;
  assign n53 = a0 & b3;
  assign n54 = a1 & b2;
  assign n55 = n53 & n54;
  assign n56 = ~n53 & ~n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = b1 & a2;
  assign n59 = b0 & a3;
  assign n60 = n44 & n45;
  assign n61 = ~n40 & ~n60;
  assign n62 = n59 & ~n61;
  assign n63 = ~n59 & n61;
  assign n64 = ~n62 & ~n63;
  assign n65 = n58 & n64;
  assign n66 = ~n58 & ~n64;
  assign n67 = ~n65 & ~n66;
  assign n68 = n57 & n67;
  assign n69 = ~n57 & ~n67;
  assign n70 = ~n68 & ~n69;
  assign n71 = n50 & n70;
  assign n72 = ~n50 & ~n70;
  assign z3 = ~n71 & ~n72;
  assign n74 = ~n68 & ~n71;
  assign n75 = a0 & b4;
  assign n76 = b2 & a2;
  assign n77 = a1 & b3;
  assign n78 = ~n43 & n77;
  assign n79 = n76 & ~n78;
  assign n80 = ~n76 & n78;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~n75 & n81;
  assign n83 = n75 & ~n81;
  assign n84 = ~n82 & ~n83;
  assign n85 = b1 & a3;
  assign n86 = b0 & a4;
  assign n87 = ~n58 & ~n62;
  assign n88 = ~n63 & ~n87;
  assign n89 = n86 & n88;
  assign n90 = ~n86 & ~n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = ~n85 & ~n91;
  assign n93 = n85 & n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = ~n84 & ~n94;
  assign n96 = n84 & n94;
  assign n97 = ~n95 & ~n96;
  assign n98 = n74 & ~n97;
  assign n99 = ~n74 & n97;
  assign z4 = ~n98 & ~n99;
  assign n101 = ~n82 & n94;
  assign n102 = ~n83 & ~n101;
  assign n103 = a0 & b5;
  assign n104 = a1 & b4;
  assign n105 = n103 & n104;
  assign n106 = ~n103 & ~n104;
  assign n107 = ~n105 & ~n106;
  assign n108 = a2 & b3;
  assign n109 = b2 & a3;
  assign n110 = n76 & n77;
  assign n111 = ~n55 & ~n110;
  assign n112 = n109 & ~n111;
  assign n113 = ~n109 & n111;
  assign n114 = ~n112 & ~n113;
  assign n115 = n108 & n114;
  assign n116 = ~n108 & ~n114;
  assign n117 = ~n115 & ~n116;
  assign n118 = n107 & n117;
  assign n119 = ~n107 & ~n117;
  assign n120 = ~n118 & ~n119;
  assign n121 = b1 & a4;
  assign n122 = b0 & a5;
  assign n123 = ~n85 & ~n89;
  assign n124 = ~n90 & ~n123;
  assign n125 = n122 & n124;
  assign n126 = ~n122 & ~n124;
  assign n127 = ~n125 & ~n126;
  assign n128 = ~n121 & ~n127;
  assign n129 = n121 & n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = n120 & ~n130;
  assign n132 = ~n120 & n130;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n102 & ~n133;
  assign n135 = n102 & n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = n99 & n136;
  assign n138 = ~n99 & ~n136;
  assign z5 = ~n137 & ~n138;
  assign n140 = ~n134 & ~n137;
  assign n141 = ~n118 & ~n130;
  assign n142 = ~n119 & ~n141;
  assign n143 = a0 & b6;
  assign n144 = a2 & b4;
  assign n145 = a1 & b5;
  assign n146 = ~n75 & n145;
  assign n147 = n144 & ~n146;
  assign n148 = ~n144 & n146;
  assign n149 = ~n147 & ~n148;
  assign n150 = n143 & ~n149;
  assign n151 = ~n143 & n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = b3 & a3;
  assign n154 = b2 & a4;
  assign n155 = ~n108 & ~n112;
  assign n156 = ~n113 & ~n155;
  assign n157 = n154 & n156;
  assign n158 = ~n154 & ~n156;
  assign n159 = ~n157 & ~n158;
  assign n160 = ~n153 & ~n159;
  assign n161 = n153 & n159;
  assign n162 = ~n160 & ~n161;
  assign n163 = n152 & n162;
  assign n164 = ~n152 & ~n162;
  assign n165 = ~n163 & ~n164;
  assign n166 = b1 & a5;
  assign n167 = b0 & a6;
  assign n168 = ~n121 & ~n125;
  assign n169 = ~n126 & ~n168;
  assign n170 = n167 & n169;
  assign n171 = ~n167 & ~n169;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~n166 & ~n172;
  assign n174 = n166 & n172;
  assign n175 = ~n173 & ~n174;
  assign n176 = n165 & ~n175;
  assign n177 = ~n165 & n175;
  assign n178 = ~n176 & ~n177;
  assign n179 = n142 & ~n178;
  assign n180 = ~n142 & n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = n140 & ~n181;
  assign n183 = ~n140 & n181;
  assign z6 = ~n182 & ~n183;
  assign n185 = ~n179 & ~n183;
  assign n186 = ~n163 & ~n175;
  assign n187 = ~n164 & ~n186;
  assign n188 = a0 & b7;
  assign n189 = a1 & b6;
  assign n190 = n188 & n189;
  assign n191 = ~n188 & ~n189;
  assign n192 = ~n190 & ~n191;
  assign n193 = a2 & b5;
  assign n194 = a3 & b4;
  assign n195 = n144 & n145;
  assign n196 = ~n105 & ~n195;
  assign n197 = n194 & ~n196;
  assign n198 = ~n194 & n196;
  assign n199 = ~n197 & ~n198;
  assign n200 = n193 & n199;
  assign n201 = ~n193 & ~n199;
  assign n202 = ~n200 & ~n201;
  assign n203 = n192 & n202;
  assign n204 = ~n192 & ~n202;
  assign n205 = ~n203 & ~n204;
  assign n206 = n150 & n205;
  assign n207 = ~n150 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = b3 & a4;
  assign n210 = b2 & a5;
  assign n211 = ~n153 & ~n157;
  assign n212 = ~n158 & ~n211;
  assign n213 = n210 & n212;
  assign n214 = ~n210 & ~n212;
  assign n215 = ~n213 & ~n214;
  assign n216 = ~n209 & ~n215;
  assign n217 = n209 & n215;
  assign n218 = ~n216 & ~n217;
  assign n219 = n208 & n218;
  assign n220 = ~n208 & ~n218;
  assign n221 = ~n219 & ~n220;
  assign n222 = b1 & a6;
  assign n223 = b0 & a7;
  assign n224 = ~n166 & ~n170;
  assign n225 = ~n171 & ~n224;
  assign n226 = n223 & n225;
  assign n227 = ~n223 & ~n225;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n222 & ~n228;
  assign n230 = n222 & n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = n221 & ~n231;
  assign n233 = ~n221 & n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = n187 & ~n234;
  assign n236 = ~n187 & n234;
  assign n237 = ~n235 & ~n236;
  assign n238 = ~n185 & n237;
  assign n239 = n185 & ~n237;
  assign z7 = ~n238 & ~n239;
  assign n241 = ~n235 & ~n238;
  assign n242 = ~n219 & ~n231;
  assign n243 = ~n220 & ~n242;
  assign n244 = ~n203 & ~n206;
  assign n245 = a0 & b8;
  assign n246 = a2 & b6;
  assign n247 = a1 & b7;
  assign n248 = ~n143 & n247;
  assign n249 = n246 & ~n248;
  assign n250 = ~n246 & n248;
  assign n251 = ~n249 & ~n250;
  assign n252 = ~n245 & n251;
  assign n253 = n245 & ~n251;
  assign n254 = ~n252 & ~n253;
  assign n255 = a3 & b5;
  assign n256 = b4 & a4;
  assign n257 = ~n193 & ~n197;
  assign n258 = ~n198 & ~n257;
  assign n259 = n256 & n258;
  assign n260 = ~n256 & ~n258;
  assign n261 = ~n259 & ~n260;
  assign n262 = ~n255 & ~n261;
  assign n263 = n255 & n261;
  assign n264 = ~n262 & ~n263;
  assign n265 = ~n254 & ~n264;
  assign n266 = n254 & n264;
  assign n267 = ~n265 & ~n266;
  assign n268 = n244 & ~n267;
  assign n269 = ~n244 & n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = b3 & a5;
  assign n272 = b2 & a6;
  assign n273 = ~n209 & ~n213;
  assign n274 = ~n214 & ~n273;
  assign n275 = n272 & n274;
  assign n276 = ~n272 & ~n274;
  assign n277 = ~n275 & ~n276;
  assign n278 = ~n271 & ~n277;
  assign n279 = n271 & n277;
  assign n280 = ~n278 & ~n279;
  assign n281 = n270 & n280;
  assign n282 = ~n270 & ~n280;
  assign n283 = ~n281 & ~n282;
  assign n284 = b1 & a7;
  assign n285 = b0 & a8;
  assign n286 = ~n222 & ~n226;
  assign n287 = ~n227 & ~n286;
  assign n288 = n285 & n287;
  assign n289 = ~n285 & ~n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n284 & ~n290;
  assign n292 = n284 & n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = n283 & ~n293;
  assign n295 = ~n283 & n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = n243 & ~n296;
  assign n298 = ~n243 & n296;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~n241 & n299;
  assign n301 = n241 & ~n299;
  assign z8 = ~n300 & ~n301;
  assign n303 = ~n297 & ~n300;
  assign n304 = ~n282 & n293;
  assign n305 = ~n281 & ~n304;
  assign n306 = b1 & a8;
  assign n307 = ~n284 & ~n288;
  assign n308 = ~n289 & ~n307;
  assign n309 = n306 & n308;
  assign n310 = ~n306 & ~n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = a1 & b8;
  assign n313 = a2 & b7;
  assign n314 = a3 & b6;
  assign n315 = n246 & n247;
  assign n316 = ~n190 & ~n315;
  assign n317 = n314 & ~n316;
  assign n318 = ~n314 & n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = n313 & n319;
  assign n321 = ~n313 & ~n319;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n312 & ~n322;
  assign n324 = n312 & n322;
  assign n325 = ~n323 & ~n324;
  assign n326 = a4 & b5;
  assign n327 = b4 & a5;
  assign n328 = ~n255 & ~n259;
  assign n329 = ~n260 & ~n328;
  assign n330 = n327 & n329;
  assign n331 = ~n327 & ~n329;
  assign n332 = ~n330 & ~n331;
  assign n333 = ~n326 & ~n332;
  assign n334 = n326 & n332;
  assign n335 = ~n333 & ~n334;
  assign n336 = ~n325 & n335;
  assign n337 = n325 & ~n335;
  assign n338 = ~n336 & ~n337;
  assign n339 = ~n252 & n264;
  assign n340 = ~n253 & ~n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = n338 & n340;
  assign n343 = ~n341 & ~n342;
  assign n344 = n269 & n343;
  assign n345 = ~n269 & ~n343;
  assign n346 = ~n344 & ~n345;
  assign n347 = b3 & a6;
  assign n348 = b2 & a7;
  assign n349 = ~n271 & ~n275;
  assign n350 = ~n276 & ~n349;
  assign n351 = n348 & n350;
  assign n352 = ~n348 & ~n350;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n347 & ~n353;
  assign n355 = n347 & n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n346 & ~n356;
  assign n358 = n346 & n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n311 & ~n359;
  assign n361 = n311 & n359;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~n305 & n362;
  assign n364 = n305 & ~n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n303 & n365;
  assign n367 = n303 & ~n365;
  assign z9 = ~n366 & ~n367;
  assign n369 = ~n363 & ~n366;
  assign n370 = ~n341 & ~n344;
  assign n371 = a2 & b8;
  assign n372 = a3 & b7;
  assign n373 = a4 & b6;
  assign n374 = ~n313 & ~n317;
  assign n375 = ~n318 & ~n374;
  assign n376 = n373 & n375;
  assign n377 = ~n373 & ~n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = ~n372 & ~n378;
  assign n380 = n372 & n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = ~n371 & ~n381;
  assign n383 = n371 & n381;
  assign n384 = ~n382 & ~n383;
  assign n385 = b5 & a5;
  assign n386 = b4 & a6;
  assign n387 = ~n326 & ~n330;
  assign n388 = ~n331 & ~n387;
  assign n389 = n386 & n388;
  assign n390 = ~n386 & ~n388;
  assign n391 = ~n389 & ~n390;
  assign n392 = ~n385 & ~n391;
  assign n393 = n385 & n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n384 & n394;
  assign n396 = n384 & ~n394;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n323 & n335;
  assign n399 = ~n324 & ~n398;
  assign n400 = ~n397 & ~n399;
  assign n401 = n397 & n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n370 & n402;
  assign n404 = n370 & ~n402;
  assign n405 = ~n403 & ~n404;
  assign n406 = b3 & a7;
  assign n407 = b2 & a8;
  assign n408 = ~n347 & ~n351;
  assign n409 = ~n352 & ~n408;
  assign n410 = n407 & n409;
  assign n411 = ~n407 & ~n409;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n406 & ~n412;
  assign n414 = n406 & n412;
  assign n415 = ~n413 & ~n414;
  assign n416 = n309 & n415;
  assign n417 = ~n309 & ~n415;
  assign n418 = ~n416 & ~n417;
  assign n419 = n405 & n418;
  assign n420 = ~n405 & ~n418;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n311 & ~n358;
  assign n423 = ~n357 & ~n422;
  assign n424 = n421 & n423;
  assign n425 = ~n421 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n369 & n426;
  assign n428 = n369 & ~n426;
  assign z10 = ~n427 & ~n428;
  assign n430 = ~n424 & ~n427;
  assign n431 = ~n400 & ~n403;
  assign n432 = a3 & b8;
  assign n433 = a4 & b7;
  assign n434 = a5 & b6;
  assign n435 = ~n372 & ~n376;
  assign n436 = ~n377 & ~n435;
  assign n437 = n434 & n436;
  assign n438 = ~n434 & ~n436;
  assign n439 = ~n437 & ~n438;
  assign n440 = ~n433 & ~n439;
  assign n441 = n433 & n439;
  assign n442 = ~n440 & ~n441;
  assign n443 = n432 & n442;
  assign n444 = ~n432 & ~n442;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n383 & ~n394;
  assign n447 = ~n382 & ~n446;
  assign n448 = n445 & n447;
  assign n449 = ~n445 & ~n447;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~n431 & n450;
  assign n452 = n431 & ~n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = b3 & a8;
  assign n455 = ~n406 & ~n410;
  assign n456 = ~n411 & ~n455;
  assign n457 = n454 & n456;
  assign n458 = ~n454 & ~n456;
  assign n459 = ~n457 & ~n458;
  assign n460 = b5 & a6;
  assign n461 = b4 & a7;
  assign n462 = ~n385 & ~n389;
  assign n463 = ~n390 & ~n462;
  assign n464 = n461 & n463;
  assign n465 = ~n461 & ~n463;
  assign n466 = ~n464 & ~n465;
  assign n467 = ~n460 & ~n466;
  assign n468 = n460 & n466;
  assign n469 = ~n467 & ~n468;
  assign n470 = n459 & n469;
  assign n471 = ~n459 & ~n469;
  assign n472 = ~n470 & ~n471;
  assign n473 = ~n453 & ~n472;
  assign n474 = n453 & n472;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n405 & ~n416;
  assign n477 = ~n417 & ~n476;
  assign n478 = n475 & n477;
  assign n479 = ~n475 & ~n477;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n430 & n480;
  assign n482 = n430 & ~n480;
  assign z11 = ~n481 & ~n482;
  assign n484 = ~n478 & ~n481;
  assign n485 = ~n448 & ~n451;
  assign n486 = a4 & b8;
  assign n487 = a5 & b7;
  assign n488 = b6 & a6;
  assign n489 = ~n433 & ~n437;
  assign n490 = ~n438 & ~n489;
  assign n491 = n488 & n490;
  assign n492 = ~n488 & ~n490;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n487 & ~n493;
  assign n495 = n487 & n493;
  assign n496 = ~n494 & ~n495;
  assign n497 = n486 & n496;
  assign n498 = ~n486 & ~n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = n443 & n499;
  assign n501 = ~n443 & ~n499;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~n485 & n502;
  assign n504 = n485 & ~n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = b5 & a7;
  assign n507 = b4 & a8;
  assign n508 = ~n460 & ~n464;
  assign n509 = ~n465 & ~n508;
  assign n510 = n507 & n509;
  assign n511 = ~n507 & ~n509;
  assign n512 = ~n510 & ~n511;
  assign n513 = ~n506 & ~n512;
  assign n514 = n506 & n512;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n457 & ~n515;
  assign n517 = n457 & n515;
  assign n518 = ~n516 & ~n517;
  assign n519 = n505 & n518;
  assign n520 = ~n505 & ~n518;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~n453 & ~n470;
  assign n523 = ~n471 & ~n522;
  assign n524 = n521 & n523;
  assign n525 = ~n521 & ~n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = n484 & ~n526;
  assign n528 = ~n484 & n526;
  assign z12 = ~n527 & ~n528;
  assign n530 = ~n524 & ~n528;
  assign n531 = ~n500 & ~n503;
  assign n532 = b5 & a8;
  assign n533 = ~n506 & ~n510;
  assign n534 = ~n511 & ~n533;
  assign n535 = n532 & n534;
  assign n536 = ~n532 & ~n534;
  assign n537 = ~n535 & ~n536;
  assign n538 = n497 & n537;
  assign n539 = ~n497 & ~n537;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~n531 & n540;
  assign n542 = n531 & ~n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = a5 & b8;
  assign n545 = a6 & b7;
  assign n546 = b6 & a7;
  assign n547 = ~n487 & ~n491;
  assign n548 = ~n492 & ~n547;
  assign n549 = n546 & n548;
  assign n550 = ~n546 & ~n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n545 & ~n551;
  assign n553 = n545 & n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = n544 & n554;
  assign n556 = ~n544 & ~n554;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~n543 & ~n557;
  assign n559 = n543 & n557;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n505 & ~n517;
  assign n562 = ~n516 & ~n561;
  assign n563 = n560 & n562;
  assign n564 = ~n560 & ~n562;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n530 & n565;
  assign n567 = n530 & ~n565;
  assign z13 = ~n566 & ~n567;
  assign n569 = ~n563 & ~n566;
  assign n570 = ~n543 & ~n555;
  assign n571 = ~n556 & ~n570;
  assign n572 = ~n538 & ~n541;
  assign n573 = n535 & ~n572;
  assign n574 = ~n535 & n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = a6 & b8;
  assign n577 = b7 & a7;
  assign n578 = b6 & a8;
  assign n579 = ~n545 & ~n549;
  assign n580 = ~n550 & ~n579;
  assign n581 = n578 & n580;
  assign n582 = ~n578 & ~n580;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n577 & ~n583;
  assign n585 = n577 & n583;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n576 & ~n586;
  assign n588 = n576 & n586;
  assign n589 = ~n587 & ~n588;
  assign n590 = n575 & n589;
  assign n591 = ~n575 & ~n589;
  assign n592 = ~n590 & ~n591;
  assign n593 = n571 & n592;
  assign n594 = ~n571 & ~n592;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n569 & n595;
  assign n597 = n569 & ~n595;
  assign z14 = ~n596 & ~n597;
  assign n599 = ~n593 & ~n596;
  assign n600 = a7 & b8;
  assign n601 = b7 & a8;
  assign n602 = ~n577 & ~n581;
  assign n603 = ~n582 & ~n602;
  assign n604 = n601 & n603;
  assign n605 = ~n601 & ~n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = n600 & n606;
  assign n608 = ~n600 & ~n606;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n573 & ~n609;
  assign n611 = n573 & n609;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n575 & ~n588;
  assign n614 = ~n587 & ~n613;
  assign n615 = n612 & n614;
  assign n616 = ~n612 & ~n614;
  assign n617 = ~n615 & ~n616;
  assign n618 = n599 & ~n617;
  assign n619 = ~n599 & n617;
  assign z15 = ~n618 & ~n619;
  assign n621 = ~n615 & ~n619;
  assign n622 = b8 & n604;
  assign n623 = b8 & a8;
  assign n624 = ~n604 & ~n623;
  assign n625 = ~n622 & ~n624;
  assign n626 = ~n573 & ~n607;
  assign n627 = ~n608 & ~n626;
  assign n628 = n625 & n627;
  assign n629 = ~n625 & ~n627;
  assign n630 = ~n628 & ~n629;
  assign n631 = ~n621 & n630;
  assign n632 = n621 & ~n630;
  assign z16 = ~n631 & ~n632;
  assign n634 = n622 & n631;
  assign n635 = ~n622 & ~n628;
  assign n636 = ~n631 & n635;
  assign z17 = ~n634 & ~n636;
endmodule


