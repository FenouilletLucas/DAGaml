// Benchmark "alu4_cl" written by ABC on Tue May 16 16:07:44 2017

module alu4_cl ( 
    a, b, c, d, e, f, g, h, i, j,
    k, l, m, n, o, p  );
  input  a, b, c, d, e, f, g, h, i, j;
  output k, l, m, n, o, p;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n164, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339;
  assign n17 = a & c;
  assign n18 = c & ~n17;
  assign n19 = ~g & ~h;
  assign n20 = ~j & n19;
  assign n21 = g & j;
  assign n22 = ~n20 & ~n21;
  assign n23 = g & n22;
  assign n24 = e & ~f;
  assign n25 = g & ~h;
  assign n26 = ~e & f;
  assign n27 = e & f;
  assign n28 = h & n24;
  assign n29 = n23 & n28;
  assign n30 = j & n26;
  assign n31 = ~n25 & n30;
  assign n32 = n25 & n27;
  assign n33 = ~n31 & ~n32;
  assign n34 = ~n29 & n33;
  assign n35 = ~f & ~j;
  assign n36 = a & ~n17;
  assign n37 = ~n18 & ~n36;
  assign n38 = ~e & ~f;
  assign n39 = h & j;
  assign n40 = n17 & n39;
  assign n41 = ~g & n35;
  assign n42 = ~j & ~n22;
  assign n43 = ~n41 & ~n42;
  assign n44 = ~n27 & ~n38;
  assign n45 = ~n22 & n44;
  assign n46 = n34 & n45;
  assign n47 = n18 & n46;
  assign n48 = n22 & ~n24;
  assign n49 = n34 & n48;
  assign n50 = n40 & n49;
  assign n51 = n30 & n36;
  assign n52 = n17 & n38;
  assign n53 = n25 & n52;
  assign n54 = ~a & ~e;
  assign n55 = ~n43 & n54;
  assign n56 = a & n24;
  assign n57 = ~n22 & n56;
  assign n58 = ~c & ~n34;
  assign n59 = ~n57 & ~n58;
  assign n60 = ~n55 & n59;
  assign n61 = ~n53 & n60;
  assign n62 = ~n51 & n61;
  assign n63 = ~n50 & n62;
  assign n64 = ~n47 & n63;
  assign n65 = n22 & n25;
  assign n66 = ~g & n24;
  assign n67 = n23 & n38;
  assign n68 = ~n22 & n66;
  assign n69 = ~n67 & ~n68;
  assign n70 = h & ~n22;
  assign n71 = j & n38;
  assign n72 = n22 & n71;
  assign n73 = ~n27 & n70;
  assign n74 = ~n72 & ~n73;
  assign n75 = ~n22 & n25;
  assign n76 = n22 & n27;
  assign n77 = n39 & n76;
  assign n78 = n26 & n75;
  assign n79 = ~n77 & ~n78;
  assign n80 = n26 & n39;
  assign n81 = j & n25;
  assign n82 = n24 & n81;
  assign n83 = a & ~n64;
  assign n84 = n27 & n81;
  assign n85 = n83 & n84;
  assign n86 = n38 & n64;
  assign n87 = n81 & n86;
  assign n88 = n17 & n82;
  assign n89 = ~n80 & ~n88;
  assign n90 = ~n87 & n89;
  assign n91 = ~n85 & n90;
  assign n92 = n82 & n91;
  assign n93 = ~g & n17;
  assign n94 = n80 & n93;
  assign n95 = ~n92 & ~n94;
  assign n96 = n24 & n75;
  assign n97 = ~n64 & n96;
  assign n98 = ~h & j;
  assign n99 = ~n25 & n98;
  assign n100 = j & ~n64;
  assign n101 = ~n27 & n100;
  assign n102 = n95 & n101;
  assign n103 = n79 & n102;
  assign n104 = n74 & n103;
  assign n105 = n75 & n79;
  assign n106 = ~n97 & n105;
  assign n107 = ~n36 & n106;
  assign n108 = j & n22;
  assign n109 = n36 & n108;
  assign n110 = ~a & n27;
  assign n111 = n70 & n110;
  assign n112 = ~a & ~n64;
  assign n113 = n70 & n112;
  assign n114 = a & n64;
  assign n115 = ~n74 & n114;
  assign n116 = j & n66;
  assign n117 = n18 & n116;
  assign n118 = a & n99;
  assign n119 = n64 & ~n79;
  assign n120 = ~n118 & ~n119;
  assign n121 = ~n117 & n120;
  assign n122 = ~n115 & n121;
  assign n123 = ~n113 & n122;
  assign n124 = ~n111 & n123;
  assign n125 = ~n109 & n124;
  assign n126 = ~n107 & n125;
  assign n127 = ~n104 & n126;
  assign n128 = n27 & n99;
  assign n129 = h & ~j;
  assign n130 = ~n27 & n129;
  assign n131 = n34 & n130;
  assign n132 = n18 & n131;
  assign n133 = ~j & ~n64;
  assign n134 = ~n37 & n133;
  assign n135 = ~n35 & n134;
  assign n136 = n17 & n129;
  assign n137 = ~n24 & n136;
  assign n138 = n22 & n35;
  assign n139 = n36 & n138;
  assign n140 = a & ~n65;
  assign n141 = n23 & n140;
  assign n142 = ~c & n65;
  assign n143 = n35 & n142;
  assign n144 = ~n64 & n69;
  assign n145 = n35 & n144;
  assign n146 = n26 & n37;
  assign n147 = n65 & n146;
  assign n148 = ~i & j;
  assign n149 = n127 & n148;
  assign n150 = n64 & ~n69;
  assign n151 = i & ~n127;
  assign n152 = ~n128 & ~n151;
  assign n153 = ~n150 & n152;
  assign n154 = ~n149 & n153;
  assign n155 = ~n147 & n154;
  assign n156 = ~n145 & n155;
  assign n157 = ~n143 & n156;
  assign n158 = ~n141 & n157;
  assign n159 = ~n139 & n158;
  assign n160 = ~n137 & n159;
  assign n161 = ~n135 & n160;
  assign k = n132 | ~n161;
  assign n = b & d;
  assign n164 = ~b & ~d;
  assign m = n | n164;
  assign n166 = ~d & m;
  assign n167 = ~n24 & n;
  assign n168 = n34 & n167;
  assign n169 = n39 & n168;
  assign n170 = ~n70 & n169;
  assign n171 = n26 & m;
  assign n172 = n18 & n171;
  assign n173 = n81 & n172;
  assign n174 = n26 & ~m;
  assign n175 = ~n18 & n174;
  assign n176 = n81 & n175;
  assign n177 = ~n22 & n24;
  assign n178 = ~n166 & n177;
  assign n179 = a & n38;
  assign n180 = n70 & n179;
  assign n181 = n38 & n;
  assign n182 = n25 & n181;
  assign n183 = ~b & ~e;
  assign n184 = ~n43 & n183;
  assign n185 = ~d & ~n34;
  assign n186 = ~n184 & ~n185;
  assign n187 = ~n182 & n186;
  assign n188 = ~n180 & n187;
  assign n189 = ~n178 & n188;
  assign n190 = ~n176 & n189;
  assign n191 = ~n173 & n190;
  assign n192 = ~n170 & n191;
  assign n193 = n66 & ~m;
  assign n194 = ~i & ~n127;
  assign n195 = a & ~n91;
  assign n196 = b & ~n192;
  assign n197 = n27 & n196;
  assign n198 = n81 & n197;
  assign n199 = n38 & n192;
  assign n200 = n81 & n199;
  assign n201 = n82 & n;
  assign n202 = n80 & ~n192;
  assign n203 = b & n80;
  assign n204 = ~n202 & ~n203;
  assign n205 = ~n201 & n204;
  assign n206 = ~n200 & n205;
  assign n207 = ~n198 & n206;
  assign n208 = ~a & ~b;
  assign n209 = n70 & n208;
  assign n210 = n91 & n207;
  assign n211 = n75 & n210;
  assign n212 = ~n209 & ~n211;
  assign n213 = n82 & n207;
  assign n214 = ~g & n;
  assign n215 = n80 & n214;
  assign n216 = ~n213 & ~n215;
  assign n217 = n192 & ~n216;
  assign n218 = ~n192 & n216;
  assign n219 = ~n217 & ~n218;
  assign n220 = ~n83 & n192;
  assign n221 = n83 & ~n192;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~b & ~n207;
  assign n224 = b & n207;
  assign n225 = ~n223 & ~n224;
  assign n226 = n64 & ~n222;
  assign n227 = n22 & n80;
  assign n228 = n207 & ~n216;
  assign n229 = ~n207 & n216;
  assign n230 = ~n228 & ~n229;
  assign n231 = n100 & ~n192;
  assign n232 = n207 & n231;
  assign n233 = ~n70 & n232;
  assign n234 = ~n195 & n233;
  assign n235 = n44 & n95;
  assign n236 = ~n219 & n235;
  assign n237 = n212 & n236;
  assign n238 = n98 & n237;
  assign n239 = a & b;
  assign n240 = j & n239;
  assign n241 = ~n222 & n240;
  assign n242 = ~n22 & n241;
  assign n243 = ~n96 & n242;
  assign n244 = n79 & ~n225;
  assign n245 = ~n96 & n244;
  assign n246 = n98 & n245;
  assign n247 = ~n195 & n246;
  assign n248 = n22 & ~n193;
  assign n249 = n226 & n248;
  assign n250 = n40 & n249;
  assign n251 = j & n193;
  assign n252 = ~n40 & n251;
  assign n253 = n95 & ~n230;
  assign n254 = n227 & n253;
  assign n255 = n64 & ~n219;
  assign n256 = n96 & n255;
  assign n257 = ~b & n222;
  assign n258 = ~n74 & n257;
  assign n259 = b & ~n222;
  assign n260 = ~n74 & n259;
  assign n261 = ~n79 & n226;
  assign n262 = n27 & ~n212;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n260 & n263;
  assign n265 = ~n258 & n264;
  assign n266 = ~n256 & n265;
  assign n267 = ~n254 & n266;
  assign n268 = ~n252 & n267;
  assign n269 = ~n250 & n268;
  assign n270 = ~n247 & n269;
  assign n271 = ~n243 & n270;
  assign n272 = ~n238 & n271;
  assign n273 = ~n234 & n272;
  assign n274 = ~j & ~m;
  assign n275 = ~n192 & n274;
  assign n276 = ~n35 & n275;
  assign n277 = n129 & n;
  assign n278 = n43 & n277;
  assign n279 = d & h;
  assign n280 = ~j & n279;
  assign n281 = n26 & n280;
  assign n282 = b & ~n65;
  assign n283 = n23 & n282;
  assign n284 = ~d & n65;
  assign n285 = n35 & n284;
  assign n286 = n22 & n193;
  assign n287 = n35 & n286;
  assign n288 = n69 & ~n192;
  assign n289 = n35 & n288;
  assign n290 = n65 & n171;
  assign n291 = h & n38;
  assign n292 = ~n43 & n291;
  assign n293 = n194 & n273;
  assign n294 = ~n194 & ~n273;
  assign n295 = ~n69 & n192;
  assign n296 = ~n128 & ~n295;
  assign n297 = ~n294 & n296;
  assign n298 = ~n293 & n297;
  assign n299 = ~n292 & n298;
  assign n300 = ~n290 & n299;
  assign n301 = ~n289 & n300;
  assign n302 = ~n287 & n301;
  assign n303 = ~n285 & n302;
  assign n304 = ~n283 & n303;
  assign n305 = ~n281 & n304;
  assign n306 = ~n278 & n305;
  assign l = n276 | ~n306;
  assign n308 = ~n95 & n227;
  assign n309 = ~n179 & ~n308;
  assign n310 = ~n27 & ~n192;
  assign n311 = ~n222 & n310;
  assign n312 = n39 & n311;
  assign n313 = ~n227 & n312;
  assign n314 = j & n27;
  assign n315 = n22 & n314;
  assign n316 = n226 & n315;
  assign n317 = ~n27 & n;
  assign n318 = n22 & n317;
  assign n319 = n39 & n318;
  assign n320 = b & n273;
  assign n321 = ~n27 & n320;
  assign n322 = n39 & n321;
  assign n323 = n78 & n226;
  assign n324 = ~n207 & ~n309;
  assign n325 = n195 & n324;
  assign n326 = ~f & n273;
  assign n327 = n75 & n326;
  assign n328 = n40 & n193;
  assign n329 = n194 & ~n273;
  assign n330 = ~n192 & ~n216;
  assign n331 = ~n262 & ~n330;
  assign n332 = ~n329 & n331;
  assign n333 = ~n328 & n332;
  assign n334 = ~n327 & n333;
  assign n335 = ~n325 & n334;
  assign n336 = ~n323 & n335;
  assign n337 = ~n322 & n336;
  assign n338 = ~n319 & n337;
  assign n339 = ~n316 & n338;
  assign o = n313 | ~n339;
  assign p = n37 & m;
endmodule


