// Benchmark "i2" written by ABC on Tue May 16 16:07:50 2017

module i2 ( 
    \V126(17) , \V144(21) , \V30(29) , \V126(1) , \V126(16) , \V144(20) ,
    \V30(28) , \V126(0) , \V126(19) , \V144(23) , \V126(18) , \V144(22) ,
    \V62(13) , \V144(25) , \V62(12) , \V191(31) , \V144(24) , \V62(15) ,
    \V94(31) , \V62(14) , \V126(7) , \V94(30) , \V126(6) , \V144(19) ,
    \V30(31) , \V201(3) , \V126(9) , \V144(18) , \V62(11) , \V30(30) ,
    \V201(2) , \V126(8) , \V126(11) , \V62(10) , \V201(5) , \V126(10) ,
    \V201(4) , \V126(13) , \V176(31) , \V126(12) , \V176(30) , \V94(2) ,
    \V126(15) , \V63(0) , \V201(1) , \V94(3) , \V126(14) , \V62(17) ,
    \V201(0) , \V94(4) , \V193(1) , \V62(16) , \V94(5) , \V193(0) ,
    \V62(19) , \V94(6) , \V62(18) , \V176(3) , \V94(7) , \V62(23) ,
    \V176(2) , \V94(8) , \V129(0) , \V62(22) , \V176(5) , \V201(7) ,
    \V94(9) , \V62(25) , \V176(4) , \V201(6) , \V62(24) , \V176(27) ,
    \V176(26) , \V176(1) , \V176(29) , \V62(21) , \V176(0) , \V176(28) ,
    \V62(20) , \V188(31) , \V176(7) , \V62(0) , \V188(30) , \V62(27) ,
    \V176(6) , \V62(1) , \V62(26) , \V176(9) , \V176(21) , \V62(2) ,
    \V62(29) , \V176(8) , \V176(20) , \V62(3) , \V62(28) , \V176(23) ,
    \V62(4) , \V176(22) , \V62(5) , \V94(13) , \V128(0) , \V176(25) ,
    \V62(6) , \V94(12) , \V176(24) , \V62(7) , \V94(15) , \V30(13) ,
    \V130(0) , \V176(17) , \V62(8) , \V94(14) , \V30(12) , \V176(16) ,
    \V62(9) , \V188(27) , \V30(15) , \V176(19) , \V188(26) , \V62(31) ,
    \V30(14) , \V126(31) , \V176(18) , \V94(11) , \V188(29) , \V62(30) ,
    \V126(30) , \V94(10) , \V188(28) , \V30(11) , \V30(10) , \V144(31) ,
    \V94(17) , \V176(11) , \V144(30) , \V94(16) , \V176(10) , \V94(19) ,
    \V30(17) , \V176(13) , \V94(18) , \V30(16) , \V176(12) , \V126(27) ,
    \V94(23) , \V188(23) , \V30(2) , \V30(19) , \V176(15) , \V126(26) ,
    \V94(22) , \V188(22) , \V30(3) , \V127(0) , \V30(18) , \V176(14) ,
    \V126(29) , \V94(25) , \V188(25) , \V30(4) , \V30(23) , \V126(28) ,
    \V94(24) , \V188(24) , \V30(5) , \V30(22) , \V30(6) , \V30(25) ,
    \V30(7) , \V30(24) , \V144(27) , \V94(21) , \V30(8) , \V144(26) ,
    \V94(20) , \V30(9) , \V178(1) , \V144(29) , \V178(0) , \V30(21) ,
    \V144(28) , \V30(20) , \V126(21) , \V126(3) , \V126(20) , \V126(2) ,
    \V126(23) , \V94(27) , \V126(5) , \V126(22) , \V94(26) , \V64(0) ,
    \V126(4) , \V126(25) , \V94(29) , \V190(1) , \V30(27) , \V126(24) ,
    \V94(28) , \V190(0) , \V30(26) ,
    \V202(0)   );
  input  \V126(17) , \V144(21) , \V30(29) , \V126(1) , \V126(16) ,
    \V144(20) , \V30(28) , \V126(0) , \V126(19) , \V144(23) , \V126(18) ,
    \V144(22) , \V62(13) , \V144(25) , \V62(12) , \V191(31) , \V144(24) ,
    \V62(15) , \V94(31) , \V62(14) , \V126(7) , \V94(30) , \V126(6) ,
    \V144(19) , \V30(31) , \V201(3) , \V126(9) , \V144(18) , \V62(11) ,
    \V30(30) , \V201(2) , \V126(8) , \V126(11) , \V62(10) , \V201(5) ,
    \V126(10) , \V201(4) , \V126(13) , \V176(31) , \V126(12) , \V176(30) ,
    \V94(2) , \V126(15) , \V63(0) , \V201(1) , \V94(3) , \V126(14) ,
    \V62(17) , \V201(0) , \V94(4) , \V193(1) , \V62(16) , \V94(5) ,
    \V193(0) , \V62(19) , \V94(6) , \V62(18) , \V176(3) , \V94(7) ,
    \V62(23) , \V176(2) , \V94(8) , \V129(0) , \V62(22) , \V176(5) ,
    \V201(7) , \V94(9) , \V62(25) , \V176(4) , \V201(6) , \V62(24) ,
    \V176(27) , \V176(26) , \V176(1) , \V176(29) , \V62(21) , \V176(0) ,
    \V176(28) , \V62(20) , \V188(31) , \V176(7) , \V62(0) , \V188(30) ,
    \V62(27) , \V176(6) , \V62(1) , \V62(26) , \V176(9) , \V176(21) ,
    \V62(2) , \V62(29) , \V176(8) , \V176(20) , \V62(3) , \V62(28) ,
    \V176(23) , \V62(4) , \V176(22) , \V62(5) , \V94(13) , \V128(0) ,
    \V176(25) , \V62(6) , \V94(12) , \V176(24) , \V62(7) , \V94(15) ,
    \V30(13) , \V130(0) , \V176(17) , \V62(8) , \V94(14) , \V30(12) ,
    \V176(16) , \V62(9) , \V188(27) , \V30(15) , \V176(19) , \V188(26) ,
    \V62(31) , \V30(14) , \V126(31) , \V176(18) , \V94(11) , \V188(29) ,
    \V62(30) , \V126(30) , \V94(10) , \V188(28) , \V30(11) , \V30(10) ,
    \V144(31) , \V94(17) , \V176(11) , \V144(30) , \V94(16) , \V176(10) ,
    \V94(19) , \V30(17) , \V176(13) , \V94(18) , \V30(16) , \V176(12) ,
    \V126(27) , \V94(23) , \V188(23) , \V30(2) , \V30(19) , \V176(15) ,
    \V126(26) , \V94(22) , \V188(22) , \V30(3) , \V127(0) , \V30(18) ,
    \V176(14) , \V126(29) , \V94(25) , \V188(25) , \V30(4) , \V30(23) ,
    \V126(28) , \V94(24) , \V188(24) , \V30(5) , \V30(22) , \V30(6) ,
    \V30(25) , \V30(7) , \V30(24) , \V144(27) , \V94(21) , \V30(8) ,
    \V144(26) , \V94(20) , \V30(9) , \V178(1) , \V144(29) , \V178(0) ,
    \V30(21) , \V144(28) , \V30(20) , \V126(21) , \V126(3) , \V126(20) ,
    \V126(2) , \V126(23) , \V94(27) , \V126(5) , \V126(22) , \V94(26) ,
    \V64(0) , \V126(4) , \V126(25) , \V94(29) , \V190(1) , \V30(27) ,
    \V126(24) , \V94(28) , \V190(0) , \V30(26) ;
  output \V202(0) ;
  wire n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732;
  assign n203 = ~\V176(31)  & ~\V178(1) ;
  assign n204 = ~\V176(29)  & n203;
  assign n205 = ~\V176(27)  & n204;
  assign n206 = ~\V176(25)  & n205;
  assign n207 = ~\V176(23)  & n206;
  assign n208 = ~\V176(21)  & n207;
  assign n209 = ~\V176(19)  & n208;
  assign n210 = ~\V176(18)  & n209;
  assign n211 = ~\V176(20)  & n210;
  assign n212 = ~\V176(22)  & n211;
  assign n213 = ~\V176(24)  & n212;
  assign n214 = ~\V176(26)  & n213;
  assign n215 = ~\V176(28)  & n214;
  assign n216 = ~\V176(30)  & n215;
  assign n217 = ~\V178(0)  & n216;
  assign n218 = \V191(31)  & \V201(7) ;
  assign n219 = \V201(6)  & n218;
  assign n220 = \V201(5)  & \V188(24) ;
  assign n221 = \V201(4)  & n220;
  assign n222 = \V201(5)  & \V188(22) ;
  assign n223 = \V201(4)  & n222;
  assign n224 = \V201(5)  & \V188(23) ;
  assign n225 = \V201(4)  & n224;
  assign n226 = \V201(5)  & \V188(25) ;
  assign n227 = \V201(4)  & n226;
  assign n228 = \V201(3)  & \V176(0) ;
  assign n229 = \V201(2)  & n228;
  assign n230 = \V201(3)  & \V144(30) ;
  assign n231 = \V201(2)  & n230;
  assign n232 = \V201(3)  & \V144(28) ;
  assign n233 = \V201(2)  & n232;
  assign n234 = \V201(3)  & \V144(26) ;
  assign n235 = \V201(2)  & n234;
  assign n236 = \V144(24)  & \V201(3) ;
  assign n237 = \V201(2)  & n236;
  assign n238 = \V144(22)  & \V201(3) ;
  assign n239 = \V201(2)  & n238;
  assign n240 = \V144(20)  & \V201(3) ;
  assign n241 = \V201(2)  & n240;
  assign n242 = \V201(3)  & \V144(18) ;
  assign n243 = \V201(2)  & n242;
  assign n244 = \V144(19)  & \V201(3) ;
  assign n245 = \V201(2)  & n244;
  assign n246 = \V144(21)  & \V201(3) ;
  assign n247 = \V201(2)  & n246;
  assign n248 = \V144(23)  & \V201(3) ;
  assign n249 = \V201(2)  & n248;
  assign n250 = \V144(25)  & \V201(3) ;
  assign n251 = \V201(2)  & n250;
  assign n252 = \V201(3)  & \V144(27) ;
  assign n253 = \V201(2)  & n252;
  assign n254 = \V201(3)  & \V144(29) ;
  assign n255 = \V201(2)  & n254;
  assign n256 = \V201(3)  & \V144(31) ;
  assign n257 = \V201(2)  & n256;
  assign n258 = \V201(3)  & \V176(1) ;
  assign n259 = \V201(2)  & n258;
  assign n260 = \V63(0)  & ~\V201(0) ;
  assign n261 = \V201(1)  & n260;
  assign n262 = ~\V201(0)  & \V62(30) ;
  assign n263 = \V201(1)  & n262;
  assign n264 = ~\V201(0)  & \V62(28) ;
  assign n265 = \V201(1)  & n264;
  assign n266 = ~\V201(0)  & \V62(26) ;
  assign n267 = \V201(1)  & n266;
  assign n268 = ~\V201(0)  & \V62(24) ;
  assign n269 = \V201(1)  & n268;
  assign n270 = ~\V201(0)  & \V62(22) ;
  assign n271 = \V201(1)  & n270;
  assign n272 = ~\V201(0)  & \V62(20) ;
  assign n273 = \V201(1)  & n272;
  assign n274 = ~\V201(0)  & \V62(18) ;
  assign n275 = \V201(1)  & n274;
  assign n276 = ~\V201(0)  & \V62(16) ;
  assign n277 = \V201(1)  & n276;
  assign n278 = \V62(14)  & ~\V201(0) ;
  assign n279 = \V201(1)  & n278;
  assign n280 = \V62(12)  & ~\V201(0) ;
  assign n281 = \V201(1)  & n280;
  assign n282 = \V62(10)  & ~\V201(0) ;
  assign n283 = \V201(1)  & n282;
  assign n284 = ~\V201(0)  & \V62(8) ;
  assign n285 = \V201(1)  & n284;
  assign n286 = ~\V201(0)  & \V62(6) ;
  assign n287 = \V201(1)  & n286;
  assign n288 = ~\V201(0)  & \V62(4) ;
  assign n289 = \V201(1)  & n288;
  assign n290 = ~\V201(0)  & \V62(2) ;
  assign n291 = \V201(1)  & n290;
  assign n292 = ~\V201(0)  & \V62(3) ;
  assign n293 = \V201(1)  & n292;
  assign n294 = ~\V201(0)  & \V62(5) ;
  assign n295 = \V201(1)  & n294;
  assign n296 = ~\V201(0)  & \V62(7) ;
  assign n297 = \V201(1)  & n296;
  assign n298 = ~\V201(0)  & \V62(9) ;
  assign n299 = \V201(1)  & n298;
  assign n300 = \V62(11)  & ~\V201(0) ;
  assign n301 = \V201(1)  & n300;
  assign n302 = \V62(13)  & ~\V201(0) ;
  assign n303 = \V201(1)  & n302;
  assign n304 = \V62(15)  & ~\V201(0) ;
  assign n305 = \V201(1)  & n304;
  assign n306 = \V62(17)  & ~\V201(0) ;
  assign n307 = \V201(1)  & n306;
  assign n308 = ~\V201(0)  & \V62(19) ;
  assign n309 = \V201(1)  & n308;
  assign n310 = ~\V201(0)  & \V62(21) ;
  assign n311 = \V201(1)  & n310;
  assign n312 = ~\V201(0)  & \V62(23) ;
  assign n313 = \V201(1)  & n312;
  assign n314 = ~\V201(0)  & \V62(25) ;
  assign n315 = \V201(1)  & n314;
  assign n316 = ~\V201(0)  & \V62(27) ;
  assign n317 = \V201(1)  & n316;
  assign n318 = ~\V201(0)  & \V62(29) ;
  assign n319 = \V201(1)  & n318;
  assign n320 = ~\V201(0)  & \V62(31) ;
  assign n321 = \V201(1)  & n320;
  assign n322 = ~\V201(0)  & \V64(0) ;
  assign n323 = \V201(1)  & n322;
  assign n324 = ~\V201(0)  & \V62(0) ;
  assign n325 = \V201(1)  & n324;
  assign n326 = \V30(30)  & ~\V201(0) ;
  assign n327 = \V201(1)  & n326;
  assign n328 = \V30(28)  & ~\V201(0) ;
  assign n329 = \V201(1)  & n328;
  assign n330 = ~\V201(0)  & \V30(26) ;
  assign n331 = \V201(1)  & n330;
  assign n332 = ~\V201(0)  & \V30(24) ;
  assign n333 = \V201(1)  & n332;
  assign n334 = ~\V201(0)  & \V30(22) ;
  assign n335 = \V201(1)  & n334;
  assign n336 = ~\V201(0)  & \V30(20) ;
  assign n337 = \V201(1)  & n336;
  assign n338 = ~\V201(0)  & \V30(18) ;
  assign n339 = \V201(1)  & n338;
  assign n340 = ~\V201(0)  & \V30(16) ;
  assign n341 = \V201(1)  & n340;
  assign n342 = ~\V201(0)  & \V30(14) ;
  assign n343 = \V201(1)  & n342;
  assign n344 = ~\V201(0)  & \V30(12) ;
  assign n345 = \V201(1)  & n344;
  assign n346 = ~\V201(0)  & \V30(10) ;
  assign n347 = \V201(1)  & n346;
  assign n348 = ~\V201(0)  & \V30(8) ;
  assign n349 = \V201(1)  & n348;
  assign n350 = ~\V201(0)  & \V30(6) ;
  assign n351 = \V201(1)  & n350;
  assign n352 = ~\V201(0)  & \V30(4) ;
  assign n353 = \V201(1)  & n352;
  assign n354 = ~\V201(0)  & \V30(2) ;
  assign n355 = \V201(1)  & n354;
  assign n356 = ~\V201(0)  & \V30(3) ;
  assign n357 = \V201(1)  & n356;
  assign n358 = ~\V201(0)  & \V30(5) ;
  assign n359 = \V201(1)  & n358;
  assign n360 = ~\V201(0)  & \V30(7) ;
  assign n361 = \V201(1)  & n360;
  assign n362 = ~\V201(0)  & \V30(9) ;
  assign n363 = \V201(1)  & n362;
  assign n364 = ~\V201(0)  & \V30(11) ;
  assign n365 = \V201(1)  & n364;
  assign n366 = ~\V201(0)  & \V30(13) ;
  assign n367 = \V201(1)  & n366;
  assign n368 = ~\V201(0)  & \V30(15) ;
  assign n369 = \V201(1)  & n368;
  assign n370 = ~\V201(0)  & \V30(17) ;
  assign n371 = \V201(1)  & n370;
  assign n372 = ~\V201(0)  & \V30(19) ;
  assign n373 = \V201(1)  & n372;
  assign n374 = ~\V201(0)  & \V30(21) ;
  assign n375 = \V201(1)  & n374;
  assign n376 = ~\V201(0)  & \V30(23) ;
  assign n377 = \V201(1)  & n376;
  assign n378 = ~\V201(0)  & \V30(25) ;
  assign n379 = \V201(1)  & n378;
  assign n380 = ~\V201(0)  & \V30(27) ;
  assign n381 = \V201(1)  & n380;
  assign n382 = \V30(29)  & ~\V201(0) ;
  assign n383 = \V201(1)  & n382;
  assign n384 = \V30(31)  & ~\V201(0) ;
  assign n385 = \V201(1)  & n384;
  assign n386 = ~\V201(0)  & \V62(1) ;
  assign n387 = \V201(1)  & n386;
  assign n388 = \V201(0)  & \V127(0) ;
  assign n389 = \V201(1)  & n388;
  assign n390 = \V201(0)  & \V126(30) ;
  assign n391 = \V201(1)  & n390;
  assign n392 = \V201(0)  & \V126(28) ;
  assign n393 = \V201(1)  & n392;
  assign n394 = \V201(0)  & \V126(26) ;
  assign n395 = \V201(1)  & n394;
  assign n396 = \V201(0)  & \V126(24) ;
  assign n397 = \V201(1)  & n396;
  assign n398 = \V201(0)  & \V126(22) ;
  assign n399 = \V201(1)  & n398;
  assign n400 = \V201(0)  & \V126(20) ;
  assign n401 = \V201(1)  & n400;
  assign n402 = \V126(18)  & \V201(0) ;
  assign n403 = \V201(1)  & n402;
  assign n404 = \V126(16)  & \V201(0) ;
  assign n405 = \V201(1)  & n404;
  assign n406 = \V126(14)  & \V201(0) ;
  assign n407 = \V201(1)  & n406;
  assign n408 = \V126(12)  & \V201(0) ;
  assign n409 = \V201(1)  & n408;
  assign n410 = \V126(10)  & \V201(0) ;
  assign n411 = \V201(1)  & n410;
  assign n412 = \V126(8)  & \V201(0) ;
  assign n413 = \V201(1)  & n412;
  assign n414 = \V126(6)  & \V201(0) ;
  assign n415 = \V201(1)  & n414;
  assign n416 = \V201(0)  & \V126(4) ;
  assign n417 = \V201(1)  & n416;
  assign n418 = \V201(0)  & \V126(2) ;
  assign n419 = \V201(1)  & n418;
  assign n420 = \V201(0)  & \V126(3) ;
  assign n421 = \V201(1)  & n420;
  assign n422 = \V201(0)  & \V126(5) ;
  assign n423 = \V201(1)  & n422;
  assign n424 = \V126(7)  & \V201(0) ;
  assign n425 = \V201(1)  & n424;
  assign n426 = \V126(9)  & \V201(0) ;
  assign n427 = \V201(1)  & n426;
  assign n428 = \V126(11)  & \V201(0) ;
  assign n429 = \V201(1)  & n428;
  assign n430 = \V126(13)  & \V201(0) ;
  assign n431 = \V201(1)  & n430;
  assign n432 = \V126(15)  & \V201(0) ;
  assign n433 = \V201(1)  & n432;
  assign n434 = \V126(17)  & \V201(0) ;
  assign n435 = \V201(1)  & n434;
  assign n436 = \V126(19)  & \V201(0) ;
  assign n437 = \V201(1)  & n436;
  assign n438 = \V201(0)  & \V126(21) ;
  assign n439 = \V201(1)  & n438;
  assign n440 = \V201(0)  & \V126(23) ;
  assign n441 = \V201(1)  & n440;
  assign n442 = \V201(0)  & \V126(25) ;
  assign n443 = \V201(1)  & n442;
  assign n444 = \V201(0)  & \V126(27) ;
  assign n445 = \V201(1)  & n444;
  assign n446 = \V201(0)  & \V126(29) ;
  assign n447 = \V201(1)  & n446;
  assign n448 = \V201(0)  & \V126(31) ;
  assign n449 = \V201(1)  & n448;
  assign n450 = \V201(0)  & \V128(0) ;
  assign n451 = \V201(1)  & n450;
  assign n452 = \V126(0)  & \V201(0) ;
  assign n453 = \V201(1)  & n452;
  assign n454 = \V94(30)  & \V201(0) ;
  assign n455 = \V201(1)  & n454;
  assign n456 = \V201(0)  & \V94(28) ;
  assign n457 = \V201(1)  & n456;
  assign n458 = \V201(0)  & \V94(26) ;
  assign n459 = \V201(1)  & n458;
  assign n460 = \V201(0)  & \V94(24) ;
  assign n461 = \V201(1)  & n460;
  assign n462 = \V201(0)  & \V94(22) ;
  assign n463 = \V201(1)  & n462;
  assign n464 = \V201(0)  & \V94(20) ;
  assign n465 = \V201(1)  & n464;
  assign n466 = \V201(0)  & \V94(18) ;
  assign n467 = \V201(1)  & n466;
  assign n468 = \V201(0)  & \V94(16) ;
  assign n469 = \V201(1)  & n468;
  assign n470 = \V201(0)  & \V94(14) ;
  assign n471 = \V201(1)  & n470;
  assign n472 = \V201(0)  & \V94(12) ;
  assign n473 = \V201(1)  & n472;
  assign n474 = \V201(0)  & \V94(10) ;
  assign n475 = \V201(1)  & n474;
  assign n476 = \V201(0)  & \V94(8) ;
  assign n477 = \V201(1)  & n476;
  assign n478 = \V201(0)  & \V94(6) ;
  assign n479 = \V201(1)  & n478;
  assign n480 = \V201(0)  & \V94(4) ;
  assign n481 = \V201(1)  & n480;
  assign n482 = \V94(2)  & \V201(0) ;
  assign n483 = \V201(1)  & n482;
  assign n484 = \V94(3)  & \V201(0) ;
  assign n485 = \V201(1)  & n484;
  assign n486 = \V201(0)  & \V94(5) ;
  assign n487 = \V201(1)  & n486;
  assign n488 = \V201(0)  & \V94(7) ;
  assign n489 = \V201(1)  & n488;
  assign n490 = \V201(0)  & \V94(9) ;
  assign n491 = \V201(1)  & n490;
  assign n492 = \V201(0)  & \V94(11) ;
  assign n493 = \V201(1)  & n492;
  assign n494 = \V201(0)  & \V94(13) ;
  assign n495 = \V201(1)  & n494;
  assign n496 = \V201(0)  & \V94(15) ;
  assign n497 = \V201(1)  & n496;
  assign n498 = \V201(0)  & \V94(17) ;
  assign n499 = \V201(1)  & n498;
  assign n500 = \V201(0)  & \V94(19) ;
  assign n501 = \V201(1)  & n500;
  assign n502 = \V201(0)  & \V94(21) ;
  assign n503 = \V201(1)  & n502;
  assign n504 = \V201(0)  & \V94(23) ;
  assign n505 = \V201(1)  & n504;
  assign n506 = \V201(0)  & \V94(25) ;
  assign n507 = \V201(1)  & n506;
  assign n508 = \V201(0)  & \V94(27) ;
  assign n509 = \V201(1)  & n508;
  assign n510 = \V201(0)  & \V94(29) ;
  assign n511 = \V201(1)  & n510;
  assign n512 = \V94(31)  & \V201(0) ;
  assign n513 = \V201(1)  & n512;
  assign n514 = \V126(1)  & \V201(0) ;
  assign n515 = \V201(1)  & n514;
  assign n516 = \V201(2)  & ~n217;
  assign n517 = \V201(3)  & ~n217;
  assign n518 = \V193(1)  & \V201(6) ;
  assign n519 = \V193(1)  & \V201(7) ;
  assign n520 = \V193(0)  & \V201(6) ;
  assign n521 = \V201(4)  & \V190(0) ;
  assign n522 = \V201(4)  & \V188(30) ;
  assign n523 = \V201(4)  & \V188(31) ;
  assign n524 = \V201(4)  & \V190(1) ;
  assign n525 = \V201(4)  & \V188(28) ;
  assign n526 = \V201(4)  & \V188(26) ;
  assign n527 = \V201(4)  & \V188(27) ;
  assign n528 = \V201(4)  & \V188(29) ;
  assign n529 = \V201(5)  & \V190(0) ;
  assign n530 = \V201(5)  & \V188(30) ;
  assign n531 = \V201(5)  & \V188(31) ;
  assign n532 = \V201(5)  & \V190(1) ;
  assign n533 = \V201(2)  & \V176(16) ;
  assign n534 = \V201(2)  & \V176(14) ;
  assign n535 = \V201(2)  & \V176(12) ;
  assign n536 = \V201(2)  & \V176(10) ;
  assign n537 = \V201(2)  & \V176(8) ;
  assign n538 = \V201(2)  & \V176(6) ;
  assign n539 = \V201(2)  & \V176(4) ;
  assign n540 = \V201(2)  & \V176(2) ;
  assign n541 = \V201(2)  & \V176(3) ;
  assign n542 = \V201(2)  & \V176(5) ;
  assign n543 = \V201(2)  & \V176(7) ;
  assign n544 = \V201(2)  & \V176(9) ;
  assign n545 = \V201(2)  & \V176(11) ;
  assign n546 = \V201(2)  & \V176(13) ;
  assign n547 = \V201(2)  & \V176(15) ;
  assign n548 = \V201(2)  & \V176(17) ;
  assign n549 = \V201(0)  & \V130(0) ;
  assign n550 = ~\V201(0)  & \V129(0) ;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n548 & n551;
  assign n553 = ~n547 & n552;
  assign n554 = ~n546 & n553;
  assign n555 = ~n545 & n554;
  assign n556 = ~n544 & n555;
  assign n557 = ~n543 & n556;
  assign n558 = ~n542 & n557;
  assign n559 = ~n541 & n558;
  assign n560 = ~n540 & n559;
  assign n561 = ~n539 & n560;
  assign n562 = ~n538 & n561;
  assign n563 = ~n537 & n562;
  assign n564 = ~n536 & n563;
  assign n565 = ~n535 & n564;
  assign n566 = ~n534 & n565;
  assign n567 = ~n533 & n566;
  assign n568 = ~n532 & n567;
  assign n569 = ~n531 & n568;
  assign n570 = ~n530 & n569;
  assign n571 = ~n529 & n570;
  assign n572 = ~n528 & n571;
  assign n573 = ~n527 & n572;
  assign n574 = ~n526 & n573;
  assign n575 = ~n525 & n574;
  assign n576 = ~n524 & n575;
  assign n577 = ~n523 & n576;
  assign n578 = ~n522 & n577;
  assign n579 = ~n521 & n578;
  assign n580 = ~n520 & n579;
  assign n581 = ~n519 & n580;
  assign n582 = ~n518 & n581;
  assign n583 = ~n517 & n582;
  assign n584 = ~n516 & n583;
  assign n585 = ~n515 & n584;
  assign n586 = ~n513 & n585;
  assign n587 = ~n511 & n586;
  assign n588 = ~n509 & n587;
  assign n589 = ~n507 & n588;
  assign n590 = ~n505 & n589;
  assign n591 = ~n503 & n590;
  assign n592 = ~n501 & n591;
  assign n593 = ~n499 & n592;
  assign n594 = ~n497 & n593;
  assign n595 = ~n495 & n594;
  assign n596 = ~n493 & n595;
  assign n597 = ~n491 & n596;
  assign n598 = ~n489 & n597;
  assign n599 = ~n487 & n598;
  assign n600 = ~n485 & n599;
  assign n601 = ~n483 & n600;
  assign n602 = ~n481 & n601;
  assign n603 = ~n479 & n602;
  assign n604 = ~n477 & n603;
  assign n605 = ~n475 & n604;
  assign n606 = ~n473 & n605;
  assign n607 = ~n471 & n606;
  assign n608 = ~n469 & n607;
  assign n609 = ~n467 & n608;
  assign n610 = ~n465 & n609;
  assign n611 = ~n463 & n610;
  assign n612 = ~n461 & n611;
  assign n613 = ~n459 & n612;
  assign n614 = ~n457 & n613;
  assign n615 = ~n455 & n614;
  assign n616 = ~n453 & n615;
  assign n617 = ~n451 & n616;
  assign n618 = ~n449 & n617;
  assign n619 = ~n447 & n618;
  assign n620 = ~n445 & n619;
  assign n621 = ~n443 & n620;
  assign n622 = ~n441 & n621;
  assign n623 = ~n439 & n622;
  assign n624 = ~n437 & n623;
  assign n625 = ~n435 & n624;
  assign n626 = ~n433 & n625;
  assign n627 = ~n431 & n626;
  assign n628 = ~n429 & n627;
  assign n629 = ~n427 & n628;
  assign n630 = ~n425 & n629;
  assign n631 = ~n423 & n630;
  assign n632 = ~n421 & n631;
  assign n633 = ~n419 & n632;
  assign n634 = ~n417 & n633;
  assign n635 = ~n415 & n634;
  assign n636 = ~n413 & n635;
  assign n637 = ~n411 & n636;
  assign n638 = ~n409 & n637;
  assign n639 = ~n407 & n638;
  assign n640 = ~n405 & n639;
  assign n641 = ~n403 & n640;
  assign n642 = ~n401 & n641;
  assign n643 = ~n399 & n642;
  assign n644 = ~n397 & n643;
  assign n645 = ~n395 & n644;
  assign n646 = ~n393 & n645;
  assign n647 = ~n391 & n646;
  assign n648 = ~n389 & n647;
  assign n649 = ~n387 & n648;
  assign n650 = ~n385 & n649;
  assign n651 = ~n383 & n650;
  assign n652 = ~n381 & n651;
  assign n653 = ~n379 & n652;
  assign n654 = ~n377 & n653;
  assign n655 = ~n375 & n654;
  assign n656 = ~n373 & n655;
  assign n657 = ~n371 & n656;
  assign n658 = ~n369 & n657;
  assign n659 = ~n367 & n658;
  assign n660 = ~n365 & n659;
  assign n661 = ~n363 & n660;
  assign n662 = ~n361 & n661;
  assign n663 = ~n359 & n662;
  assign n664 = ~n357 & n663;
  assign n665 = ~n355 & n664;
  assign n666 = ~n353 & n665;
  assign n667 = ~n351 & n666;
  assign n668 = ~n349 & n667;
  assign n669 = ~n347 & n668;
  assign n670 = ~n345 & n669;
  assign n671 = ~n343 & n670;
  assign n672 = ~n341 & n671;
  assign n673 = ~n339 & n672;
  assign n674 = ~n337 & n673;
  assign n675 = ~n335 & n674;
  assign n676 = ~n333 & n675;
  assign n677 = ~n331 & n676;
  assign n678 = ~n329 & n677;
  assign n679 = ~n327 & n678;
  assign n680 = ~n325 & n679;
  assign n681 = ~n323 & n680;
  assign n682 = ~n321 & n681;
  assign n683 = ~n319 & n682;
  assign n684 = ~n317 & n683;
  assign n685 = ~n315 & n684;
  assign n686 = ~n313 & n685;
  assign n687 = ~n311 & n686;
  assign n688 = ~n309 & n687;
  assign n689 = ~n307 & n688;
  assign n690 = ~n305 & n689;
  assign n691 = ~n303 & n690;
  assign n692 = ~n301 & n691;
  assign n693 = ~n299 & n692;
  assign n694 = ~n297 & n693;
  assign n695 = ~n295 & n694;
  assign n696 = ~n293 & n695;
  assign n697 = ~n291 & n696;
  assign n698 = ~n289 & n697;
  assign n699 = ~n287 & n698;
  assign n700 = ~n285 & n699;
  assign n701 = ~n283 & n700;
  assign n702 = ~n281 & n701;
  assign n703 = ~n279 & n702;
  assign n704 = ~n277 & n703;
  assign n705 = ~n275 & n704;
  assign n706 = ~n273 & n705;
  assign n707 = ~n271 & n706;
  assign n708 = ~n269 & n707;
  assign n709 = ~n267 & n708;
  assign n710 = ~n265 & n709;
  assign n711 = ~n263 & n710;
  assign n712 = ~n261 & n711;
  assign n713 = ~n259 & n712;
  assign n714 = ~n257 & n713;
  assign n715 = ~n255 & n714;
  assign n716 = ~n253 & n715;
  assign n717 = ~n251 & n716;
  assign n718 = ~n249 & n717;
  assign n719 = ~n247 & n718;
  assign n720 = ~n245 & n719;
  assign n721 = ~n243 & n720;
  assign n722 = ~n241 & n721;
  assign n723 = ~n239 & n722;
  assign n724 = ~n237 & n723;
  assign n725 = ~n235 & n724;
  assign n726 = ~n233 & n725;
  assign n727 = ~n231 & n726;
  assign n728 = ~n229 & n727;
  assign n729 = ~n227 & n728;
  assign n730 = ~n225 & n729;
  assign n731 = ~n223 & n730;
  assign n732 = ~n221 & n731;
  assign \V202(0)  = n219 | ~n732;
endmodule


