// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:02 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_;
  wire n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
    n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1436, n1437, n1438, n1439, n1440, n1441,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1467, n1468, n1469, n1470, n1471, n1472, n1474,
    n1475, n1476, n1478, n1479, n1480;
  assign n30 = ~i_3_ & i_4_;
  assign n31 = ~i_5_ & n30;
  assign n32 = i_0_ & ~i_1_;
  assign n33 = ~i_2_ & n32;
  assign n34 = i_6_ & ~i_7_;
  assign n35 = ~i_8_ & n34;
  assign n36 = n33 & n35;
  assign n37 = n31 & n36;
  assign n38 = ~i_4_ & i_5_;
  assign n39 = ~i_3_ & n38;
  assign n40 = i_7_ & ~i_8_;
  assign n41 = i_0_ & i_1_;
  assign n42 = ~i_2_ & n41;
  assign n43 = ~i_6_ & n42;
  assign n44 = n40 & n43;
  assign n45 = n39 & n44;
  assign n46 = ~n37 & ~n45;
  assign n47 = ~i_6_ & i_7_;
  assign n48 = i_8_ & n47;
  assign n49 = n33 & n48;
  assign n50 = n31 & n49;
  assign n51 = i_5_ & n30;
  assign n52 = i_6_ & i_8_;
  assign n53 = ~i_7_ & n52;
  assign n54 = n33 & n53;
  assign n55 = n51 & n54;
  assign n56 = ~n50 & ~n55;
  assign n57 = i_4_ & i_5_;
  assign n58 = i_7_ & n57;
  assign n59 = i_0_ & ~i_2_;
  assign n60 = ~i_6_ & i_8_;
  assign n61 = i_3_ & n60;
  assign n62 = n59 & n61;
  assign n63 = n58 & n62;
  assign n64 = n56 & ~n63;
  assign n65 = n46 & n64;
  assign n66 = ~i_3_ & i_5_;
  assign n67 = i_2_ & n41;
  assign n68 = n66 & n67;
  assign n69 = ~i_4_ & n68;
  assign n70 = n35 & n69;
  assign n71 = ~i_6_ & ~i_7_;
  assign n72 = n30 & n41;
  assign n73 = i_2_ & i_5_;
  assign n74 = n72 & n73;
  assign n75 = n71 & n74;
  assign n76 = i_3_ & ~i_5_;
  assign n77 = ~i_4_ & n76;
  assign n78 = ~i_6_ & ~i_8_;
  assign n79 = ~i_7_ & n78;
  assign n80 = n33 & n79;
  assign n81 = n77 & n80;
  assign n82 = ~n75 & ~n81;
  assign n83 = ~n70 & n82;
  assign n84 = n65 & n83;
  assign n85 = i_3_ & ~i_4_;
  assign n86 = i_5_ & n85;
  assign n87 = n33 & n40;
  assign n88 = i_6_ & n87;
  assign n89 = n86 & n88;
  assign n90 = ~i_6_ & n40;
  assign n91 = n33 & n90;
  assign n92 = i_3_ & i_4_;
  assign n93 = n91 & n92;
  assign n94 = ~i_7_ & i_8_;
  assign n95 = ~i_6_ & n94;
  assign n96 = n33 & n95;
  assign n97 = n85 & n96;
  assign n98 = ~n93 & ~n97;
  assign n99 = ~n89 & n98;
  assign n100 = i_6_ & i_7_;
  assign n101 = i_8_ & n100;
  assign n102 = n33 & n101;
  assign n103 = n86 & n102;
  assign n104 = n53 & n69;
  assign n105 = ~n103 & ~n104;
  assign n106 = n39 & n59;
  assign n107 = n95 & n106;
  assign n108 = n105 & ~n107;
  assign n109 = n99 & n108;
  assign n110 = n84 & n109;
  assign n111 = ~i_3_ & ~i_5_;
  assign n112 = ~i_4_ & n111;
  assign n113 = n67 & n112;
  assign n114 = n53 & n113;
  assign n115 = ~i_8_ & n100;
  assign n116 = ~i_0_ & i_1_;
  assign n117 = i_2_ & n116;
  assign n118 = n31 & n117;
  assign n119 = n115 & n118;
  assign n120 = ~i_2_ & n116;
  assign n121 = n39 & n120;
  assign n122 = n115 & n121;
  assign n123 = ~n119 & ~n122;
  assign n124 = ~n114 & n123;
  assign n125 = n69 & n115;
  assign n126 = n77 & n102;
  assign n127 = ~i_5_ & n92;
  assign n128 = i_2_ & n32;
  assign n129 = n115 & n128;
  assign n130 = n127 & n129;
  assign n131 = ~n126 & ~n130;
  assign n132 = ~n125 & n131;
  assign n133 = n124 & n132;
  assign n134 = ~i_6_ & n38;
  assign n135 = n87 & n134;
  assign n136 = n86 & n117;
  assign n137 = n35 & n136;
  assign n138 = ~n135 & ~n137;
  assign n139 = n31 & n67;
  assign n140 = n79 & n139;
  assign n141 = n120 & n127;
  assign n142 = n48 & n141;
  assign n143 = n42 & n112;
  assign n144 = n95 & n143;
  assign n145 = ~n142 & ~n144;
  assign n146 = ~n140 & n145;
  assign n147 = n138 & n146;
  assign n148 = i_5_ & n92;
  assign n149 = n128 & n148;
  assign n150 = n41 & n148;
  assign n151 = ~i_2_ & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = n100 & ~n152;
  assign n154 = n79 & n127;
  assign n155 = n32 & n154;
  assign n156 = ~n153 & ~n155;
  assign n157 = n147 & n156;
  assign n158 = n133 & n157;
  assign n159 = n110 & n158;
  assign n160 = n77 & n88;
  assign n161 = n53 & n128;
  assign n162 = n127 & n161;
  assign n163 = n48 & n136;
  assign n164 = n35 & n113;
  assign n165 = ~n163 & ~n164;
  assign n166 = ~n162 & n165;
  assign n167 = ~n160 & n166;
  assign n168 = n101 & n113;
  assign n169 = n71 & n149;
  assign n170 = ~n168 & ~n169;
  assign n171 = n112 & n120;
  assign n172 = n53 & n171;
  assign n173 = n112 & n117;
  assign n174 = n53 & n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = n170 & n175;
  assign n177 = n167 & n176;
  assign n178 = n111 & n117;
  assign n179 = i_4_ & n101;
  assign n180 = n178 & n179;
  assign n181 = n92 & n120;
  assign n182 = i_5_ & n181;
  assign n183 = n35 & n182;
  assign n184 = n117 & n148;
  assign n185 = n115 & n184;
  assign n186 = ~i_3_ & ~i_4_;
  assign n187 = n117 & n186;
  assign n188 = i_5_ & n187;
  assign n189 = n115 & n188;
  assign n190 = ~n185 & ~n189;
  assign n191 = ~n183 & n190;
  assign n192 = ~n180 & n191;
  assign n193 = n177 & n192;
  assign n194 = n69 & n79;
  assign n195 = n101 & n128;
  assign n196 = n86 & n195;
  assign n197 = n35 & n128;
  assign n198 = n86 & n197;
  assign n199 = n53 & n57;
  assign n200 = i_2_ & i_3_;
  assign n201 = ~i_1_ & n200;
  assign n202 = n199 & n201;
  assign n203 = ~n198 & ~n202;
  assign n204 = ~n196 & n203;
  assign n205 = ~n194 & n204;
  assign n206 = n193 & n205;
  assign o_1_ = ~n159 | ~n206;
  assign n208 = ~i_0_ & ~i_1_;
  assign n209 = i_2_ & n208;
  assign n210 = n127 & n209;
  assign n211 = n115 & n210;
  assign n212 = n31 & n54;
  assign n213 = ~n211 & ~n212;
  assign n214 = n53 & n86;
  assign n215 = n42 & n214;
  assign n216 = n213 & ~n215;
  assign n217 = n117 & n127;
  assign n218 = n95 & n217;
  assign n219 = n148 & n209;
  assign n220 = n35 & n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = n48 & n210;
  assign n223 = n221 & ~n222;
  assign n224 = n216 & n223;
  assign n225 = n209 & n214;
  assign n226 = n90 & n184;
  assign n227 = ~n225 & ~n226;
  assign n228 = n69 & n101;
  assign n229 = n94 & n184;
  assign n230 = n54 & n77;
  assign n231 = n112 & n129;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n229 & n232;
  assign n234 = ~n228 & n233;
  assign n235 = n227 & n234;
  assign n236 = n224 & n235;
  assign n237 = ~i_7_ & ~i_8_;
  assign n238 = ~n106 & ~n150;
  assign n239 = n237 & ~n238;
  assign n240 = n31 & n209;
  assign n241 = n79 & n240;
  assign n242 = n35 & n171;
  assign n243 = ~n241 & ~n242;
  assign n244 = ~n239 & n243;
  assign n245 = n95 & n128;
  assign n246 = n86 & n245;
  assign n247 = n51 & n91;
  assign n248 = ~n246 & ~n247;
  assign n249 = i_4_ & ~i_5_;
  assign n250 = n42 & n249;
  assign n251 = i_3_ & n250;
  assign n252 = n40 & n251;
  assign n253 = n248 & ~n252;
  assign n254 = n35 & n173;
  assign n255 = i_7_ & i_8_;
  assign n256 = n77 & n128;
  assign n257 = n255 & n256;
  assign n258 = ~n254 & ~n257;
  assign n259 = n39 & n209;
  assign n260 = n101 & n259;
  assign n261 = n36 & n148;
  assign n262 = ~n260 & ~n261;
  assign n263 = n258 & n262;
  assign n264 = n253 & n263;
  assign n265 = n39 & n94;
  assign n266 = n117 & n265;
  assign n267 = i_0_ & i_2_;
  assign n268 = n58 & n267;
  assign n269 = ~i_3_ & n268;
  assign n270 = ~n266 & ~n269;
  assign n271 = n264 & n270;
  assign n272 = n244 & n271;
  assign n273 = n236 & n272;
  assign n274 = n61 & n249;
  assign n275 = i_5_ & n79;
  assign n276 = ~i_4_ & ~i_5_;
  assign n277 = n95 & n276;
  assign n278 = i_3_ & n277;
  assign n279 = ~n275 & ~n278;
  assign n280 = ~n274 & n279;
  assign n281 = n33 & ~n280;
  assign n282 = n79 & n121;
  assign n283 = n90 & n136;
  assign n284 = ~n282 & ~n283;
  assign n285 = n115 & n219;
  assign n286 = n284 & ~n285;
  assign n287 = i_3_ & i_5_;
  assign n288 = n101 & n287;
  assign n289 = n41 & n288;
  assign n290 = n51 & n117;
  assign n291 = n35 & n290;
  assign n292 = n39 & n48;
  assign n293 = n41 & n292;
  assign n294 = ~n291 & ~n293;
  assign n295 = ~n289 & n294;
  assign n296 = n286 & n295;
  assign n297 = ~n281 & n296;
  assign n298 = n48 & n276;
  assign n299 = n267 & n298;
  assign n300 = n79 & n287;
  assign n301 = n117 & n300;
  assign n302 = i_4_ & n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = n115 & n139;
  assign n305 = n67 & n148;
  assign n306 = n100 & n305;
  assign n307 = ~i_5_ & n197;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~n304 & n308;
  assign n310 = n303 & n309;
  assign n311 = n297 & n310;
  assign n312 = n273 & n311;
  assign n313 = n53 & n182;
  assign n314 = n245 & n249;
  assign n315 = ~n313 & ~n314;
  assign n316 = n31 & n120;
  assign n317 = n90 & n316;
  assign n318 = n33 & n214;
  assign n319 = n42 & n115;
  assign n320 = n31 & n319;
  assign n321 = ~n318 & ~n320;
  assign n322 = ~n317 & n321;
  assign n323 = n90 & n151;
  assign n324 = i_2_ & ~i_3_;
  assign n325 = n32 & n38;
  assign n326 = n324 & n325;
  assign n327 = n47 & n326;
  assign n328 = ~n323 & ~n327;
  assign n329 = n322 & n328;
  assign n330 = n315 & n329;
  assign n331 = n101 & n184;
  assign n332 = n53 & n305;
  assign n333 = n42 & n101;
  assign n334 = n39 & n333;
  assign n335 = n67 & n127;
  assign n336 = n95 & n335;
  assign n337 = ~n334 & ~n336;
  assign n338 = ~n332 & n337;
  assign n339 = n101 & n120;
  assign n340 = n31 & n339;
  assign n341 = n338 & ~n340;
  assign n342 = ~n331 & n341;
  assign n343 = n330 & n342;
  assign n344 = n35 & n149;
  assign n345 = n90 & n128;
  assign n346 = n86 & n345;
  assign n347 = n39 & n339;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n344 & n348;
  assign n350 = n57 & n95;
  assign n351 = n77 & n237;
  assign n352 = n40 & n86;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n350 & n353;
  assign n355 = n42 & ~n354;
  assign n356 = n349 & ~n355;
  assign n357 = n85 & n90;
  assign n358 = n41 & n357;
  assign n359 = i_1_ & ~i_2_;
  assign n360 = n79 & n359;
  assign n361 = n111 & n360;
  assign n362 = ~n358 & ~n361;
  assign n363 = n112 & n195;
  assign n364 = n117 & n154;
  assign n365 = ~n363 & ~n364;
  assign n366 = n30 & n42;
  assign n367 = n77 & n209;
  assign n368 = ~n366 & ~n367;
  assign n369 = n47 & ~n368;
  assign n370 = n365 & ~n369;
  assign n371 = n362 & n370;
  assign n372 = n356 & n371;
  assign n373 = n36 & n51;
  assign n374 = n86 & n209;
  assign n375 = n35 & n374;
  assign n376 = n90 & n290;
  assign n377 = i_0_ & n200;
  assign n378 = n38 & n377;
  assign n379 = n48 & n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~n375 & n380;
  assign n382 = ~n373 & n381;
  assign n383 = n71 & n287;
  assign n384 = ~i_3_ & n179;
  assign n385 = ~n383 & ~n384;
  assign n386 = n67 & ~n385;
  assign n387 = n116 & n127;
  assign n388 = ~i_3_ & n32;
  assign n389 = ~i_4_ & n388;
  assign n390 = ~n387 & ~n389;
  assign n391 = n35 & ~n390;
  assign n392 = n92 & n96;
  assign n393 = ~n391 & ~n392;
  assign n394 = ~n386 & n393;
  assign n395 = n382 & n394;
  assign n396 = n372 & n395;
  assign n397 = n90 & n118;
  assign n398 = n112 & n115;
  assign n399 = n59 & n398;
  assign n400 = ~n397 & ~n399;
  assign n401 = n94 & n139;
  assign n402 = n51 & n209;
  assign n403 = n71 & n402;
  assign n404 = ~n401 & ~n403;
  assign n405 = n400 & n404;
  assign n406 = n77 & n91;
  assign n407 = n102 & n127;
  assign n408 = ~n406 & ~n407;
  assign n409 = n53 & n118;
  assign n410 = n79 & n113;
  assign n411 = ~n409 & ~n410;
  assign n412 = n408 & n411;
  assign n413 = n405 & n412;
  assign n414 = n112 & n128;
  assign n415 = n71 & n414;
  assign n416 = n120 & n265;
  assign n417 = ~n415 & ~n416;
  assign n418 = n31 & n161;
  assign n419 = n47 & n217;
  assign n420 = ~n418 & ~n419;
  assign n421 = n48 & n128;
  assign n422 = ~i_3_ & n421;
  assign n423 = n59 & n78;
  assign n424 = n31 & n423;
  assign n425 = ~n422 & ~n424;
  assign n426 = n420 & n425;
  assign n427 = n417 & n426;
  assign n428 = n101 & n117;
  assign n429 = n66 & n428;
  assign n430 = n67 & n77;
  assign n431 = n53 & n430;
  assign n432 = n116 & n398;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n429 & n433;
  assign n435 = n48 & n249;
  assign n436 = ~n277 & ~n435;
  assign n437 = i_1_ & n200;
  assign n438 = ~n436 & n437;
  assign n439 = n43 & n287;
  assign n440 = n94 & n439;
  assign n441 = ~n438 & ~n440;
  assign n442 = n434 & n441;
  assign n443 = n427 & n442;
  assign n444 = n413 & n443;
  assign n445 = n396 & n444;
  assign n446 = n343 & n445;
  assign n447 = n48 & n184;
  assign n448 = n44 & n112;
  assign n449 = ~n447 & ~n448;
  assign n450 = n47 & n120;
  assign n451 = n86 & n450;
  assign n452 = ~i_8_ & n451;
  assign n453 = n449 & ~n452;
  assign n454 = n67 & n154;
  assign n455 = n42 & n77;
  assign n456 = n95 & n455;
  assign n457 = ~n454 & ~n456;
  assign n458 = n53 & n388;
  assign n459 = n276 & n458;
  assign n460 = n95 & n290;
  assign n461 = n77 & n117;
  assign n462 = n79 & n461;
  assign n463 = ~n460 & ~n462;
  assign n464 = ~n459 & n463;
  assign n465 = n457 & n464;
  assign n466 = n48 & n182;
  assign n467 = n71 & n136;
  assign n468 = ~n466 & ~n467;
  assign n469 = n47 & n461;
  assign n470 = n95 & n316;
  assign n471 = ~n469 & ~n470;
  assign n472 = n31 & n42;
  assign n473 = n34 & n472;
  assign n474 = n31 & n345;
  assign n475 = ~n473 & ~n474;
  assign n476 = n471 & n475;
  assign n477 = n468 & n476;
  assign n478 = n465 & n477;
  assign n479 = n53 & n251;
  assign n480 = n77 & n129;
  assign n481 = n31 & n102;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n479 & n482;
  assign n484 = n101 & n217;
  assign n485 = n86 & n120;
  assign n486 = n95 & n485;
  assign n487 = ~n484 & ~n486;
  assign n488 = n483 & n487;
  assign n489 = n49 & n57;
  assign n490 = ~i_3_ & n489;
  assign n491 = n276 & n377;
  assign n492 = n35 & n491;
  assign n493 = ~n490 & ~n492;
  assign n494 = n113 & n115;
  assign n495 = n127 & n195;
  assign n496 = ~n494 & ~n495;
  assign n497 = n493 & n496;
  assign n498 = n488 & n497;
  assign n499 = n478 & n498;
  assign n500 = n453 & n499;
  assign n501 = n53 & n141;
  assign n502 = n34 & n485;
  assign n503 = ~i_8_ & n502;
  assign n504 = ~n501 & ~n503;
  assign n505 = n54 & n148;
  assign n506 = n112 & n333;
  assign n507 = n35 & n42;
  assign n508 = n66 & n507;
  assign n509 = ~n506 & ~n508;
  assign n510 = ~n505 & n509;
  assign n511 = n76 & n450;
  assign n512 = ~i_8_ & n511;
  assign n513 = n510 & ~n512;
  assign n514 = n504 & n513;
  assign n515 = n90 & n335;
  assign n516 = n38 & n161;
  assign n517 = n39 & n49;
  assign n518 = ~n516 & ~n517;
  assign n519 = n48 & n251;
  assign n520 = n518 & ~n519;
  assign n521 = n48 & n455;
  assign n522 = n39 & n102;
  assign n523 = ~n521 & ~n522;
  assign n524 = n101 & n219;
  assign n525 = n148 & n339;
  assign n526 = ~n524 & ~n525;
  assign n527 = n523 & n526;
  assign n528 = n520 & n527;
  assign n529 = ~n515 & n528;
  assign n530 = n514 & n529;
  assign n531 = n79 & n128;
  assign n532 = n76 & n531;
  assign n533 = n51 & n88;
  assign n534 = n101 & n210;
  assign n535 = n35 & n210;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n533 & n536;
  assign n538 = ~n532 & n537;
  assign n539 = n530 & n538;
  assign n540 = n500 & n539;
  assign n541 = n446 & n540;
  assign o_2_ = ~n312 | ~n541;
  assign n543 = n30 & n275;
  assign n544 = n116 & n543;
  assign n545 = i_6_ & ~i_8_;
  assign n546 = n67 & n85;
  assign n547 = n545 & n546;
  assign n548 = ~n544 & ~n547;
  assign n549 = n58 & n60;
  assign n550 = n201 & n549;
  assign n551 = n101 & n335;
  assign n552 = ~n550 & ~n551;
  assign n553 = n95 & n118;
  assign n554 = n53 & n72;
  assign n555 = ~n553 & ~n554;
  assign n556 = n552 & n555;
  assign n557 = n548 & n556;
  assign n558 = ~n364 & n557;
  assign n559 = n36 & n86;
  assign n560 = n48 & n290;
  assign n561 = n115 & n181;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n559 & n562;
  assign n564 = n112 & n339;
  assign n565 = i_1_ & n324;
  assign n566 = n298 & n565;
  assign n567 = ~n564 & ~n566;
  assign n568 = n100 & n461;
  assign n569 = n567 & ~n568;
  assign n570 = n563 & n569;
  assign n571 = n31 & n91;
  assign n572 = ~i_2_ & n389;
  assign n573 = n48 & n572;
  assign n574 = ~n571 & ~n573;
  assign n575 = n570 & n574;
  assign n576 = n234 & n575;
  assign n577 = n558 & n576;
  assign n578 = n53 & n209;
  assign n579 = n127 & n578;
  assign n580 = n79 & n485;
  assign n581 = i_6_ & n266;
  assign n582 = n48 & n171;
  assign n583 = n100 & n143;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n581 & n584;
  assign n586 = ~n580 & n585;
  assign n587 = n101 & n240;
  assign n588 = n35 & n118;
  assign n589 = ~n587 & ~n588;
  assign n590 = n586 & n589;
  assign n591 = n167 & n590;
  assign n592 = ~n579 & n591;
  assign n593 = n577 & n592;
  assign n594 = n38 & n47;
  assign n595 = n565 & n594;
  assign n596 = ~i_8_ & n595;
  assign n597 = n38 & n48;
  assign n598 = n201 & n597;
  assign n599 = ~n226 & ~n598;
  assign n600 = n221 & n599;
  assign n601 = ~n596 & n600;
  assign n602 = n129 & n148;
  assign n603 = n115 & n259;
  assign n604 = ~n602 & ~n603;
  assign n605 = n105 & n604;
  assign n606 = ~n331 & n605;
  assign n607 = n601 & n606;
  assign n608 = n51 & n360;
  assign n609 = ~n304 & ~n608;
  assign n610 = ~n81 & n609;
  assign n611 = ~n151 & ~n290;
  assign n612 = n115 & ~n611;
  assign n613 = n101 & n430;
  assign n614 = n73 & n388;
  assign n615 = n71 & n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n196 & n616;
  assign n618 = ~n612 & n617;
  assign n619 = n610 & n618;
  assign n620 = n249 & n333;
  assign n621 = n350 & n388;
  assign n622 = n128 & n237;
  assign n623 = n134 & n622;
  assign n624 = ~n621 & ~n623;
  assign n625 = ~n620 & n624;
  assign n626 = n619 & n625;
  assign n627 = n607 & n626;
  assign n628 = n201 & n277;
  assign n629 = n35 & n188;
  assign n630 = n38 & n129;
  assign n631 = n42 & n199;
  assign n632 = ~n630 & ~n631;
  assign n633 = n51 & n102;
  assign n634 = n632 & ~n633;
  assign n635 = ~n629 & n634;
  assign n636 = n100 & n217;
  assign n637 = ~i_8_ & n636;
  assign n638 = n635 & ~n637;
  assign n639 = ~n628 & n638;
  assign n640 = n95 & n472;
  assign n641 = ~n430 & ~n572;
  assign n642 = n79 & ~n641;
  assign n643 = n112 & n345;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~n640 & n644;
  assign n646 = n80 & n148;
  assign n647 = n53 & n485;
  assign n648 = n35 & n184;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n646 & n649;
  assign n651 = n645 & n650;
  assign n652 = n639 & n651;
  assign n653 = n627 & n652;
  assign n654 = n39 & n319;
  assign n655 = n127 & n507;
  assign n656 = ~n654 & ~n655;
  assign n657 = n102 & n148;
  assign n658 = n53 & n256;
  assign n659 = n187 & n275;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n657 & n660;
  assign n662 = ~n181 & ~n210;
  assign n663 = n90 & ~n662;
  assign n664 = n31 & n88;
  assign n665 = ~n663 & ~n664;
  assign n666 = n661 & n665;
  assign n667 = n656 & n666;
  assign n668 = n92 & n307;
  assign n669 = n86 & n507;
  assign n670 = n53 & n217;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n668 & n671;
  assign n673 = ~n462 & n672;
  assign n674 = n95 & n141;
  assign n675 = n51 & n161;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n178 & ~n305;
  assign n678 = n48 & ~n677;
  assign n679 = n96 & n249;
  assign n680 = ~n347 & ~n679;
  assign n681 = ~n678 & n680;
  assign n682 = n676 & n681;
  assign n683 = n673 & n682;
  assign n684 = n51 & n333;
  assign n685 = n31 & n531;
  assign n686 = ~n684 & ~n685;
  assign n687 = n48 & n485;
  assign n688 = ~n407 & ~n687;
  assign n689 = n686 & n688;
  assign n690 = n112 & n423;
  assign n691 = ~i_7_ & n690;
  assign n692 = n77 & n120;
  assign n693 = n60 & n692;
  assign n694 = ~n691 & ~n693;
  assign n695 = n115 & n316;
  assign n696 = ~n254 & ~n695;
  assign n697 = n694 & n696;
  assign n698 = n689 & n697;
  assign n699 = n683 & n698;
  assign n700 = n667 & n699;
  assign n701 = n71 & n251;
  assign n702 = n32 & n39;
  assign n703 = n115 & n702;
  assign n704 = n77 & n345;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~n701 & n705;
  assign n707 = n42 & n300;
  assign n708 = ~i_4_ & n707;
  assign n709 = ~n323 & ~n373;
  assign n710 = ~n708 & n709;
  assign n711 = n77 & n333;
  assign n712 = n67 & n100;
  assign n713 = ~i_8_ & n712;
  assign n714 = n127 & n713;
  assign n715 = ~n711 & ~n714;
  assign n716 = n120 & n398;
  assign n717 = n52 & n290;
  assign n718 = n79 & n173;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n716 & n719;
  assign n721 = n715 & n720;
  assign n722 = n710 & n721;
  assign n723 = n706 & n722;
  assign n724 = n468 & n723;
  assign n725 = n700 & n724;
  assign n726 = n653 & n725;
  assign o_3_ = ~n593 | ~n726;
  assign n728 = n35 & n151;
  assign n729 = n85 & n428;
  assign n730 = ~n533 & ~n729;
  assign n731 = ~n728 & n730;
  assign n732 = n90 & n171;
  assign n733 = n49 & n287;
  assign n734 = ~n732 & ~n733;
  assign n735 = n731 & n734;
  assign n736 = n34 & n414;
  assign n737 = n86 & n161;
  assign n738 = n115 & n461;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = i_2_ & n543;
  assign n742 = ~i_0_ & i_2_;
  assign n743 = n357 & n742;
  assign n744 = ~n741 & ~n743;
  assign n745 = n740 & n744;
  assign n746 = n735 & n745;
  assign n747 = n95 & n173;
  assign n748 = ~n517 & ~n747;
  assign n749 = n33 & n71;
  assign n750 = n112 & n749;
  assign n751 = ~n107 & ~n750;
  assign n752 = n748 & n751;
  assign n753 = n746 & n752;
  assign n754 = n35 & n472;
  assign n755 = n115 & n209;
  assign n756 = ~n161 & ~n755;
  assign n757 = ~n87 & n756;
  assign n758 = n148 & ~n757;
  assign n759 = ~n754 & ~n758;
  assign n760 = n79 & n692;
  assign n761 = n74 & n237;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n70 & ~n89;
  assign n764 = ~i_8_ & n701;
  assign n765 = n763 & ~n764;
  assign n766 = n762 & n765;
  assign n767 = n42 & n265;
  assign n768 = ~n581 & ~n648;
  assign n769 = ~n767 & n768;
  assign n770 = n53 & n316;
  assign n771 = ~n459 & ~n770;
  assign n772 = n53 & n461;
  assign n773 = n771 & ~n772;
  assign n774 = n769 & n773;
  assign n775 = n766 & n774;
  assign n776 = n759 & n775;
  assign n777 = n141 & n545;
  assign n778 = n483 & ~n777;
  assign n779 = n95 & n182;
  assign n780 = n39 & n54;
  assign n781 = ~n779 & ~n780;
  assign n782 = n778 & n781;
  assign n783 = n619 & n782;
  assign n784 = ~n182 & ~n250;
  assign n785 = n90 & ~n784;
  assign n786 = n303 & ~n785;
  assign n787 = n683 & n786;
  assign n788 = n783 & n787;
  assign n789 = n776 & n788;
  assign n790 = n753 & n789;
  assign n791 = n298 & n388;
  assign n792 = i_8_ & n75;
  assign n793 = ~n791 & ~n792;
  assign n794 = n48 & n219;
  assign n795 = n39 & n578;
  assign n796 = ~n551 & ~n795;
  assign n797 = ~n794 & n796;
  assign n798 = n793 & n797;
  assign n799 = n31 & n195;
  assign n800 = n77 & n319;
  assign n801 = ~n799 & ~n800;
  assign n802 = n255 & n472;
  assign n803 = n40 & n430;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n45 & n804;
  assign n806 = n801 & n805;
  assign n807 = n79 & n141;
  assign n808 = n277 & n377;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n506 & ~n646;
  assign n811 = n809 & n810;
  assign n812 = ~n172 & ~n707;
  assign n813 = n811 & n812;
  assign n814 = n806 & n813;
  assign n815 = n798 & n814;
  assign n816 = n95 & n210;
  assign n817 = n51 & n197;
  assign n818 = ~n691 & ~n817;
  assign n819 = ~n816 & n818;
  assign n820 = n276 & n428;
  assign n821 = n48 & n692;
  assign n822 = ~n716 & ~n821;
  assign n823 = ~n820 & n822;
  assign n824 = n819 & n823;
  assign n825 = n33 & n543;
  assign n826 = n53 & n335;
  assign n827 = ~n825 & ~n826;
  assign n828 = i_5_ & n547;
  assign n829 = n79 & n178;
  assign n830 = ~n484 & ~n829;
  assign n831 = ~n828 & n830;
  assign n832 = n827 & n831;
  assign n833 = n824 & n832;
  assign n834 = n686 & n833;
  assign n835 = ~n637 & ~n647;
  assign n836 = n35 & n121;
  assign n837 = ~i_1_ & n690;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n228 & n838;
  assign n840 = n835 & n839;
  assign n841 = n90 & n219;
  assign n842 = n42 & n597;
  assign n843 = n77 & n339;
  assign n844 = n58 & n78;
  assign n845 = n67 & n844;
  assign n846 = ~n843 & ~n845;
  assign n847 = ~n842 & n846;
  assign n848 = ~n841 & n847;
  assign n849 = n840 & n848;
  assign n850 = n264 & n849;
  assign n851 = n834 & n850;
  assign n852 = n815 & n851;
  assign n853 = n69 & n95;
  assign n854 = n90 & n149;
  assign n855 = ~n853 & ~n854;
  assign n856 = n100 & n326;
  assign n857 = n51 & n319;
  assign n858 = ~n856 & ~n857;
  assign n859 = n53 & n143;
  assign n860 = ~n230 & ~n859;
  assign n861 = n858 & n860;
  assign n862 = n855 & n861;
  assign n863 = n88 & n127;
  assign n864 = n47 & n187;
  assign n865 = ~n331 & ~n864;
  assign n866 = ~n863 & n865;
  assign n867 = ~n466 & n866;
  assign n868 = n862 & n867;
  assign n869 = i_5_ & n546;
  assign n870 = n53 & n869;
  assign n871 = n35 & n139;
  assign n872 = ~n870 & ~n871;
  assign n873 = n31 & n755;
  assign n874 = ~n460 & ~n873;
  assign n875 = n79 & n367;
  assign n876 = n874 & ~n875;
  assign n877 = n872 & n876;
  assign n878 = n635 & n877;
  assign n879 = n868 & n878;
  assign n880 = n715 & n879;
  assign n881 = ~i_7_ & n717;
  assign n882 = n880 & ~n881;
  assign n883 = n852 & n882;
  assign o_4_ = ~n790 | ~n883;
  assign n885 = n79 & n182;
  assign n886 = n801 & ~n885;
  assign n887 = ~n587 & n886;
  assign n888 = n79 & n210;
  assign n889 = n95 & n219;
  assign n890 = n90 & n276;
  assign n891 = n565 & n890;
  assign n892 = n35 & n316;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n889 & n893;
  assign n895 = ~n888 & n894;
  assign n896 = n887 & n895;
  assign n897 = ~n841 & n896;
  assign n898 = n213 & n349;
  assign n899 = i_3_ & n421;
  assign n900 = n35 & n461;
  assign n901 = ~n899 & ~n900;
  assign n902 = n51 & n339;
  assign n903 = n100 & n141;
  assign n904 = ~n902 & ~n903;
  assign n905 = n901 & n904;
  assign n906 = n54 & n127;
  assign n907 = n35 & n143;
  assign n908 = n435 & n565;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n906 & n909;
  assign n911 = n905 & n910;
  assign n912 = n898 & n911;
  assign n913 = ~n551 & n731;
  assign n914 = ~n282 & n913;
  assign n915 = n912 & n914;
  assign n916 = n897 & n915;
  assign n917 = n48 & n121;
  assign n918 = ~n340 & ~n917;
  assign n919 = n35 & n335;
  assign n920 = n102 & n112;
  assign n921 = ~n919 & ~n920;
  assign n922 = n53 & n455;
  assign n923 = ~n670 & ~n922;
  assign n924 = n921 & n923;
  assign n925 = n918 & n924;
  assign n926 = ~n285 & ~n674;
  assign n927 = n925 & n926;
  assign n928 = n79 & n305;
  assign n929 = n48 & n430;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n242 & n930;
  assign n932 = ~n440 & n931;
  assign n933 = ~n318 & n932;
  assign n934 = n723 & n933;
  assign n935 = n927 & n934;
  assign n936 = n916 & n935;
  assign n937 = i_8_ & n864;
  assign n938 = ~n779 & ~n937;
  assign n939 = n100 & n485;
  assign n940 = n40 & n692;
  assign n941 = ~n939 & ~n940;
  assign n942 = n793 & n941;
  assign n943 = n938 & n942;
  assign n944 = ~n489 & ~n836;
  assign n945 = ~n772 & ~n826;
  assign n946 = n944 & n945;
  assign n947 = n858 & n946;
  assign n948 = n943 & n947;
  assign n949 = n101 & n402;
  assign n950 = n31 & n545;
  assign n951 = ~i_3_ & n844;
  assign n952 = ~n950 & ~n951;
  assign n953 = n128 & ~n952;
  assign n954 = n95 & n374;
  assign n955 = ~n953 & ~n954;
  assign n956 = ~n949 & n955;
  assign n957 = n32 & n85;
  assign n958 = n35 & n957;
  assign n959 = ~n777 & ~n958;
  assign n960 = ~n754 & n959;
  assign n961 = n956 & n960;
  assign n962 = n948 & n961;
  assign n963 = n95 & n111;
  assign n964 = n120 & n963;
  assign n965 = ~n544 & ~n964;
  assign n966 = n809 & n965;
  assign n967 = ~n785 & n966;
  assign n968 = n77 & n713;
  assign n969 = ~n837 & ~n968;
  assign n970 = ~n313 & n969;
  assign n971 = n65 & n970;
  assign n972 = n34 & n378;
  assign n973 = n48 & n68;
  assign n974 = ~n972 & ~n973;
  assign n975 = n35 & n259;
  assign n976 = n974 & ~n975;
  assign n977 = n115 & n136;
  assign n978 = n53 & n414;
  assign n979 = ~n977 & ~n978;
  assign n980 = n53 & n240;
  assign n981 = ~n821 & ~n980;
  assign n982 = n979 & n981;
  assign n983 = n976 & n982;
  assign n984 = n381 & n983;
  assign n985 = n971 & n984;
  assign n986 = n967 & n985;
  assign n987 = n530 & n986;
  assign n988 = n962 & n987;
  assign n989 = n653 & n988;
  assign o_5_ = ~n936 | ~n989;
  assign n991 = ~n135 & n925;
  assign n992 = n248 & ~n519;
  assign n993 = ~n313 & n992;
  assign n994 = n224 & n993;
  assign n995 = n991 & n994;
  assign n996 = n597 & n742;
  assign n997 = ~n129 & ~n996;
  assign n998 = ~i_3_ & ~n997;
  assign n999 = n434 & ~n998;
  assign n1000 = n117 & n435;
  assign n1001 = n67 & n287;
  assign n1002 = n35 & n1001;
  assign n1003 = ~n1000 & ~n1002;
  assign n1004 = ~n185 & n1003;
  assign n1005 = ~n885 & n1004;
  assign n1006 = n999 & n1005;
  assign n1007 = ~n470 & ~n817;
  assign n1008 = ~n484 & ~n515;
  assign n1009 = n400 & n1008;
  assign n1010 = n1007 & n1009;
  assign n1011 = n1006 & n1010;
  assign n1012 = ~n194 & ~n564;
  assign n1013 = ~n486 & ~n579;
  assign n1014 = n96 & n127;
  assign n1015 = n1013 & ~n1014;
  assign n1016 = n38 & n339;
  assign n1017 = ~n363 & ~n1016;
  assign n1018 = n1015 & n1017;
  assign n1019 = n1012 & n1018;
  assign n1020 = n78 & n121;
  assign n1021 = n79 & n219;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = n719 & n1022;
  assign n1024 = n698 & n1023;
  assign n1025 = n1019 & n1024;
  assign n1026 = n1011 & n1025;
  assign n1027 = n645 & n782;
  assign n1028 = n1026 & n1027;
  assign n1029 = n995 & n1028;
  assign n1030 = ~n561 & ~n889;
  assign n1031 = ~n334 & n1030;
  assign n1032 = ~n266 & n1031;
  assign n1033 = ~n44 & ~n713;
  assign n1034 = n30 & ~n1033;
  assign n1035 = n53 & n136;
  assign n1036 = n79 & n374;
  assign n1037 = n57 & n755;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = ~n1035 & n1038;
  assign n1040 = ~n1034 & n1039;
  assign n1041 = n1032 & n1040;
  assign n1042 = n95 & n869;
  assign n1043 = ~n55 & ~n198;
  assign n1044 = ~n1042 & n1043;
  assign n1045 = n504 & n1044;
  assign n1046 = n35 & n240;
  assign n1047 = n34 & n184;
  assign n1048 = n53 & n692;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = ~n1046 & n1049;
  assign n1051 = n706 & n1050;
  assign n1052 = n1045 & n1051;
  assign n1053 = n1041 & n1052;
  assign n1054 = n90 & n305;
  assign n1055 = n51 & n245;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n86 & n333;
  assign n1058 = n36 & n127;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = n53 & n139;
  assign n1061 = ~n373 & ~n1060;
  assign n1062 = n1059 & n1061;
  assign n1063 = n1056 & n1062;
  assign n1064 = n40 & n41;
  assign n1065 = n31 & n1064;
  assign n1066 = n90 & n374;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~n63 & ~n376;
  assign n1069 = n1067 & n1068;
  assign n1070 = i_1_ & n276;
  assign n1071 = ~n325 & ~n1070;
  assign n1072 = n48 & ~n1071;
  assign n1073 = ~n323 & ~n1072;
  assign n1074 = n1069 & n1073;
  assign n1075 = n1063 & n1074;
  assign n1076 = n170 & n1075;
  assign n1077 = n1053 & n1076;
  assign n1078 = n548 & n840;
  assign n1079 = n66 & n531;
  assign n1080 = ~n580 & ~n1079;
  assign n1081 = ~n375 & n1080;
  assign n1082 = ~n826 & n1081;
  assign n1083 = n1078 & n1082;
  assign n1084 = n815 & n1083;
  assign n1085 = n1077 & n1084;
  assign n1086 = n209 & n288;
  assign n1087 = ~n301 & ~n1086;
  assign n1088 = n255 & n439;
  assign n1089 = n1087 & ~n1088;
  assign n1090 = ~n900 & n1089;
  assign n1091 = n86 & n96;
  assign n1092 = n1090 & ~n1091;
  assign n1093 = n979 & n1092;
  assign n1094 = n880 & n1093;
  assign n1095 = n276 & n531;
  assign n1096 = ~n473 & ~n1095;
  assign n1097 = n308 & n1096;
  assign n1098 = ~n512 & ~n568;
  assign n1099 = n1097 & n1098;
  assign n1100 = n1094 & n1099;
  assign n1101 = n1085 & n1100;
  assign o_6_ = ~n1029 | ~n1101;
  assign n1103 = n849 & n1029;
  assign n1104 = n35 & n692;
  assign n1105 = ~n346 & ~n1104;
  assign n1106 = ~n50 & ~n375;
  assign n1107 = ~n226 & n1106;
  assign n1108 = n1105 & n1107;
  assign n1109 = n51 & n120;
  assign n1110 = n115 & n1109;
  assign n1111 = ~i_0_ & n324;
  assign n1112 = n134 & n1111;
  assign n1113 = n40 & n1112;
  assign n1114 = ~n1110 & ~n1113;
  assign n1115 = ~n344 & ~n474;
  assign n1116 = n1114 & n1115;
  assign n1117 = ~n525 & n1116;
  assign n1118 = n1108 & n1117;
  assign n1119 = n667 & n1118;
  assign n1120 = n49 & n77;
  assign n1121 = n48 & n316;
  assign n1122 = n95 & n113;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = n127 & n345;
  assign n1125 = n1123 & ~n1124;
  assign n1126 = ~n1120 & n1125;
  assign n1127 = n457 & n625;
  assign n1128 = n95 & n149;
  assign n1129 = n321 & ~n1128;
  assign n1130 = ~n975 & n1129;
  assign n1131 = n1127 & n1130;
  assign n1132 = n1126 & n1131;
  assign n1133 = n1119 & n1132;
  assign n1134 = n776 & n1133;
  assign n1135 = n94 & n1112;
  assign n1136 = ~n119 & ~n1135;
  assign n1137 = ~n524 & n1136;
  assign n1138 = n493 & n1137;
  assign n1139 = n1134 & n1138;
  assign n1140 = n47 & n240;
  assign n1141 = n30 & n578;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = n116 & n890;
  assign n1144 = n115 & n374;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = n1142 & n1145;
  assign n1147 = ~n521 & ~n707;
  assign n1148 = ~n261 & n1147;
  assign n1149 = n1146 & n1148;
  assign n1150 = n956 & n1149;
  assign n1151 = n932 & ~n940;
  assign n1152 = n557 & n1151;
  assign n1153 = n1150 & n1152;
  assign n1154 = i_6_ & n77;
  assign n1155 = n742 & n1154;
  assign n1156 = n255 & n1155;
  assign n1157 = n128 & n278;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = ~n559 & ~n595;
  assign n1160 = n1158 & n1159;
  assign n1161 = n1153 & n1160;
  assign n1162 = n1139 & n1161;
  assign o_7_ = ~n1103 | ~n1162;
  assign n1164 = n237 & n414;
  assign n1165 = ~n582 & ~n1164;
  assign n1166 = ~n241 & n1165;
  assign n1167 = n79 & n259;
  assign n1168 = ~n489 & ~n1167;
  assign n1169 = ~n522 & n1168;
  assign n1170 = n1166 & n1169;
  assign n1171 = n60 & n240;
  assign n1172 = n40 & n1155;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n494 & n1173;
  assign n1175 = n1170 & n1174;
  assign n1176 = ~n137 & ~n364;
  assign n1177 = ~n409 & n1176;
  assign n1178 = ~n122 & n1177;
  assign n1179 = n605 & n1178;
  assign n1180 = n1175 & n1179;
  assign n1181 = n1053 & n1180;
  assign n1182 = n852 & n1181;
  assign n1183 = n112 & n209;
  assign n1184 = i_6_ & n1183;
  assign n1185 = n78 & n86;
  assign n1186 = n33 & n1185;
  assign n1187 = ~n1184 & ~n1186;
  assign n1188 = n255 & n1183;
  assign n1189 = ~n588 & ~n1188;
  assign n1190 = n1187 & n1189;
  assign n1191 = n910 & n1190;
  assign n1192 = n1019 & n1191;
  assign n1193 = n48 & n402;
  assign n1194 = n71 & n1109;
  assign n1195 = n35 & n402;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1193 & n1196;
  assign n1198 = ~n291 & ~n431;
  assign n1199 = ~n495 & ~n920;
  assign n1200 = n1198 & n1199;
  assign n1201 = n60 & n151;
  assign n1202 = ~n885 & ~n1201;
  assign n1203 = n1200 & n1202;
  assign n1204 = n1197 & n1203;
  assign n1205 = n66 & n450;
  assign n1206 = n267 & n292;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = i_1_ & ~i_3_;
  assign n1209 = n199 & n1208;
  assign n1210 = n1207 & ~n1209;
  assign n1211 = n965 & n1210;
  assign n1212 = n1204 & n1211;
  assign n1213 = n1192 & n1212;
  assign n1214 = n1133 & n1213;
  assign o_8_ = ~n1182 | ~n1214;
  assign n1216 = n193 & n500;
  assign n1217 = n819 & n1160;
  assign n1218 = n413 & n1190;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1083 & n1219;
  assign n1221 = n36 & n77;
  assign n1222 = ~i_1_ & n324;
  assign n1223 = n844 & n1222;
  assign n1224 = ~n1221 & ~n1223;
  assign n1225 = n855 & n1224;
  assign n1226 = n1126 & n1225;
  assign n1227 = ~n695 & ~n1167;
  assign n1228 = n138 & n1227;
  assign n1229 = ~n685 & n1228;
  assign n1230 = ~n770 & ~n1141;
  assign n1231 = ~n1021 & n1230;
  assign n1232 = n1229 & n1231;
  assign n1233 = n1226 & n1232;
  assign n1234 = ~n553 & n1012;
  assign n1235 = n32 & n274;
  assign n1236 = n1050 & ~n1235;
  assign n1237 = n1234 & n1236;
  assign n1238 = n1233 & n1237;
  assign n1239 = n1056 & n1114;
  assign n1240 = n52 & n366;
  assign n1241 = n120 & n351;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = n35 & n1109;
  assign n1244 = n1242 & ~n1243;
  assign n1245 = n1239 & n1244;
  assign n1246 = n115 & n1222;
  assign n1247 = ~n578 & ~n1246;
  assign n1248 = ~i_5_ & ~n1247;
  assign n1249 = n804 & ~n1248;
  assign n1250 = n740 & n1249;
  assign n1251 = n1245 & n1250;
  assign n1252 = n38 & n62;
  assign n1253 = n127 & n359;
  assign n1254 = n47 & n1253;
  assign n1255 = ~n1252 & ~n1254;
  assign n1256 = ~n1000 & ~n1195;
  assign n1257 = n1255 & n1256;
  assign n1258 = ~n693 & ~n1035;
  assign n1259 = n1257 & n1258;
  assign n1260 = n574 & n1259;
  assign n1261 = n1251 & n1260;
  assign n1262 = n1238 & n1261;
  assign n1263 = n1220 & n1262;
  assign n1264 = n936 & n1263;
  assign o_9_ = ~n1216 | ~n1264;
  assign n1266 = n423 & n1208;
  assign n1267 = ~n828 & ~n1266;
  assign n1268 = n1173 & n1267;
  assign n1269 = ~n613 & ~n870;
  assign n1270 = n734 & n1269;
  assign n1271 = n1268 & n1270;
  assign n1272 = n896 & n1271;
  assign n1273 = n1238 & n1272;
  assign n1274 = ~n507 & ~n712;
  assign n1275 = n51 & ~n1274;
  assign n1276 = ~n873 & ~n1275;
  assign n1277 = ~n750 & n1276;
  assign n1278 = n639 & n1277;
  assign n1279 = n35 & n367;
  assign n1280 = ~n684 & ~n1279;
  assign n1281 = n1087 & n1280;
  assign n1282 = n133 & n1281;
  assign n1283 = ~i_1_ & n179;
  assign n1284 = i_1_ & n255;
  assign n1285 = ~i_4_ & n1284;
  assign n1286 = ~n1283 & ~n1285;
  assign n1287 = n73 & ~n1286;
  assign n1288 = n32 & n265;
  assign n1289 = ~n1037 & ~n1288;
  assign n1290 = ~n1135 & n1289;
  assign n1291 = n59 & n154;
  assign n1292 = ~n1128 & ~n1291;
  assign n1293 = ~n875 & ~n1020;
  assign n1294 = n1292 & n1293;
  assign n1295 = n1290 & n1294;
  assign n1296 = ~n1287 & n1295;
  assign n1297 = n1282 & n1296;
  assign n1298 = n948 & n1297;
  assign n1299 = n1278 & n1298;
  assign n1300 = n446 & n1299;
  assign o_10_ = ~n1273 | ~n1300;
  assign n1302 = ~i_2_ & n208;
  assign n1303 = ~n1144 & ~n1302;
  assign n1304 = ~n222 & ~n903;
  assign n1305 = n1303 & n1304;
  assign n1306 = n38 & n1222;
  assign n1307 = ~n210 & ~n1306;
  assign n1308 = n35 & ~n1307;
  assign n1309 = n131 & ~n1308;
  assign n1310 = n1305 & n1309;
  assign n1311 = n42 & n549;
  assign n1312 = ~n196 & ~n1311;
  assign n1313 = ~n230 & ~n410;
  assign n1314 = n1123 & n1313;
  assign n1315 = n1312 & n1314;
  assign n1316 = n1310 & n1315;
  assign n1317 = ~n881 & n969;
  assign n1318 = ~n160 & ~n642;
  assign n1319 = n1317 & n1318;
  assign n1320 = n1204 & n1319;
  assign n1321 = n1316 & n1320;
  assign n1322 = n563 & n1277;
  assign n1323 = n330 & n1322;
  assign n1324 = n476 & n1323;
  assign n1325 = n1321 & n1324;
  assign n1326 = ~n306 & ~n917;
  assign n1327 = ~n409 & n1326;
  assign n1328 = n186 & n208;
  assign n1329 = ~i_6_ & n1328;
  assign n1330 = ~n711 & ~n1329;
  assign n1331 = n676 & n1330;
  assign n1332 = n1327 & n1331;
  assign n1333 = ~n646 & ~n807;
  assign n1334 = ~n246 & ~n633;
  assign n1335 = n1333 & n1334;
  assign n1336 = ~n836 & n1335;
  assign n1337 = n1332 & n1336;
  assign n1338 = n83 & ~n977;
  assign n1339 = ~n519 & n656;
  assign n1340 = n1338 & n1339;
  assign n1341 = n1337 & n1340;
  assign n1342 = n338 & ~n1046;
  assign n1343 = n449 & n1137;
  assign n1344 = n1108 & n1343;
  assign n1345 = n1342 & n1344;
  assign n1346 = n1341 & n1345;
  assign n1347 = ~n736 & n1346;
  assign n1348 = n1325 & n1347;
  assign n1349 = ~n843 & ~n919;
  assign n1350 = ~n225 & n1349;
  assign n1351 = n43 & n352;
  assign n1352 = ~n629 & ~n1351;
  assign n1353 = n1350 & n1352;
  assign n1354 = ~n228 & ~n664;
  assign n1355 = ~n218 & ~n859;
  assign n1356 = ~n732 & ~n980;
  assign n1357 = n1355 & n1356;
  assign n1358 = n1354 & n1357;
  assign n1359 = n1353 & n1358;
  assign n1360 = ~n532 & n1359;
  assign n1361 = ~n1184 & n1360;
  assign n1362 = ~n63 & n1361;
  assign o_11_ = ~n1348 | ~n1362;
  assign n1364 = ~n490 & ~n978;
  assign n1365 = ~n502 & ~n760;
  assign n1366 = ~n1302 & n1365;
  assign n1367 = n95 & n305;
  assign n1368 = ~n415 & ~n1367;
  assign n1369 = ~n480 & n1368;
  assign n1370 = n872 & n1369;
  assign n1371 = n1366 & n1370;
  assign n1372 = ~n397 & ~n602;
  assign n1373 = ~n794 & n1372;
  assign n1374 = ~n636 & n1373;
  assign n1375 = ~n658 & n1374;
  assign n1376 = n1371 & n1375;
  assign n1377 = n1063 & n1234;
  assign n1378 = ~n45 & n523;
  assign n1379 = n284 & n1378;
  assign n1380 = ~n975 & ~n1184;
  assign n1381 = ~n241 & ~n1036;
  assign n1382 = ~n174 & n1381;
  assign n1383 = n1380 & n1382;
  assign n1384 = n1379 & n1383;
  assign n1385 = n1377 & n1384;
  assign n1386 = n1376 & n1385;
  assign n1387 = n1364 & n1386;
  assign n1388 = n208 & n963;
  assign n1389 = ~n144 & ~n821;
  assign n1390 = ~n1388 & n1389;
  assign n1391 = ~n571 & ~n817;
  assign n1392 = ~n800 & ~n1035;
  assign n1393 = ~n659 & ~n954;
  assign n1394 = n1392 & n1393;
  assign n1395 = n1391 & n1394;
  assign n1396 = ~n285 & ~n454;
  assign n1397 = ~n407 & n1396;
  assign n1398 = n1395 & n1397;
  assign n1399 = n1390 & n1398;
  assign n1400 = ~n293 & ~n1164;
  assign n1401 = ~n764 & n1400;
  assign n1402 = n1399 & n1401;
  assign n1403 = n1346 & n1402;
  assign o_12_ = ~n1387 | ~n1403;
  assign n1405 = n420 & n748;
  assign n1406 = ~n242 & ~n481;
  assign n1407 = ~n261 & ~n486;
  assign n1408 = ~n1157 & n1407;
  assign n1409 = n1406 & n1408;
  assign n1410 = ~n1042 & n1280;
  assign n1411 = n1409 & n1410;
  assign n1412 = ~n854 & ~n1243;
  assign n1413 = n112 & n208;
  assign n1414 = ~i_6_ & n1413;
  assign n1415 = n1412 & ~n1414;
  assign n1416 = n71 & n139;
  assign n1417 = ~n164 & ~n1416;
  assign n1418 = ~n189 & n1417;
  assign n1419 = n827 & n1418;
  assign n1420 = n1415 & n1419;
  assign n1421 = n1411 & n1420;
  assign n1422 = ~n669 & ~n704;
  assign n1423 = ~n505 & n1422;
  assign n1424 = ~n534 & ~n738;
  assign n1425 = ~n714 & n1424;
  assign n1426 = n1423 & n1425;
  assign n1427 = n586 & n1426;
  assign n1428 = n1421 & n1427;
  assign n1429 = n1405 & n1428;
  assign n1430 = n1168 & n1386;
  assign n1431 = n1429 & n1430;
  assign n1432 = ~n1291 & n1359;
  assign n1433 = ~n1095 & n1432;
  assign n1434 = ~n842 & n1433;
  assign o_13_ = ~n1431 | ~n1434;
  assign n1436 = ~n155 & n1399;
  assign n1437 = n237 & n1413;
  assign n1438 = n1436 & ~n1437;
  assign n1439 = n1429 & n1438;
  assign n1440 = ~n1088 & ~n1206;
  assign n1441 = n1325 & n1440;
  assign o_14_ = ~n1439 | ~n1441;
  assign n1443 = ~n795 & n1380;
  assign n1444 = ~n1329 & n1443;
  assign n1445 = n1382 & n1444;
  assign n1446 = ~n260 & ~n1388;
  assign n1447 = ~n1110 & n1446;
  assign n1448 = ~n71 & ~n100;
  assign n1449 = n240 & n1448;
  assign n1450 = ~n603 & ~n1449;
  assign n1451 = n1447 & n1450;
  assign n1452 = n1445 & n1451;
  assign n1453 = ~n902 & ~n954;
  assign n1454 = ~n451 & ~n841;
  assign n1455 = ~n807 & ~n873;
  assign n1456 = n1454 & n1455;
  assign n1457 = n71 & n219;
  assign n1458 = ~n1066 & ~n1457;
  assign n1459 = ~n939 & n1458;
  assign n1460 = n1456 & n1459;
  assign n1461 = ~n211 & ~n579;
  assign n1462 = n536 & n1461;
  assign n1463 = n1366 & n1462;
  assign n1464 = n1460 & n1463;
  assign n1465 = n1453 & n1464;
  assign o_15_ = ~n1452 | ~n1465;
  assign n1467 = ~n873 & ~n1302;
  assign n1468 = ~n770 & ~n949;
  assign n1469 = ~n183 & n1468;
  assign n1470 = n1467 & n1469;
  assign n1471 = ~n695 & ~n875;
  assign n1472 = n1470 & n1471;
  assign o_16_ = ~n1452 | ~n1472;
  assign n1474 = ~n142 & ~n836;
  assign n1475 = n1470 & n1474;
  assign n1476 = n1444 & n1453;
  assign o_17_ = ~n1475 | ~n1476;
  assign n1478 = n1471 & n1474;
  assign n1479 = ~n1414 & n1478;
  assign n1480 = ~n1437 & n1479;
  assign o_18_ = ~n1464 | ~n1480;
  assign o_0_ = 1'b0;
endmodule


