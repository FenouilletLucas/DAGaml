// Benchmark "t481" written by ABC on Tue May 16 16:07:52 2017

module t481 ( 
    v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9,
    \v16.0   );
  input  v10, v11, v12, v13, v14, v15, v0, v1, v2, v3, v4, v5, v6, v7,
    v8, v9;
  output \v16.0 ;
  wire n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639;
  assign n18 = v10 & v9;
  assign n19 = ~v12 & v13;
  assign n20 = v15 & n19;
  assign n21 = ~v5 & v7;
  assign n22 = ~v8 & n21;
  assign n23 = v0 & v2;
  assign n24 = ~v3 & n23;
  assign n25 = n22 & n24;
  assign n26 = n20 & n25;
  assign n27 = ~v11 & n26;
  assign n28 = n18 & n27;
  assign n29 = ~v1 & v2;
  assign n30 = ~v3 & n29;
  assign n31 = n22 & n30;
  assign n32 = n20 & n31;
  assign n33 = ~v11 & n32;
  assign n34 = n18 & n33;
  assign n35 = v5 & v6;
  assign n36 = ~v4 & n24;
  assign n37 = ~v8 & v9;
  assign n38 = v10 & n37;
  assign n39 = ~v11 & n38;
  assign n40 = n20 & n39;
  assign n41 = n36 & n40;
  assign n42 = ~v7 & n41;
  assign n43 = n35 & n42;
  assign n44 = ~v4 & n30;
  assign n45 = ~v7 & n35;
  assign n46 = n44 & n45;
  assign n47 = n40 & n46;
  assign n48 = ~n43 & ~n47;
  assign n49 = ~n34 & n48;
  assign n50 = ~n28 & n49;
  assign n51 = v4 & ~v6;
  assign n52 = ~v8 & n51;
  assign n53 = n24 & n52;
  assign n54 = n20 & n53;
  assign n55 = ~v11 & n54;
  assign n56 = n18 & n55;
  assign n57 = n30 & n52;
  assign n58 = n20 & n57;
  assign n59 = ~v11 & n58;
  assign n60 = n18 & n59;
  assign n61 = ~v5 & ~v8;
  assign n62 = ~v6 & n61;
  assign n63 = n24 & n62;
  assign n64 = n20 & n63;
  assign n65 = ~v11 & n64;
  assign n66 = n18 & n65;
  assign n67 = n30 & n62;
  assign n68 = n20 & n67;
  assign n69 = ~v11 & n68;
  assign n70 = n18 & n69;
  assign n71 = ~n66 & ~n70;
  assign n72 = ~n60 & n71;
  assign n73 = ~n56 & n72;
  assign n74 = ~v0 & v1;
  assign n75 = v3 & n74;
  assign n76 = ~v4 & n75;
  assign n77 = ~v14 & n19;
  assign n78 = n39 & n77;
  assign n79 = n76 & n78;
  assign n80 = ~v7 & n79;
  assign n81 = n35 & n80;
  assign n82 = ~v2 & n74;
  assign n83 = ~v4 & n82;
  assign n84 = n45 & n83;
  assign n85 = n39 & n84;
  assign n86 = ~v14 & n85;
  assign n87 = n19 & n86;
  assign n88 = n62 & n82;
  assign n89 = n77 & n88;
  assign n90 = ~v11 & n89;
  assign n91 = n18 & n90;
  assign n92 = ~v11 & n18;
  assign n93 = n77 & n92;
  assign n94 = v4 & v7;
  assign n95 = ~v8 & n94;
  assign n96 = n75 & n95;
  assign n97 = n93 & n96;
  assign n98 = n20 & n92;
  assign n99 = n24 & n95;
  assign n100 = n98 & n99;
  assign n101 = n30 & n95;
  assign n102 = n98 & n101;
  assign n103 = n82 & n95;
  assign n104 = n93 & n103;
  assign n105 = ~n102 & ~n104;
  assign n106 = ~n100 & n105;
  assign n107 = ~n97 & n106;
  assign n108 = ~n91 & n107;
  assign n109 = ~n87 & n108;
  assign n110 = ~n81 & n109;
  assign n111 = n30 & n93;
  assign n112 = n52 & n111;
  assign n113 = ~v8 & n24;
  assign n114 = ~v5 & n113;
  assign n115 = ~v6 & n114;
  assign n116 = n93 & n115;
  assign n117 = n62 & n111;
  assign n118 = n22 & n93;
  assign n119 = v3 & n118;
  assign n120 = n74 & n119;
  assign n121 = ~n117 & ~n120;
  assign n122 = ~n116 & n121;
  assign n123 = ~n112 & n122;
  assign n124 = n82 & n93;
  assign n125 = n22 & n124;
  assign n126 = n52 & n93;
  assign n127 = v3 & n126;
  assign n128 = n74 & n127;
  assign n129 = n52 & n124;
  assign n130 = n62 & n93;
  assign n131 = v3 & n130;
  assign n132 = n74 & n131;
  assign n133 = ~n129 & ~n132;
  assign n134 = ~n128 & n133;
  assign n135 = ~n125 & n134;
  assign n136 = n93 & n101;
  assign n137 = n25 & n93;
  assign n138 = n93 & n99;
  assign n139 = n31 & n77;
  assign n140 = ~v11 & n139;
  assign n141 = n18 & n140;
  assign n142 = n36 & n78;
  assign n143 = ~v7 & n142;
  assign n144 = n35 & n143;
  assign n145 = n39 & n46;
  assign n146 = ~v14 & n145;
  assign n147 = n19 & n146;
  assign n148 = n53 & n77;
  assign n149 = ~v11 & n148;
  assign n150 = n18 & n149;
  assign n151 = ~n147 & ~n150;
  assign n152 = ~n144 & n151;
  assign n153 = ~n141 & n152;
  assign n154 = ~n138 & n153;
  assign n155 = ~n137 & n154;
  assign n156 = ~n136 & n155;
  assign n157 = n135 & n156;
  assign n158 = n123 & n157;
  assign n159 = n110 & n158;
  assign n160 = n73 & n159;
  assign n161 = n50 & n160;
  assign n162 = n40 & n84;
  assign n163 = n20 & n96;
  assign n164 = ~v11 & n163;
  assign n165 = n18 & n164;
  assign n166 = n20 & n103;
  assign n167 = ~v11 & n166;
  assign n168 = n18 & n167;
  assign n169 = ~v10 & v8;
  assign n170 = ~v12 & n169;
  assign n171 = v7 & n24;
  assign n172 = v4 & n171;
  assign n173 = v13 & ~v14;
  assign n174 = n172 & n173;
  assign n175 = n170 & n174;
  assign n176 = ~n168 & ~n175;
  assign n177 = ~n165 & n176;
  assign n178 = ~n162 & n177;
  assign n179 = v7 & n30;
  assign n180 = v4 & n179;
  assign n181 = n173 & n180;
  assign n182 = n170 & n181;
  assign n183 = n170 & n173;
  assign n184 = n21 & n183;
  assign n185 = n24 & n184;
  assign n186 = n30 & n184;
  assign n187 = ~v4 & v5;
  assign n188 = v6 & n187;
  assign n189 = ~v7 & v8;
  assign n190 = ~v10 & n189;
  assign n191 = n77 & n190;
  assign n192 = n188 & n191;
  assign n193 = ~v3 & n192;
  assign n194 = n23 & n193;
  assign n195 = ~n186 & ~n194;
  assign n196 = ~n185 & n195;
  assign n197 = ~n182 & n196;
  assign n198 = n22 & n82;
  assign n199 = n20 & n198;
  assign n200 = ~v11 & n199;
  assign n201 = n18 & n200;
  assign n202 = n52 & n75;
  assign n203 = n20 & n202;
  assign n204 = ~v11 & n203;
  assign n205 = n18 & n204;
  assign n206 = n22 & n75;
  assign n207 = n20 & n206;
  assign n208 = ~v11 & n207;
  assign n209 = n18 & n208;
  assign n210 = n82 & n98;
  assign n211 = n52 & n210;
  assign n212 = n62 & n98;
  assign n213 = v3 & n212;
  assign n214 = n74 & n213;
  assign n215 = n62 & n210;
  assign n216 = n45 & n76;
  assign n217 = n39 & n216;
  assign n218 = v15 & n217;
  assign n219 = n19 & n218;
  assign n220 = ~n215 & ~n219;
  assign n221 = ~n214 & n220;
  assign n222 = ~n211 & n221;
  assign n223 = ~n209 & n222;
  assign n224 = ~n205 & n223;
  assign n225 = ~n201 & n224;
  assign n226 = ~v3 & v4;
  assign n227 = ~v6 & n226;
  assign n228 = n23 & n227;
  assign n229 = n173 & n228;
  assign n230 = n170 & n229;
  assign n231 = n30 & n51;
  assign n232 = n173 & n231;
  assign n233 = n170 & n232;
  assign n234 = n30 & n188;
  assign n235 = n190 & n234;
  assign n236 = n77 & n235;
  assign n237 = ~n233 & ~n236;
  assign n238 = ~n230 & n237;
  assign n239 = ~v5 & n24;
  assign n240 = ~v6 & n239;
  assign n241 = n173 & n240;
  assign n242 = n170 & n241;
  assign n243 = ~v5 & n30;
  assign n244 = ~v6 & n243;
  assign n245 = n173 & n244;
  assign n246 = n170 & n245;
  assign n247 = n21 & n75;
  assign n248 = n173 & n247;
  assign n249 = n170 & n248;
  assign n250 = n21 & n82;
  assign n251 = n173 & n250;
  assign n252 = n170 & n251;
  assign n253 = ~n249 & ~n252;
  assign n254 = ~n246 & n253;
  assign n255 = ~n242 & n254;
  assign n256 = n51 & n75;
  assign n257 = n173 & n256;
  assign n258 = n170 & n257;
  assign n259 = n51 & n82;
  assign n260 = n173 & n259;
  assign n261 = n170 & n260;
  assign n262 = ~v5 & n75;
  assign n263 = ~v6 & n262;
  assign n264 = n173 & n263;
  assign n265 = n170 & n264;
  assign n266 = ~v5 & n82;
  assign n267 = ~v6 & n266;
  assign n268 = n173 & n267;
  assign n269 = n170 & n268;
  assign n270 = ~n265 & ~n269;
  assign n271 = ~n261 & n270;
  assign n272 = ~n258 & n271;
  assign n273 = n75 & n188;
  assign n274 = n190 & n273;
  assign n275 = n77 & n274;
  assign n276 = n82 & n188;
  assign n277 = n190 & n276;
  assign n278 = n77 & n277;
  assign n279 = n75 & n94;
  assign n280 = n173 & n279;
  assign n281 = n170 & n280;
  assign n282 = v11 & v8;
  assign n283 = n77 & n282;
  assign n284 = n24 & n283;
  assign n285 = v7 & n284;
  assign n286 = v4 & n285;
  assign n287 = ~n281 & ~n286;
  assign n288 = ~n278 & n287;
  assign n289 = ~n275 & n288;
  assign n290 = n272 & n289;
  assign n291 = n255 & n290;
  assign n292 = n238 & n291;
  assign n293 = n225 & n292;
  assign n294 = n197 & n293;
  assign n295 = n178 & n294;
  assign n296 = v11 & ~v9;
  assign n297 = ~v12 & n296;
  assign n298 = v13 & n297;
  assign n299 = v15 & n298;
  assign n300 = n21 & n299;
  assign n301 = n24 & n300;
  assign n302 = n30 & n300;
  assign n303 = ~v7 & ~v9;
  assign n304 = v11 & n303;
  assign n305 = n20 & n304;
  assign n306 = n188 & n305;
  assign n307 = ~v3 & n306;
  assign n308 = n23 & n307;
  assign n309 = n29 & n307;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~n302 & n310;
  assign n312 = ~n301 & n311;
  assign n313 = n51 & n299;
  assign n314 = n24 & n313;
  assign n315 = n30 & n313;
  assign n316 = n24 & n299;
  assign n317 = ~v5 & n316;
  assign n318 = ~v6 & n317;
  assign n319 = n30 & n299;
  assign n320 = ~v5 & n319;
  assign n321 = ~v6 & n320;
  assign n322 = ~n318 & ~n321;
  assign n323 = ~n315 & n322;
  assign n324 = ~n314 & n323;
  assign n325 = v11 & n189;
  assign n326 = n77 & n325;
  assign n327 = n75 & n326;
  assign n328 = n188 & n327;
  assign n329 = n276 & n326;
  assign n330 = ~v12 & n282;
  assign n331 = ~v5 & ~v6;
  assign n332 = n82 & n331;
  assign n333 = n173 & n332;
  assign n334 = n330 & n333;
  assign n335 = n75 & n283;
  assign n336 = v7 & n335;
  assign n337 = v4 & n336;
  assign n338 = n82 & n283;
  assign n339 = v7 & n338;
  assign n340 = v4 & n339;
  assign n341 = v13 & v15;
  assign n342 = n297 & n341;
  assign n343 = n24 & n342;
  assign n344 = v7 & n343;
  assign n345 = v4 & n344;
  assign n346 = n30 & n342;
  assign n347 = v7 & n346;
  assign n348 = v4 & n347;
  assign n349 = ~n345 & ~n348;
  assign n350 = ~n340 & n349;
  assign n351 = ~n337 & n350;
  assign n352 = ~n334 & n351;
  assign n353 = ~n329 & n352;
  assign n354 = ~n328 & n353;
  assign n355 = n51 & n283;
  assign n356 = n30 & n355;
  assign n357 = n241 & n330;
  assign n358 = n283 & n331;
  assign n359 = n30 & n358;
  assign n360 = n21 & n283;
  assign n361 = n75 & n360;
  assign n362 = ~n359 & ~n361;
  assign n363 = ~n357 & n362;
  assign n364 = ~n356 & n363;
  assign n365 = n82 & n360;
  assign n366 = n75 & n355;
  assign n367 = n82 & n355;
  assign n368 = n264 & n330;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & n369;
  assign n371 = ~n365 & n370;
  assign n372 = n82 & n94;
  assign n373 = n173 & n372;
  assign n374 = n170 & n373;
  assign n375 = n24 & n360;
  assign n376 = n30 & n283;
  assign n377 = v7 & n376;
  assign n378 = v4 & n377;
  assign n379 = n21 & n30;
  assign n380 = n173 & n379;
  assign n381 = n330 & n380;
  assign n382 = n188 & n326;
  assign n383 = ~v3 & n382;
  assign n384 = n23 & n383;
  assign n385 = n234 & n326;
  assign n386 = n24 & n51;
  assign n387 = n173 & n386;
  assign n388 = n330 & n387;
  assign n389 = ~n385 & ~n388;
  assign n390 = ~n384 & n389;
  assign n391 = ~n381 & n390;
  assign n392 = ~n378 & n391;
  assign n393 = ~n375 & n392;
  assign n394 = ~n374 & n393;
  assign n395 = n371 & n394;
  assign n396 = n364 & n395;
  assign n397 = n354 & n396;
  assign n398 = n324 & n397;
  assign n399 = n312 & n398;
  assign n400 = ~v12 & ~v9;
  assign n401 = ~v10 & n400;
  assign n402 = v13 & n401;
  assign n403 = v15 & n402;
  assign n404 = n51 & n403;
  assign n405 = n75 & n404;
  assign n406 = n82 & n404;
  assign n407 = n75 & n403;
  assign n408 = ~v5 & n407;
  assign n409 = ~v6 & n408;
  assign n410 = n82 & n403;
  assign n411 = ~v5 & n410;
  assign n412 = ~v6 & n411;
  assign n413 = ~n409 & ~n412;
  assign n414 = ~n406 & n413;
  assign n415 = ~n405 & n414;
  assign n416 = ~v10 & ~v7;
  assign n417 = ~v9 & n416;
  assign n418 = n20 & n417;
  assign n419 = n75 & n418;
  assign n420 = n188 & n419;
  assign n421 = n188 & n418;
  assign n422 = ~v2 & n421;
  assign n423 = n74 & n422;
  assign n424 = n94 & n403;
  assign n425 = n75 & n424;
  assign n426 = v13 & n170;
  assign n427 = v15 & n426;
  assign n428 = n94 & n427;
  assign n429 = n24 & n428;
  assign n430 = ~n425 & ~n429;
  assign n431 = ~n423 & n430;
  assign n432 = ~n420 & n431;
  assign n433 = n24 & n404;
  assign n434 = n30 & n404;
  assign n435 = ~v3 & n421;
  assign n436 = n29 & n435;
  assign n437 = n240 & n401;
  assign n438 = v13 & n437;
  assign n439 = v15 & n438;
  assign n440 = n244 & n401;
  assign n441 = v13 & n440;
  assign n442 = v15 & n441;
  assign n443 = n247 & n401;
  assign n444 = v13 & n443;
  assign n445 = v15 & n444;
  assign n446 = ~v12 & n341;
  assign n447 = ~v9 & n446;
  assign n448 = ~v10 & n447;
  assign n449 = n21 & n448;
  assign n450 = n82 & n449;
  assign n451 = ~n445 & ~n450;
  assign n452 = ~n442 & n451;
  assign n453 = ~n439 & n452;
  assign n454 = ~n436 & n453;
  assign n455 = ~n434 & n454;
  assign n456 = ~n433 & n455;
  assign n457 = n21 & n342;
  assign n458 = n82 & n457;
  assign n459 = n256 & n297;
  assign n460 = v13 & n459;
  assign n461 = v15 & n460;
  assign n462 = n247 & n297;
  assign n463 = v13 & n462;
  assign n464 = v15 & n463;
  assign n465 = ~n461 & ~n464;
  assign n466 = ~n458 & n465;
  assign n467 = n51 & n342;
  assign n468 = n82 & n467;
  assign n469 = n263 & n297;
  assign n470 = v13 & n469;
  assign n471 = v15 & n470;
  assign n472 = n267 & n297;
  assign n473 = v13 & n472;
  assign n474 = v15 & n473;
  assign n475 = n20 & n273;
  assign n476 = v11 & n475;
  assign n477 = n303 & n476;
  assign n478 = ~n474 & ~n477;
  assign n479 = ~n471 & n478;
  assign n480 = ~n468 & n479;
  assign n481 = n20 & n276;
  assign n482 = v11 & n481;
  assign n483 = n303 & n482;
  assign n484 = n75 & n342;
  assign n485 = v7 & n484;
  assign n486 = v4 & n485;
  assign n487 = n82 & n342;
  assign n488 = v7 & n487;
  assign n489 = v4 & n488;
  assign n490 = n24 & n448;
  assign n491 = v7 & n490;
  assign n492 = v4 & n491;
  assign n493 = ~n489 & ~n492;
  assign n494 = ~n486 & n493;
  assign n495 = ~n483 & n494;
  assign n496 = n30 & n448;
  assign n497 = v7 & n496;
  assign n498 = v4 & n497;
  assign n499 = ~v3 & ~v5;
  assign n500 = v7 & n499;
  assign n501 = n23 & n500;
  assign n502 = n401 & n501;
  assign n503 = v13 & n502;
  assign n504 = v15 & n503;
  assign n505 = n30 & n449;
  assign n506 = ~v10 & n20;
  assign n507 = ~v7 & n506;
  assign n508 = ~v9 & n507;
  assign n509 = n24 & n508;
  assign n510 = v6 & n509;
  assign n511 = n187 & n510;
  assign n512 = ~n505 & ~n511;
  assign n513 = ~n504 & n512;
  assign n514 = ~n498 & n513;
  assign n515 = n495 & n514;
  assign n516 = n480 & n515;
  assign n517 = n466 & n516;
  assign n518 = n456 & n517;
  assign n519 = n432 & n518;
  assign n520 = n415 & n519;
  assign n521 = n399 & n520;
  assign n522 = n295 & n521;
  assign n523 = n161 & n522;
  assign n524 = v13 & n330;
  assign n525 = v15 & n524;
  assign n526 = n21 & n525;
  assign n527 = n24 & n526;
  assign n528 = n341 & n379;
  assign n529 = n330 & n528;
  assign n530 = n24 & n188;
  assign n531 = n325 & n530;
  assign n532 = n20 & n531;
  assign n533 = n234 & n325;
  assign n534 = n20 & n533;
  assign n535 = ~n532 & ~n534;
  assign n536 = ~n529 & n535;
  assign n537 = ~n527 & n536;
  assign n538 = n51 & n525;
  assign n539 = n24 & n538;
  assign n540 = n231 & n341;
  assign n541 = n330 & n540;
  assign n542 = n24 & n525;
  assign n543 = ~v5 & n542;
  assign n544 = ~v6 & n543;
  assign n545 = n30 & n525;
  assign n546 = ~v5 & n545;
  assign n547 = ~v6 & n546;
  assign n548 = ~n544 & ~n547;
  assign n549 = ~n541 & n548;
  assign n550 = ~n539 & n549;
  assign n551 = n20 & n190;
  assign n552 = n75 & n551;
  assign n553 = n188 & n552;
  assign n554 = n188 & n551;
  assign n555 = ~v2 & n554;
  assign n556 = n74 & n555;
  assign n557 = n82 & n427;
  assign n558 = ~v5 & n557;
  assign n559 = ~v6 & n558;
  assign n560 = n170 & n341;
  assign n561 = n75 & n560;
  assign n562 = v7 & n561;
  assign n563 = v4 & n562;
  assign n564 = n20 & n282;
  assign n565 = n24 & n564;
  assign n566 = v7 & n565;
  assign n567 = v4 & n566;
  assign n568 = n30 & n564;
  assign n569 = v7 & n568;
  assign n570 = v4 & n569;
  assign n571 = n82 & n560;
  assign n572 = v7 & n571;
  assign n573 = v4 & n572;
  assign n574 = ~n570 & ~n573;
  assign n575 = ~n567 & n574;
  assign n576 = ~n563 & n575;
  assign n577 = ~n559 & n576;
  assign n578 = ~n556 & n577;
  assign n579 = ~n553 & n578;
  assign n580 = n82 & n448;
  assign n581 = v7 & n580;
  assign n582 = v4 & n581;
  assign n583 = n170 & n501;
  assign n584 = v13 & n583;
  assign n585 = v15 & n584;
  assign n586 = n30 & n560;
  assign n587 = v7 & n586;
  assign n588 = v4 & n587;
  assign n589 = ~n585 & ~n588;
  assign n590 = ~n582 & n589;
  assign n591 = n21 & n560;
  assign n592 = n30 & n591;
  assign n593 = n190 & n530;
  assign n594 = v15 & n593;
  assign n595 = n19 & n594;
  assign n596 = v15 & n235;
  assign n597 = n19 & n596;
  assign n598 = n170 & n228;
  assign n599 = v13 & n598;
  assign n600 = v15 & n599;
  assign n601 = ~n597 & ~n600;
  assign n602 = ~n595 & n601;
  assign n603 = ~n592 & n602;
  assign n604 = n51 & n560;
  assign n605 = n30 & n604;
  assign n606 = n170 & n240;
  assign n607 = v13 & n606;
  assign n608 = v15 & n607;
  assign n609 = n170 & n244;
  assign n610 = v13 & n609;
  assign n611 = v15 & n610;
  assign n612 = n170 & n247;
  assign n613 = v13 & n612;
  assign n614 = v15 & n613;
  assign n615 = ~n611 & ~n614;
  assign n616 = ~n608 & n615;
  assign n617 = ~n605 & n616;
  assign n618 = n82 & n591;
  assign n619 = n170 & n256;
  assign n620 = v13 & n619;
  assign n621 = v15 & n620;
  assign n622 = n82 & n604;
  assign n623 = n170 & n263;
  assign n624 = v13 & n623;
  assign n625 = v15 & n624;
  assign n626 = ~n622 & ~n625;
  assign n627 = ~n621 & n626;
  assign n628 = ~n618 & n627;
  assign n629 = n617 & n628;
  assign n630 = n603 & n629;
  assign n631 = n590 & n630;
  assign n632 = n579 & n631;
  assign n633 = n550 & n632;
  assign n634 = n537 & n633;
  assign n635 = ~v13 & v14;
  assign n636 = ~v15 & n635;
  assign n637 = n202 & n636;
  assign n638 = ~v11 & n637;
  assign n639 = n18 & n638;
  assign n640 = n52 & n82;
  assign n641 = n636 & n640;
  assign n642 = ~v11 & n641;
  assign n643 = n18 & n642;
  assign n644 = n62 & n75;
  assign n645 = n636 & n644;
  assign n646 = ~v11 & n645;
  assign n647 = n18 & n646;
  assign n648 = n88 & n636;
  assign n649 = ~v11 & n648;
  assign n650 = n18 & n649;
  assign n651 = ~n647 & ~n650;
  assign n652 = ~n643 & n651;
  assign n653 = ~n639 & n652;
  assign n654 = n39 & n636;
  assign n655 = n76 & n654;
  assign n656 = ~v7 & n655;
  assign n657 = n35 & n656;
  assign n658 = ~v15 & n85;
  assign n659 = n635 & n658;
  assign n660 = n92 & n636;
  assign n661 = n75 & n660;
  assign n662 = ~v8 & n661;
  assign n663 = n94 & n662;
  assign n664 = v12 & v14;
  assign n665 = ~v15 & n664;
  assign n666 = n99 & n665;
  assign n667 = ~v11 & n666;
  assign n668 = n18 & n667;
  assign n669 = ~n663 & ~n668;
  assign n670 = ~n659 & n669;
  assign n671 = ~n657 & n670;
  assign n672 = n53 & n636;
  assign n673 = ~v11 & n672;
  assign n674 = n18 & n673;
  assign n675 = n57 & n636;
  assign n676 = ~v11 & n675;
  assign n677 = n18 & n676;
  assign n678 = ~v15 & n145;
  assign n679 = n635 & n678;
  assign n680 = n115 & n660;
  assign n681 = n30 & n660;
  assign n682 = n62 & n681;
  assign n683 = n22 & n660;
  assign n684 = v3 & n683;
  assign n685 = n74 & n684;
  assign n686 = n82 & n660;
  assign n687 = n22 & n686;
  assign n688 = ~n685 & ~n687;
  assign n689 = ~n682 & n688;
  assign n690 = ~n680 & n689;
  assign n691 = ~n679 & n690;
  assign n692 = ~n677 & n691;
  assign n693 = ~n674 & n692;
  assign n694 = n21 & n564;
  assign n695 = n82 & n694;
  assign n696 = n256 & n330;
  assign n697 = v13 & n696;
  assign n698 = v15 & n697;
  assign n699 = n247 & n330;
  assign n700 = v13 & n699;
  assign n701 = v15 & n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = ~n695 & n702;
  assign n704 = n51 & n564;
  assign n705 = n82 & n704;
  assign n706 = n263 & n330;
  assign n707 = v13 & n706;
  assign n708 = v15 & n707;
  assign n709 = n267 & n330;
  assign n710 = v13 & n709;
  assign n711 = v15 & n710;
  assign n712 = n20 & n325;
  assign n713 = n273 & n712;
  assign n714 = ~n711 & ~n713;
  assign n715 = ~n708 & n714;
  assign n716 = ~n705 & n715;
  assign n717 = n276 & n712;
  assign n718 = n75 & n564;
  assign n719 = v7 & n718;
  assign n720 = v4 & n719;
  assign n721 = n82 & n564;
  assign n722 = v7 & n721;
  assign n723 = v4 & n722;
  assign n724 = n99 & n660;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n720 & n725;
  assign n727 = ~n717 & n726;
  assign n728 = n101 & n660;
  assign n729 = n25 & n660;
  assign n730 = n22 & n681;
  assign n731 = n36 & n654;
  assign n732 = n45 & n731;
  assign n733 = ~n730 & ~n732;
  assign n734 = ~n729 & n733;
  assign n735 = ~n728 & n734;
  assign n736 = n727 & n735;
  assign n737 = n716 & n736;
  assign n738 = n703 & n737;
  assign n739 = n693 & n738;
  assign n740 = n671 & n739;
  assign n741 = n653 & n740;
  assign n742 = n57 & n665;
  assign n743 = ~v11 & n742;
  assign n744 = n18 & n743;
  assign n745 = n63 & n665;
  assign n746 = ~v11 & n745;
  assign n747 = n18 & n746;
  assign n748 = n67 & n665;
  assign n749 = ~v11 & n748;
  assign n750 = n18 & n749;
  assign n751 = n206 & n665;
  assign n752 = ~v11 & n751;
  assign n753 = n18 & n752;
  assign n754 = ~n750 & ~n753;
  assign n755 = ~n747 & n754;
  assign n756 = ~n744 & n755;
  assign n757 = n198 & n665;
  assign n758 = ~v11 & n757;
  assign n759 = n18 & n758;
  assign n760 = n202 & n665;
  assign n761 = ~v11 & n760;
  assign n762 = n18 & n761;
  assign n763 = n640 & n665;
  assign n764 = ~v11 & n763;
  assign n765 = n18 & n764;
  assign n766 = n644 & n665;
  assign n767 = ~v11 & n766;
  assign n768 = n18 & n767;
  assign n769 = ~n765 & ~n768;
  assign n770 = ~n762 & n769;
  assign n771 = ~n759 & n770;
  assign n772 = n103 & n636;
  assign n773 = ~v11 & n772;
  assign n774 = n18 & n773;
  assign n775 = n25 & n665;
  assign n776 = ~v11 & n775;
  assign n777 = n18 & n776;
  assign n778 = n101 & n665;
  assign n779 = ~v11 & n778;
  assign n780 = n18 & n779;
  assign n781 = n92 & n665;
  assign n782 = n30 & n781;
  assign n783 = n22 & n782;
  assign n784 = n39 & n665;
  assign n785 = n36 & n784;
  assign n786 = n45 & n785;
  assign n787 = n44 & n784;
  assign n788 = n45 & n787;
  assign n789 = n53 & n781;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n786 & n790;
  assign n792 = ~n783 & n791;
  assign n793 = ~n780 & n792;
  assign n794 = ~n777 & n793;
  assign n795 = ~n774 & n794;
  assign n796 = n173 & n501;
  assign n797 = n297 & n796;
  assign n798 = n297 & n380;
  assign n799 = n77 & n530;
  assign n800 = v11 & n799;
  assign n801 = n303 & n800;
  assign n802 = n77 & n234;
  assign n803 = v11 & n802;
  assign n804 = n303 & n803;
  assign n805 = ~n801 & ~n804;
  assign n806 = ~n798 & n805;
  assign n807 = ~n797 & n806;
  assign n808 = n229 & n297;
  assign n809 = n232 & n297;
  assign n810 = n241 & n297;
  assign n811 = n245 & n297;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n809 & n812;
  assign n814 = ~n808 & n813;
  assign n815 = n76 & n784;
  assign n816 = n45 & n815;
  assign n817 = n83 & n784;
  assign n818 = n45 & n817;
  assign n819 = n82 & n781;
  assign n820 = n62 & n819;
  assign n821 = n96 & n665;
  assign n822 = ~v11 & n821;
  assign n823 = n18 & n822;
  assign n824 = n103 & n665;
  assign n825 = ~v11 & n824;
  assign n826 = n18 & n825;
  assign n827 = n174 & n297;
  assign n828 = n181 & n297;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n826 & n829;
  assign n831 = ~n823 & n830;
  assign n832 = ~n820 & n831;
  assign n833 = ~n818 & n832;
  assign n834 = ~n816 & n833;
  assign n835 = n814 & n834;
  assign n836 = n807 & n835;
  assign n837 = n795 & n836;
  assign n838 = n771 & n837;
  assign n839 = n756 & n838;
  assign n840 = n77 & n304;
  assign n841 = n188 & n840;
  assign n842 = ~v2 & n841;
  assign n843 = n74 & n842;
  assign n844 = v7 & n75;
  assign n845 = v4 & n844;
  assign n846 = n173 & n845;
  assign n847 = n297 & n846;
  assign n848 = ~v13 & n296;
  assign n849 = v14 & ~v15;
  assign n850 = n172 & n849;
  assign n851 = n848 & n850;
  assign n852 = n180 & n849;
  assign n853 = n848 & n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = ~n847 & n854;
  assign n856 = ~n843 & n855;
  assign n857 = v7 & n82;
  assign n858 = v4 & n857;
  assign n859 = n173 & n858;
  assign n860 = n297 & n859;
  assign n861 = n848 & n849;
  assign n862 = n21 & n861;
  assign n863 = n24 & n862;
  assign n864 = n30 & n862;
  assign n865 = n304 & n636;
  assign n866 = n188 & n865;
  assign n867 = ~v3 & n866;
  assign n868 = n23 & n867;
  assign n869 = ~n864 & ~n868;
  assign n870 = ~n863 & n869;
  assign n871 = ~n860 & n870;
  assign n872 = n173 & n297;
  assign n873 = n21 & n872;
  assign n874 = n82 & n873;
  assign n875 = n51 & n872;
  assign n876 = n75 & n875;
  assign n877 = n75 & n873;
  assign n878 = n260 & n297;
  assign n879 = n264 & n297;
  assign n880 = n268 & n297;
  assign n881 = n77 & n273;
  assign n882 = v11 & n881;
  assign n883 = n303 & n882;
  assign n884 = ~n880 & ~n883;
  assign n885 = ~n879 & n884;
  assign n886 = ~n878 & n885;
  assign n887 = ~n877 & n886;
  assign n888 = ~n876 & n887;
  assign n889 = ~n874 & n888;
  assign n890 = n228 & n849;
  assign n891 = n848 & n890;
  assign n892 = n231 & n849;
  assign n893 = n848 & n892;
  assign n894 = n234 & n636;
  assign n895 = v11 & n894;
  assign n896 = n303 & n895;
  assign n897 = ~n893 & ~n896;
  assign n898 = ~n891 & n897;
  assign n899 = n240 & n849;
  assign n900 = n848 & n899;
  assign n901 = n244 & n849;
  assign n902 = n848 & n901;
  assign n903 = n247 & n849;
  assign n904 = n848 & n903;
  assign n905 = n250 & n849;
  assign n906 = n848 & n905;
  assign n907 = ~n904 & ~n906;
  assign n908 = ~n902 & n907;
  assign n909 = ~n900 & n908;
  assign n910 = n256 & n849;
  assign n911 = n848 & n910;
  assign n912 = n259 & n849;
  assign n913 = n848 & n912;
  assign n914 = n263 & n849;
  assign n915 = n848 & n914;
  assign n916 = n267 & n849;
  assign n917 = n848 & n916;
  assign n918 = ~n915 & ~n917;
  assign n919 = ~n913 & n918;
  assign n920 = ~n911 & n919;
  assign n921 = n273 & n636;
  assign n922 = v11 & n921;
  assign n923 = n303 & n922;
  assign n924 = n276 & n636;
  assign n925 = v11 & n924;
  assign n926 = n303 & n925;
  assign n927 = n279 & n849;
  assign n928 = n848 & n927;
  assign n929 = n372 & n849;
  assign n930 = n848 & n929;
  assign n931 = ~n928 & ~n930;
  assign n932 = ~n926 & n931;
  assign n933 = ~n923 & n932;
  assign n934 = n920 & n933;
  assign n935 = n909 & n934;
  assign n936 = n898 & n935;
  assign n937 = n889 & n936;
  assign n938 = n871 & n937;
  assign n939 = n856 & n938;
  assign n940 = n839 & n939;
  assign n941 = n741 & n940;
  assign n942 = n634 & n941;
  assign n943 = ~v13 & n282;
  assign n944 = n21 & n24;
  assign n945 = n849 & n944;
  assign n946 = n943 & n945;
  assign n947 = n379 & n849;
  assign n948 = n943 & n947;
  assign n949 = n325 & n636;
  assign n950 = n188 & n949;
  assign n951 = ~v3 & n950;
  assign n952 = n23 & n951;
  assign n953 = n234 & n949;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~n948 & n954;
  assign n956 = ~n946 & n955;
  assign n957 = n386 & n849;
  assign n958 = n943 & n957;
  assign n959 = n892 & n943;
  assign n960 = n24 & n331;
  assign n961 = n849 & n960;
  assign n962 = n943 & n961;
  assign n963 = n30 & n331;
  assign n964 = n849 & n963;
  assign n965 = n943 & n964;
  assign n966 = ~n962 & ~n965;
  assign n967 = ~n959 & n966;
  assign n968 = ~n958 & n967;
  assign n969 = n190 & n636;
  assign n970 = n75 & n969;
  assign n971 = n188 & n970;
  assign n972 = n188 & n969;
  assign n973 = ~v2 & n972;
  assign n974 = n74 & n973;
  assign n975 = ~v13 & n169;
  assign n976 = n849 & n975;
  assign n977 = n82 & n976;
  assign n978 = ~v5 & n977;
  assign n979 = ~v6 & n978;
  assign n980 = n927 & n975;
  assign n981 = n282 & n636;
  assign n982 = n24 & n981;
  assign n983 = v7 & n982;
  assign n984 = v4 & n983;
  assign n985 = n30 & n981;
  assign n986 = v7 & n985;
  assign n987 = v4 & n986;
  assign n988 = n929 & n975;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~n984 & n989;
  assign n991 = ~n980 & n990;
  assign n992 = ~n979 & n991;
  assign n993 = ~n974 & n992;
  assign n994 = ~n971 & n993;
  assign n995 = n30 & n94;
  assign n996 = n849 & n995;
  assign n997 = n975 & n996;
  assign n998 = n501 & n849;
  assign n999 = n975 & n998;
  assign n1000 = n24 & n94;
  assign n1001 = n849 & n1000;
  assign n1002 = n975 & n1001;
  assign n1003 = ~n999 & ~n1002;
  assign n1004 = ~n997 & n1003;
  assign n1005 = n947 & n975;
  assign n1006 = n593 & n636;
  assign n1007 = n235 & n636;
  assign n1008 = n890 & n975;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~n1006 & n1009;
  assign n1011 = ~n1005 & n1010;
  assign n1012 = n892 & n975;
  assign n1013 = n899 & n975;
  assign n1014 = n901 & n975;
  assign n1015 = n903 & n975;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n1013 & n1016;
  assign n1018 = ~n1012 & n1017;
  assign n1019 = n905 & n975;
  assign n1020 = n910 & n975;
  assign n1021 = n912 & n975;
  assign n1022 = n914 & n975;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n1020 & n1023;
  assign n1025 = ~n1019 & n1024;
  assign n1026 = n1018 & n1025;
  assign n1027 = n1011 & n1026;
  assign n1028 = n1004 & n1027;
  assign n1029 = n994 & n1028;
  assign n1030 = n968 & n1029;
  assign n1031 = n956 & n1030;
  assign n1032 = v12 & n296;
  assign n1033 = n910 & n1032;
  assign n1034 = n912 & n1032;
  assign n1035 = n75 & n331;
  assign n1036 = n849 & n1035;
  assign n1037 = n1032 & n1036;
  assign n1038 = n332 & n849;
  assign n1039 = n1032 & n1038;
  assign n1040 = ~n1037 & ~n1039;
  assign n1041 = ~n1034 & n1040;
  assign n1042 = ~n1033 & n1041;
  assign n1043 = n304 & n665;
  assign n1044 = n75 & n1043;
  assign n1045 = n188 & n1044;
  assign n1046 = n188 & n1043;
  assign n1047 = ~v2 & n1046;
  assign n1048 = n74 & n1047;
  assign n1049 = n845 & n849;
  assign n1050 = n1032 & n1049;
  assign n1051 = n849 & n858;
  assign n1052 = n1032 & n1051;
  assign n1053 = ~n1050 & ~n1052;
  assign n1054 = ~n1048 & n1053;
  assign n1055 = ~n1045 & n1054;
  assign n1056 = n957 & n1032;
  assign n1057 = n892 & n1032;
  assign n1058 = ~v3 & n1046;
  assign n1059 = n29 & n1058;
  assign n1060 = n899 & n1032;
  assign n1061 = n901 & n1032;
  assign n1062 = n849 & n1032;
  assign n1063 = n21 & n1062;
  assign n1064 = n75 & n1063;
  assign n1065 = n82 & n1063;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~n1061 & n1066;
  assign n1068 = ~n1060 & n1067;
  assign n1069 = ~n1059 & n1068;
  assign n1070 = ~n1057 & n1069;
  assign n1071 = ~n1056 & n1070;
  assign n1072 = n276 & n949;
  assign n1073 = n75 & n981;
  assign n1074 = v7 & n1073;
  assign n1075 = v4 & n1074;
  assign n1076 = n82 & n981;
  assign n1077 = v7 & n1076;
  assign n1078 = v4 & n1077;
  assign n1079 = n24 & n1062;
  assign n1080 = v7 & n1079;
  assign n1081 = v4 & n1080;
  assign n1082 = ~n1078 & ~n1081;
  assign n1083 = ~n1075 & n1082;
  assign n1084 = ~n1072 & n1083;
  assign n1085 = n30 & n1062;
  assign n1086 = v7 & n1085;
  assign n1087 = v4 & n1086;
  assign n1088 = n998 & n1032;
  assign n1089 = n30 & n1063;
  assign n1090 = n530 & n665;
  assign n1091 = v11 & n1090;
  assign n1092 = n303 & n1091;
  assign n1093 = ~n1089 & ~n1092;
  assign n1094 = ~n1088 & n1093;
  assign n1095 = ~n1087 & n1094;
  assign n1096 = n21 & n981;
  assign n1097 = n82 & n1096;
  assign n1098 = n51 & n981;
  assign n1099 = n75 & n1098;
  assign n1100 = n75 & n1096;
  assign n1101 = n912 & n943;
  assign n1102 = n943 & n1036;
  assign n1103 = n943 & n1038;
  assign n1104 = n75 & n949;
  assign n1105 = n188 & n1104;
  assign n1106 = ~n1103 & ~n1105;
  assign n1107 = ~n1102 & n1106;
  assign n1108 = ~n1101 & n1107;
  assign n1109 = ~n1100 & n1108;
  assign n1110 = ~n1099 & n1109;
  assign n1111 = ~n1097 & n1110;
  assign n1112 = n1095 & n1111;
  assign n1113 = n1084 & n1112;
  assign n1114 = n1071 & n1113;
  assign n1115 = n1055 & n1114;
  assign n1116 = n1042 & n1115;
  assign n1117 = ~v13 & ~v9;
  assign n1118 = ~v10 & n1117;
  assign n1119 = n849 & n1118;
  assign n1120 = n21 & n1119;
  assign n1121 = n24 & n1120;
  assign n1122 = n30 & n1120;
  assign n1123 = n417 & n636;
  assign n1124 = n188 & n1123;
  assign n1125 = ~v3 & n1124;
  assign n1126 = n23 & n1125;
  assign n1127 = n29 & n1125;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1122 & n1128;
  assign n1130 = ~n1121 & n1129;
  assign n1131 = n51 & n1119;
  assign n1132 = n24 & n1131;
  assign n1133 = n30 & n1131;
  assign n1134 = n24 & n1119;
  assign n1135 = ~v5 & n1134;
  assign n1136 = ~v6 & n1135;
  assign n1137 = n30 & n1119;
  assign n1138 = ~v5 & n1137;
  assign n1139 = ~v6 & n1138;
  assign n1140 = ~n1136 & ~n1139;
  assign n1141 = ~n1133 & n1140;
  assign n1142 = ~n1132 & n1141;
  assign n1143 = n77 & n417;
  assign n1144 = n75 & n1143;
  assign n1145 = n188 & n1144;
  assign n1146 = n188 & n1143;
  assign n1147 = ~v2 & n1146;
  assign n1148 = n74 & n1147;
  assign n1149 = n173 & n401;
  assign n1150 = n82 & n1149;
  assign n1151 = ~v5 & n1150;
  assign n1152 = ~v6 & n1151;
  assign n1153 = n280 & n401;
  assign n1154 = n1001 & n1118;
  assign n1155 = n996 & n1118;
  assign n1156 = n373 & n401;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1154 & n1157;
  assign n1159 = ~n1153 & n1158;
  assign n1160 = ~n1152 & n1159;
  assign n1161 = ~n1148 & n1160;
  assign n1162 = ~n1145 & n1161;
  assign n1163 = n173 & n995;
  assign n1164 = n401 & n1163;
  assign n1165 = n401 & n796;
  assign n1166 = n173 & n1000;
  assign n1167 = n401 & n1166;
  assign n1168 = ~n1165 & ~n1167;
  assign n1169 = ~n1164 & n1168;
  assign n1170 = n380 & n401;
  assign n1171 = n417 & n530;
  assign n1172 = n77 & n1171;
  assign n1173 = n234 & n417;
  assign n1174 = n77 & n1173;
  assign n1175 = n229 & n401;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~n1172 & n1176;
  assign n1178 = ~n1170 & n1177;
  assign n1179 = n232 & n401;
  assign n1180 = n241 & n401;
  assign n1181 = n245 & n401;
  assign n1182 = n248 & n401;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n1180 & n1183;
  assign n1185 = ~n1179 & n1184;
  assign n1186 = n251 & n401;
  assign n1187 = n257 & n401;
  assign n1188 = n260 & n401;
  assign n1189 = n264 & n401;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = ~n1187 & n1190;
  assign n1192 = ~n1186 & n1191;
  assign n1193 = n1185 & n1192;
  assign n1194 = n1178 & n1193;
  assign n1195 = n1169 & n1194;
  assign n1196 = n1162 & n1195;
  assign n1197 = n1142 & n1196;
  assign n1198 = n1130 & n1197;
  assign n1199 = ~v10 & ~v9;
  assign n1200 = n665 & n1199;
  assign n1201 = n51 & n1200;
  assign n1202 = n75 & n1201;
  assign n1203 = n82 & n1201;
  assign n1204 = n75 & n1200;
  assign n1205 = ~v5 & n1204;
  assign n1206 = ~v6 & n1205;
  assign n1207 = n82 & n1200;
  assign n1208 = ~v5 & n1207;
  assign n1209 = ~v6 & n1208;
  assign n1210 = ~n1206 & ~n1209;
  assign n1211 = ~n1203 & n1210;
  assign n1212 = ~n1202 & n1211;
  assign n1213 = n417 & n665;
  assign n1214 = n75 & n1213;
  assign n1215 = n188 & n1214;
  assign n1216 = n188 & n1213;
  assign n1217 = ~v2 & n1216;
  assign n1218 = n74 & n1217;
  assign n1219 = n94 & n1200;
  assign n1220 = n75 & n1219;
  assign n1221 = v12 & n169;
  assign n1222 = n850 & n1221;
  assign n1223 = ~n1220 & ~n1222;
  assign n1224 = ~n1218 & n1223;
  assign n1225 = ~n1215 & n1224;
  assign n1226 = n24 & n1201;
  assign n1227 = n30 & n1201;
  assign n1228 = ~v3 & n1216;
  assign n1229 = n29 & n1228;
  assign n1230 = v12 & n1199;
  assign n1231 = n899 & n1230;
  assign n1232 = n901 & n1230;
  assign n1233 = n903 & n1230;
  assign n1234 = n905 & n1230;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1232 & n1235;
  assign n1237 = ~n1231 & n1236;
  assign n1238 = ~n1229 & n1237;
  assign n1239 = ~n1227 & n1238;
  assign n1240 = ~n1226 & n1239;
  assign n1241 = n905 & n1118;
  assign n1242 = n910 & n1118;
  assign n1243 = n903 & n1118;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1241 & n1244;
  assign n1246 = n912 & n1118;
  assign n1247 = n914 & n1118;
  assign n1248 = n916 & n1118;
  assign n1249 = n273 & n417;
  assign n1250 = n636 & n1249;
  assign n1251 = ~n1248 & ~n1250;
  assign n1252 = ~n1247 & n1251;
  assign n1253 = ~n1246 & n1252;
  assign n1254 = n276 & n417;
  assign n1255 = n636 & n1254;
  assign n1256 = n927 & n1118;
  assign n1257 = n1001 & n1230;
  assign n1258 = n996 & n1230;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1256 & n1259;
  assign n1261 = ~n1255 & n1260;
  assign n1262 = n929 & n1118;
  assign n1263 = n998 & n1230;
  assign n1264 = n947 & n1230;
  assign n1265 = ~v10 & n665;
  assign n1266 = ~v7 & n1265;
  assign n1267 = ~v9 & n1266;
  assign n1268 = n24 & n1267;
  assign n1269 = v6 & n1268;
  assign n1270 = n187 & n1269;
  assign n1271 = ~n1264 & ~n1270;
  assign n1272 = ~n1263 & n1271;
  assign n1273 = ~n1262 & n1272;
  assign n1274 = n1261 & n1273;
  assign n1275 = n1253 & n1274;
  assign n1276 = n1245 & n1275;
  assign n1277 = n1240 & n1276;
  assign n1278 = n1225 & n1277;
  assign n1279 = n1212 & n1278;
  assign n1280 = n1198 & n1279;
  assign n1281 = n1116 & n1280;
  assign n1282 = n1031 & n1281;
  assign n1283 = v12 & v8;
  assign n1284 = v11 & n1283;
  assign n1285 = n945 & n1284;
  assign n1286 = n947 & n1284;
  assign n1287 = n531 & n665;
  assign n1288 = ~v15 & n533;
  assign n1289 = n664 & n1288;
  assign n1290 = ~n1287 & ~n1289;
  assign n1291 = ~n1286 & n1290;
  assign n1292 = ~n1285 & n1291;
  assign n1293 = n957 & n1284;
  assign n1294 = n892 & n1284;
  assign n1295 = n961 & n1284;
  assign n1296 = n964 & n1284;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = ~n1294 & n1297;
  assign n1299 = ~n1293 & n1298;
  assign n1300 = n190 & n665;
  assign n1301 = n75 & n1300;
  assign n1302 = n188 & n1301;
  assign n1303 = n188 & n1300;
  assign n1304 = ~v2 & n1303;
  assign n1305 = n74 & n1304;
  assign n1306 = n1038 & n1221;
  assign n1307 = n849 & n1221;
  assign n1308 = n75 & n1307;
  assign n1309 = v7 & n1308;
  assign n1310 = v4 & n1309;
  assign n1311 = n849 & n1284;
  assign n1312 = n24 & n1311;
  assign n1313 = v7 & n1312;
  assign n1314 = v4 & n1313;
  assign n1315 = n30 & n1311;
  assign n1316 = v7 & n1315;
  assign n1317 = v4 & n1316;
  assign n1318 = n82 & n1307;
  assign n1319 = v7 & n1318;
  assign n1320 = v4 & n1319;
  assign n1321 = ~n1317 & ~n1320;
  assign n1322 = ~n1314 & n1321;
  assign n1323 = ~n1310 & n1322;
  assign n1324 = ~n1306 & n1323;
  assign n1325 = ~n1305 & n1324;
  assign n1326 = ~n1302 & n1325;
  assign n1327 = n51 & n1307;
  assign n1328 = n30 & n1327;
  assign n1329 = n899 & n1221;
  assign n1330 = n901 & n1221;
  assign n1331 = n21 & n1307;
  assign n1332 = n75 & n1331;
  assign n1333 = ~n1330 & ~n1332;
  assign n1334 = ~n1329 & n1333;
  assign n1335 = ~n1328 & n1334;
  assign n1336 = n82 & n1331;
  assign n1337 = n75 & n1327;
  assign n1338 = n82 & n1327;
  assign n1339 = n914 & n1221;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = ~n1337 & n1340;
  assign n1342 = ~n1336 & n1341;
  assign n1343 = n929 & n1230;
  assign n1344 = n998 & n1221;
  assign n1345 = n30 & n1307;
  assign n1346 = v7 & n1345;
  assign n1347 = v4 & n1346;
  assign n1348 = n947 & n1221;
  assign n1349 = ~v3 & n1303;
  assign n1350 = n23 & n1349;
  assign n1351 = n29 & n1349;
  assign n1352 = n957 & n1221;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n1350 & n1353;
  assign n1355 = ~n1348 & n1354;
  assign n1356 = ~n1347 & n1355;
  assign n1357 = ~n1344 & n1356;
  assign n1358 = ~n1343 & n1357;
  assign n1359 = n1342 & n1358;
  assign n1360 = n1335 & n1359;
  assign n1361 = n1326 & n1360;
  assign n1362 = n1299 & n1361;
  assign n1363 = n1292 & n1362;
  assign n1364 = v7 & n187;
  assign n1365 = v11 & n37;
  assign n1366 = n1364 & n1365;
  assign n1367 = v10 & v8;
  assign n1368 = ~v11 & n1367;
  assign n1369 = n1364 & n1368;
  assign n1370 = ~v13 & v15;
  assign n1371 = n1364 & n1370;
  assign n1372 = ~v13 & n1364;
  assign n1373 = ~v14 & n1372;
  assign n1374 = ~n1371 & ~n1373;
  assign n1375 = ~n1369 & n1374;
  assign n1376 = ~n1366 & n1375;
  assign n1377 = v10 & ~v9;
  assign n1378 = ~v11 & n1377;
  assign n1379 = n1364 & n1378;
  assign n1380 = ~v10 & n37;
  assign n1381 = n1364 & n1380;
  assign n1382 = v12 & ~v6;
  assign n1383 = ~v14 & n1382;
  assign n1384 = n187 & n1383;
  assign n1385 = ~v6 & n187;
  assign n1386 = ~v12 & n1385;
  assign n1387 = v13 & v14;
  assign n1388 = ~v15 & n1387;
  assign n1389 = n1386 & n1388;
  assign n1390 = ~n1384 & ~n1389;
  assign n1391 = ~n1381 & n1390;
  assign n1392 = ~n1379 & n1391;
  assign n1393 = v2 & n74;
  assign n1394 = ~v14 & n1393;
  assign n1395 = ~v3 & n1394;
  assign n1396 = ~v13 & n1395;
  assign n1397 = ~v3 & n1393;
  assign n1398 = n1378 & n1397;
  assign n1399 = ~v13 & ~v3;
  assign n1400 = v15 & n1399;
  assign n1401 = n1393 & n1400;
  assign n1402 = n1380 & n1397;
  assign n1403 = v12 & v7;
  assign n1404 = ~v14 & n1403;
  assign n1405 = n187 & n1404;
  assign n1406 = ~v12 & n1364;
  assign n1407 = n1388 & n1406;
  assign n1408 = v15 & n1364;
  assign n1409 = v12 & n1408;
  assign n1410 = ~n1407 & ~n1409;
  assign n1411 = ~n1405 & n1410;
  assign n1412 = ~n1402 & n1411;
  assign n1413 = ~n1401 & n1412;
  assign n1414 = ~n1398 & n1413;
  assign n1415 = ~n1396 & n1414;
  assign n1416 = n325 & n665;
  assign n1417 = n276 & n1416;
  assign n1418 = n75 & n1311;
  assign n1419 = v7 & n1418;
  assign n1420 = v4 & n1419;
  assign n1421 = n82 & n1311;
  assign n1422 = v7 & n1421;
  assign n1423 = v4 & n1422;
  assign n1424 = v12 & ~v3;
  assign n1425 = ~v14 & n1424;
  assign n1426 = n1393 & n1425;
  assign n1427 = ~n1423 & ~n1426;
  assign n1428 = ~n1420 & n1427;
  assign n1429 = ~n1417 & n1428;
  assign n1430 = v14 & n19;
  assign n1431 = ~v15 & n1430;
  assign n1432 = n1397 & n1431;
  assign n1433 = v15 & n1424;
  assign n1434 = n1393 & n1433;
  assign n1435 = n1365 & n1397;
  assign n1436 = n1368 & n1397;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1434 & n1437;
  assign n1439 = ~n1432 & n1438;
  assign n1440 = n21 & n1311;
  assign n1441 = n82 & n1440;
  assign n1442 = n51 & n1311;
  assign n1443 = n75 & n1442;
  assign n1444 = n75 & n1440;
  assign n1445 = n912 & n1284;
  assign n1446 = n1036 & n1284;
  assign n1447 = n1038 & n1284;
  assign n1448 = n273 & n325;
  assign n1449 = n665 & n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = ~n1446 & n1450;
  assign n1452 = ~n1445 & n1451;
  assign n1453 = ~n1444 & n1452;
  assign n1454 = ~n1443 & n1453;
  assign n1455 = ~n1441 & n1454;
  assign n1456 = n1439 & n1455;
  assign n1457 = n1429 & n1456;
  assign n1458 = n1415 & n1457;
  assign n1459 = n1392 & n1458;
  assign n1460 = n1376 & n1459;
  assign n1461 = v0 & v3;
  assign n1462 = ~v13 & n1461;
  assign n1463 = ~v14 & n1462;
  assign n1464 = n1378 & n1461;
  assign n1465 = n1380 & n1461;
  assign n1466 = ~v1 & v3;
  assign n1467 = v12 & n1466;
  assign n1468 = ~v14 & n1467;
  assign n1469 = ~n1465 & ~n1468;
  assign n1470 = ~n1464 & n1469;
  assign n1471 = ~n1463 & n1470;
  assign n1472 = ~v12 & n1466;
  assign n1473 = n1388 & n1472;
  assign n1474 = v15 & n1467;
  assign n1475 = v11 & v9;
  assign n1476 = ~v8 & n1466;
  assign n1477 = n1475 & n1476;
  assign n1478 = v8 & n1466;
  assign n1479 = v10 & ~v11;
  assign n1480 = n1478 & n1479;
  assign n1481 = ~n1477 & ~n1480;
  assign n1482 = ~n1474 & n1481;
  assign n1483 = ~n1473 & n1482;
  assign n1484 = v12 & n1461;
  assign n1485 = ~v14 & n1484;
  assign n1486 = ~v12 & n1461;
  assign n1487 = n1388 & n1486;
  assign n1488 = ~v5 & v6;
  assign n1489 = ~v7 & n1488;
  assign n1490 = n1380 & n1489;
  assign n1491 = v15 & n1461;
  assign n1492 = v12 & n1491;
  assign n1493 = ~v8 & n1461;
  assign n1494 = v9 & n1493;
  assign n1495 = v11 & n1494;
  assign n1496 = v8 & n1479;
  assign n1497 = v0 & n1496;
  assign n1498 = v3 & n1497;
  assign n1499 = v15 & n1462;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1495 & n1500;
  assign n1502 = ~n1492 & n1501;
  assign n1503 = ~n1490 & n1502;
  assign n1504 = ~n1487 & n1503;
  assign n1505 = ~n1485 & n1504;
  assign n1506 = v12 & ~v14;
  assign n1507 = n1489 & n1506;
  assign n1508 = ~v12 & n1489;
  assign n1509 = n1388 & n1508;
  assign n1510 = v15 & n1489;
  assign n1511 = v12 & n1510;
  assign n1512 = n1365 & n1489;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = ~n1509 & n1513;
  assign n1515 = ~n1507 & n1514;
  assign n1516 = n1368 & n1489;
  assign n1517 = n1370 & n1489;
  assign n1518 = ~v13 & ~v14;
  assign n1519 = n1489 & n1518;
  assign n1520 = n1378 & n1489;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n1517 & n1521;
  assign n1523 = ~n1516 & n1522;
  assign n1524 = n1365 & n1385;
  assign n1525 = n1368 & n1385;
  assign n1526 = v15 & n1385;
  assign n1527 = v12 & n1526;
  assign n1528 = ~v13 & ~v6;
  assign n1529 = v15 & n1528;
  assign n1530 = n187 & n1529;
  assign n1531 = ~v13 & n1385;
  assign n1532 = ~v14 & n1531;
  assign n1533 = n1378 & n1385;
  assign n1534 = n1380 & n1385;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = ~n1532 & n1535;
  assign n1537 = ~n1530 & n1536;
  assign n1538 = ~n1527 & n1537;
  assign n1539 = ~n1525 & n1538;
  assign n1540 = ~n1524 & n1539;
  assign n1541 = n1523 & n1540;
  assign n1542 = n1515 & n1541;
  assign n1543 = n1505 & n1542;
  assign n1544 = n1483 & n1543;
  assign n1545 = n1471 & n1544;
  assign n1546 = v4 & v6;
  assign n1547 = ~v7 & n1546;
  assign n1548 = n1365 & n1547;
  assign n1549 = n1368 & n1547;
  assign n1550 = ~v13 & ~v7;
  assign n1551 = v15 & n1550;
  assign n1552 = n1546 & n1551;
  assign n1553 = ~v13 & n1547;
  assign n1554 = ~v14 & n1553;
  assign n1555 = ~n1552 & ~n1554;
  assign n1556 = ~n1549 & n1555;
  assign n1557 = ~n1548 & n1556;
  assign n1558 = n1378 & n1547;
  assign n1559 = n1380 & n1547;
  assign n1560 = v0 & ~v2;
  assign n1561 = v12 & n1560;
  assign n1562 = ~v14 & n1561;
  assign n1563 = ~v12 & n1560;
  assign n1564 = n1388 & n1563;
  assign n1565 = ~n1562 & ~n1564;
  assign n1566 = ~n1559 & n1565;
  assign n1567 = ~n1558 & n1566;
  assign n1568 = ~v13 & n1466;
  assign n1569 = ~v14 & n1568;
  assign n1570 = ~v9 & n1466;
  assign n1571 = n1479 & n1570;
  assign n1572 = v15 & n1568;
  assign n1573 = ~v10 & v9;
  assign n1574 = n1476 & n1573;
  assign n1575 = n1506 & n1547;
  assign n1576 = ~v12 & n1547;
  assign n1577 = n1388 & n1576;
  assign n1578 = v15 & n1547;
  assign n1579 = v12 & n1578;
  assign n1580 = ~n1577 & ~n1579;
  assign n1581 = ~n1575 & n1580;
  assign n1582 = ~n1574 & n1581;
  assign n1583 = ~n1572 & n1582;
  assign n1584 = ~n1571 & n1583;
  assign n1585 = ~n1569 & n1584;
  assign n1586 = v15 & n1561;
  assign n1587 = ~v8 & n1560;
  assign n1588 = v9 & n1587;
  assign n1589 = v11 & n1588;
  assign n1590 = v8 & n1560;
  assign n1591 = n1479 & n1590;
  assign n1592 = ~v13 & n1560;
  assign n1593 = v15 & n1592;
  assign n1594 = ~n1591 & ~n1593;
  assign n1595 = ~n1589 & n1594;
  assign n1596 = ~n1586 & n1595;
  assign n1597 = ~v14 & n1592;
  assign n1598 = ~v9 & n1560;
  assign n1599 = n1479 & n1598;
  assign n1600 = n1573 & n1587;
  assign n1601 = ~v1 & ~v2;
  assign n1602 = v12 & n1601;
  assign n1603 = ~v14 & n1602;
  assign n1604 = ~n1600 & ~n1603;
  assign n1605 = ~n1599 & n1604;
  assign n1606 = ~n1597 & n1605;
  assign n1607 = ~v12 & ~v1;
  assign n1608 = ~v2 & n1607;
  assign n1609 = n1388 & n1608;
  assign n1610 = v15 & n1602;
  assign n1611 = ~v1 & ~v8;
  assign n1612 = ~v2 & n1611;
  assign n1613 = v9 & n1612;
  assign n1614 = v11 & n1613;
  assign n1615 = n1368 & n1601;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~n1610 & n1616;
  assign n1618 = ~n1609 & n1617;
  assign n1619 = ~v13 & n1601;
  assign n1620 = v15 & n1619;
  assign n1621 = ~v14 & n1619;
  assign n1622 = ~v1 & ~v9;
  assign n1623 = ~v2 & n1622;
  assign n1624 = n1479 & n1623;
  assign n1625 = n1573 & n1612;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~n1621 & n1626;
  assign n1628 = ~n1620 & n1627;
  assign n1629 = n1618 & n1628;
  assign n1630 = n1606 & n1629;
  assign n1631 = n1596 & n1630;
  assign n1632 = n1585 & n1631;
  assign n1633 = n1567 & n1632;
  assign n1634 = n1557 & n1633;
  assign n1635 = n1545 & n1634;
  assign n1636 = n1460 & n1635;
  assign n1637 = n1363 & n1636;
  assign n1638 = n1282 & n1637;
  assign n1639 = n942 & n1638;
  assign \v16.0  = ~n523 | ~n1639;
endmodule


