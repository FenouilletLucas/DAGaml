// Benchmark "i10" written by ABC on Tue May 16 16:07:49 2017

module i10 ( 
    \V223(1) , \V223(0) , \V100(3) , \V100(2) , \V100(5) , \V100(4) ,
    \V100(1) , \V100(0) , \V60(0) , \V247(0) , \V7(0) , \V124(3) ,
    \V124(2) , \V124(5) , \V124(4) , \V11(0) , \V124(1) , \V124(0) ,
    \V259(0) , \V84(0) , \V84(1) , \V84(2) , \V84(3) , \V84(4) , \V84(5) ,
    \V35(0) , \V302(0) , \V59(0) , \V240(0) , \V203(0) , \V288(3) ,
    \V215(0) , \V288(2) , \V288(5) , \V288(4) , \V40(0) , \V288(1) ,
    \V288(0) , \V165(3) , \V165(2) , \V165(5) , \V165(4) , \V239(3) ,
    \V288(7) , \V239(2) , \V288(6) , \V52(0) , \V165(1) , \V239(4) ,
    \V165(0) , \V239(1) , \V239(0) , \V165(7) , \V165(6) , \V177(0) ,
    \V189(3) , \V189(2) , \V189(5) , \V189(4) , \V189(1) , \V189(0) ,
    \V15(0) , \V88(0) , \V88(1) , \V88(2) , \V88(3) , \V39(0) , \V293(0) ,
    \V244(0) , \V4(0) , \V194(3) , \V194(2) , \V194(4) , \V268(3) ,
    \V268(2) , \V268(5) , \V194(1) , \V268(4) , \V194(0) , \V268(1) ,
    \V268(0) , \V207(0) , \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V32(4) ,
    \V32(5) , \V32(6) , \V32(7) , \V32(8) , \V44(0) , \V32(9) , \V108(3) ,
    \V108(2) , \V56(0) , \V108(5) , \V108(4) , \V169(1) , \V169(0) ,
    \V108(1) , \V108(0) , \V68(0) , \V261(0) , \V101(0) , \V174(0) ,
    \V248(0) , \V8(0) , \V12(0) , \V149(3) , \V149(2) , \V149(5) ,
    \V149(4) , \V149(1) , \V149(0) , \V149(7) , \V149(6) , \V48(0) ,
    \V290(0) , \V32(11) , \V32(10) , \V241(0) , \V1(0) , \V204(0) ,
    \V277(0) , \V216(0) , \V41(0) , \V289(0) , \V53(0) , \V65(0) ,
    \V16(0) , \V270(0) , \V294(0) , \V171(0) , \V183(3) , \V110(0) ,
    \V183(2) , \V245(0) , \V183(5) , \V5(0) , \V183(4) , \V257(3) ,
    \V257(2) , \V70(0) , \V257(5) , \V183(1) , \V257(4) , \V183(0) ,
    \V257(1) , \V257(0) , \V257(7) , \V257(6) , \V134(1) , \V134(0) ,
    \V269(0) , \V94(0) , \V94(1) , \V33(0) , \V45(0) , \V57(0) , \V109(0) ,
    \V69(0) , \V262(0) , \V213(3) , \V213(2) , \V213(5) , \V213(4) ,
    \V274(0) , \V213(1) , \V213(0) , \V50(0) , \V102(0) , \V62(0) ,
    \V175(0) , \V249(0) , \V9(0) , \V13(0) , \V199(3) , \V199(2) ,
    \V199(4) , \V199(1) , \V199(0) , \V37(0) , \V291(0) , \V242(0) ,
    \V2(0) , \V205(0) , \V91(0) , \V91(1) , \V278(0) , \V229(3) ,
    \V229(2) , \V42(0) , \V229(5) , \V229(4) , \V229(1) , \V229(0) ,
    \V118(3) , \V118(2) , \V66(0) , \V118(5) , \V118(4) , \V118(1) ,
    \V118(0) , \V78(0) , \V78(1) , \V118(7) , \V78(2) , \V118(6) ,
    \V78(3) , \V78(4) , \V78(5) , \V271(0) , \V234(3) , \V234(2) ,
    \V234(4) , \V295(0) , \V234(1) , \V234(0) , \V172(0) , \V246(0) ,
    \V6(0) , \V71(0) , \V10(0) , \V258(0) , \V34(0) , \V46(0) , \V301(0) ,
    \V202(0) , \V275(0) , \V214(0) , \V51(0) , \V63(0) , \V14(0) ,
    \V38(0) , \V280(0) , \V292(0) , \V243(0) , \V3(0) , \V132(3) ,
    \V132(2) , \V132(5) , \V132(4) , \V132(1) , \V132(0) , \V132(7) ,
    \V132(6) , \V279(0) , \V43(0) , \V55(0) , \V67(0) , \V260(0) ,
    \V272(0) , \V223(3) , \V223(2) , \V223(5) , \V223(4) ,
    \V1243(7) , \V500(0) , \V1243(6) , \V1243(9) , \V1243(8) , \V1243(1) ,
    \V1243(0) , \V1717(0) , \V1243(3) , \V1243(2) , \V1243(5) , \V1243(4) ,
    \V585(0) , \V597(0) , \V1679(0) , \V1833(0) , \V1968(0) , \V1771(1) ,
    \V1771(0) , \V640(0) , \V375(0) , \V603(0) , \V1758(0) , \V1900(0) ,
    \V1709(1) , \V1709(0) , \V1709(3) , \V1709(2) , \V1709(4) , \V1512(1) ,
    \V1512(3) , \V1512(2) , \V1536(0) , \V1898(0) , \V1652(0) , \V1726(0) ,
    \V1953(7) , \V1953(6) , \V410(0) , \V1953(1) , \V1953(0) , \V1953(3) ,
    \V1953(2) , \V1953(5) , \V1953(4) , \V508(0) , \V1392(0) , \V1829(7) ,
    \V1829(6) , \V1829(9) , \V1829(8) , \V1281(0) , \V1620(0) , \V1829(1) ,
    \V1829(0) , \V1829(3) , \V1829(2) , \V1693(0) , \V1829(5) , \V1829(4) ,
    \V1921(1) , \V1921(0) , \V1921(3) , \V1921(2) , \V1921(5) , \V1921(4) ,
    \V802(0) , \V826(0) , \V1213(10) , \V1213(11) , \V1760(0) , \V1495(0) ,
    \V591(0) , \V1759(0) , \V1901(0) , \V1297(1) , \V1297(0) , \V1297(3) ,
    \V1297(2) , \V1297(4) , \V1451(0) , \V1863(0) , \V393(0) , \V1899(0) ,
    \V1480(0) , \V423(0) , \V1492(0) , \V435(0) , \V1781(1) , \V1781(0) ,
    V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265,
    V1266, V1267, \V1467(0) , V1365, V1370, V1371, V1372, V1373, V1374,
    V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1423, V1426, V1428,
    V1429, V1431, V1432, V1470, \V1645(0) , V1537, V1539, V1669, V1719,
    \V1896(0) , V1736, V1832, \V1459(0) , \V1213(7) , \V1213(6) ,
    \V1213(9) , \V1213(8) , \V1613(1) , \V1274(0) , \V1613(0) , \V1213(1) ,
    \V1213(0) , \V1213(3) , \V1213(2) , \V1213(5) , \V1213(4) , \V1440(0) ,
    \V321(2) , \V1864(0) , \V1741(0) , \V572(3) , \V572(2) , \V634(0) ,
    \V572(5) , \V572(4) , \V1439(0) , \V572(1) , \V572(0) , \V511(0) ,
    \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) , \V1992(0) ,
    \V609(0) , \V1481(0) , \V1629(0) , \V798(0) , \V398(0) , \V1671(0) ,
    \V1745(0) , \V1757(0) , \V1960(1) , \V1960(0) , V356, V357, V373, V377,
    \V1897(0) , V432, V512, V527, V537, V538, V539, V540, V541, V542, V543,
    V544, V545, V546, V547, V548, V587, V620, V621, V630, V650, V651, V652,
    V653, V654, V655, V656, V657, \V821(0) , \V1552(1) , \V1552(0) , V707,
    V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V801,
    V966, V986  );
  input  \V223(1) , \V223(0) , \V100(3) , \V100(2) , \V100(5) ,
    \V100(4) , \V100(1) , \V100(0) , \V60(0) , \V247(0) , \V7(0) ,
    \V124(3) , \V124(2) , \V124(5) , \V124(4) , \V11(0) , \V124(1) ,
    \V124(0) , \V259(0) , \V84(0) , \V84(1) , \V84(2) , \V84(3) , \V84(4) ,
    \V84(5) , \V35(0) , \V302(0) , \V59(0) , \V240(0) , \V203(0) ,
    \V288(3) , \V215(0) , \V288(2) , \V288(5) , \V288(4) , \V40(0) ,
    \V288(1) , \V288(0) , \V165(3) , \V165(2) , \V165(5) , \V165(4) ,
    \V239(3) , \V288(7) , \V239(2) , \V288(6) , \V52(0) , \V165(1) ,
    \V239(4) , \V165(0) , \V239(1) , \V239(0) , \V165(7) , \V165(6) ,
    \V177(0) , \V189(3) , \V189(2) , \V189(5) , \V189(4) , \V189(1) ,
    \V189(0) , \V15(0) , \V88(0) , \V88(1) , \V88(2) , \V88(3) , \V39(0) ,
    \V293(0) , \V244(0) , \V4(0) , \V194(3) , \V194(2) , \V194(4) ,
    \V268(3) , \V268(2) , \V268(5) , \V194(1) , \V268(4) , \V194(0) ,
    \V268(1) , \V268(0) , \V207(0) , \V32(0) , \V32(1) , \V32(2) ,
    \V32(3) , \V32(4) , \V32(5) , \V32(6) , \V32(7) , \V32(8) , \V44(0) ,
    \V32(9) , \V108(3) , \V108(2) , \V56(0) , \V108(5) , \V108(4) ,
    \V169(1) , \V169(0) , \V108(1) , \V108(0) , \V68(0) , \V261(0) ,
    \V101(0) , \V174(0) , \V248(0) , \V8(0) , \V12(0) , \V149(3) ,
    \V149(2) , \V149(5) , \V149(4) , \V149(1) , \V149(0) , \V149(7) ,
    \V149(6) , \V48(0) , \V290(0) , \V32(11) , \V32(10) , \V241(0) ,
    \V1(0) , \V204(0) , \V277(0) , \V216(0) , \V41(0) , \V289(0) ,
    \V53(0) , \V65(0) , \V16(0) , \V270(0) , \V294(0) , \V171(0) ,
    \V183(3) , \V110(0) , \V183(2) , \V245(0) , \V183(5) , \V5(0) ,
    \V183(4) , \V257(3) , \V257(2) , \V70(0) , \V257(5) , \V183(1) ,
    \V257(4) , \V183(0) , \V257(1) , \V257(0) , \V257(7) , \V257(6) ,
    \V134(1) , \V134(0) , \V269(0) , \V94(0) , \V94(1) , \V33(0) ,
    \V45(0) , \V57(0) , \V109(0) , \V69(0) , \V262(0) , \V213(3) ,
    \V213(2) , \V213(5) , \V213(4) , \V274(0) , \V213(1) , \V213(0) ,
    \V50(0) , \V102(0) , \V62(0) , \V175(0) , \V249(0) , \V9(0) , \V13(0) ,
    \V199(3) , \V199(2) , \V199(4) , \V199(1) , \V199(0) , \V37(0) ,
    \V291(0) , \V242(0) , \V2(0) , \V205(0) , \V91(0) , \V91(1) ,
    \V278(0) , \V229(3) , \V229(2) , \V42(0) , \V229(5) , \V229(4) ,
    \V229(1) , \V229(0) , \V118(3) , \V118(2) , \V66(0) , \V118(5) ,
    \V118(4) , \V118(1) , \V118(0) , \V78(0) , \V78(1) , \V118(7) ,
    \V78(2) , \V118(6) , \V78(3) , \V78(4) , \V78(5) , \V271(0) ,
    \V234(3) , \V234(2) , \V234(4) , \V295(0) , \V234(1) , \V234(0) ,
    \V172(0) , \V246(0) , \V6(0) , \V71(0) , \V10(0) , \V258(0) , \V34(0) ,
    \V46(0) , \V301(0) , \V202(0) , \V275(0) , \V214(0) , \V51(0) ,
    \V63(0) , \V14(0) , \V38(0) , \V280(0) , \V292(0) , \V243(0) , \V3(0) ,
    \V132(3) , \V132(2) , \V132(5) , \V132(4) , \V132(1) , \V132(0) ,
    \V132(7) , \V132(6) , \V279(0) , \V43(0) , \V55(0) , \V67(0) ,
    \V260(0) , \V272(0) , \V223(3) , \V223(2) , \V223(5) , \V223(4) ;
  output \V1243(7) , \V500(0) , \V1243(6) , \V1243(9) , \V1243(8) ,
    \V1243(1) , \V1243(0) , \V1717(0) , \V1243(3) , \V1243(2) , \V1243(5) ,
    \V1243(4) , \V585(0) , \V597(0) , \V1679(0) , \V1833(0) , \V1968(0) ,
    \V1771(1) , \V1771(0) , \V640(0) , \V375(0) , \V603(0) , \V1758(0) ,
    \V1900(0) , \V1709(1) , \V1709(0) , \V1709(3) , \V1709(2) , \V1709(4) ,
    \V1512(1) , \V1512(3) , \V1512(2) , \V1536(0) , \V1898(0) , \V1652(0) ,
    \V1726(0) , \V1953(7) , \V1953(6) , \V410(0) , \V1953(1) , \V1953(0) ,
    \V1953(3) , \V1953(2) , \V1953(5) , \V1953(4) , \V508(0) , \V1392(0) ,
    \V1829(7) , \V1829(6) , \V1829(9) , \V1829(8) , \V1281(0) , \V1620(0) ,
    \V1829(1) , \V1829(0) , \V1829(3) , \V1829(2) , \V1693(0) , \V1829(5) ,
    \V1829(4) , \V1921(1) , \V1921(0) , \V1921(3) , \V1921(2) , \V1921(5) ,
    \V1921(4) , \V802(0) , \V826(0) , \V1213(10) , \V1213(11) , \V1760(0) ,
    \V1495(0) , \V591(0) , \V1759(0) , \V1901(0) , \V1297(1) , \V1297(0) ,
    \V1297(3) , \V1297(2) , \V1297(4) , \V1451(0) , \V1863(0) , \V393(0) ,
    \V1899(0) , \V1480(0) , \V423(0) , \V1492(0) , \V435(0) , \V1781(1) ,
    \V1781(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1467(0) , V1365, V1370, V1371, V1372,
    V1373, V1374, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1423,
    V1426, V1428, V1429, V1431, V1432, V1470, \V1645(0) , V1537, V1539,
    V1669, V1719, \V1896(0) , V1736, V1832, \V1459(0) , \V1213(7) ,
    \V1213(6) , \V1213(9) , \V1213(8) , \V1613(1) , \V1274(0) , \V1613(0) ,
    \V1213(1) , \V1213(0) , \V1213(3) , \V1213(2) , \V1213(5) , \V1213(4) ,
    \V1440(0) , \V321(2) , \V1864(0) , \V1741(0) , \V572(3) , \V572(2) ,
    \V634(0) , \V572(5) , \V572(4) , \V1439(0) , \V572(1) , \V572(0) ,
    \V511(0) , \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) ,
    \V1992(0) , \V609(0) , \V1481(0) , \V1629(0) , \V798(0) , \V398(0) ,
    \V1671(0) , \V1745(0) , \V1757(0) , \V1960(1) , \V1960(0) , V356, V357,
    V373, V377, \V1897(0) , V432, V512, V527, V537, V538, V539, V540, V541,
    V542, V543, V544, V545, V546, V547, V548, V587, V620, V621, V630, V650,
    V651, V652, V653, V654, V655, V656, V657, \V821(0) , \V1552(1) ,
    \V1552(0) , V707, V763, V775, V778, V779, V780, V781, V782, V783, V784,
    V787, V789, V801, V966, V986;
  wire n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n947, n948, n949, n950, n951,
    n952, n954, n955, n956, n957, n958, n960, n961, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n974, n975, n976, n977, n979, n980,
    n981, n982, n984, n985, n989, n997, n998, n999, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1011, n1012, n1013, n1014,
    n1015, n1017, n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1040, n1041, n1042, n1043, n1044, n1046, n1047, n1048,
    n1049, n1050, n1052, n1053, n1054, n1055, n1056, n1058, n1059, n1060,
    n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1532, n1533, n1534, n1535, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1706, n1707, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1741, n1742, n1743,
    n1744, n1745, n1746, n1748, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1759, n1760, n1762, n1763, n1764, n1765, n1766, n1767,
    n1769, n1770, n1771, n1772, n1773, n1774, n1776, n1777, n1778, n1779,
    n1780, n1781, n1783, n1784, n1785, n1786, n1787, n1788, n1790, n1791,
    n1792, n1793, n1794, n1795, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1910, n1911, n1912, n1913, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1940, n1941, n1942, n1943, n1945, n1946, n1947, n1948,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1976, n1977, n1978, n1979, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2012,
    n2013, n2014, n2015, n2016, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2034,
    n2035, n2036, n2037, n2039, n2040, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2064, n2065, n2066, n2067,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2091, n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2132,
    n2133, n2134, n2135, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2162, n2163, n2164,
    n2165, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2284, n2285, n2286, n2287, n2289, n2290, n2291, n2292, n2293,
    n2294, n2296, n2298, n2299, n2300, n2301, n2302, n2304, n2305, n2306,
    n2307, n2308, n2310, n2311, n2312, n2313, n2314, n2316, n2317, n2318,
    n2319, n2320, n2322, n2323, n2324, n2325, n2326, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2342, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2395, n2396, n2398, n2399, n2400, n2401, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2503, n2504, n2505, n2506, n2508, n2509, n2510, n2511,
    n2513, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2555, n2556, n2558, n2559, n2560, n2561, n2563, n2564, n2565,
    n2567, n2568, n2569, n2571, n2572, n2574, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2598, n2599, n2600, n2602,
    n2603, n2604, n2605, n2607, n2612, n2614, n2615, n2617, n2618, n2620,
    n2622, n2623, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2666, n2667, n2668, n2669, n2671, n2672, n2674, n2675,
    n2677, n2678, n2679, n2680, n2682, n2683, n2684, n2685, n2686, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2705, n2706, n2707, n2708, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2831, n2832, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2870, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2934, n2935, n2936, n2937, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2998, n2999, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3019, n3021, n3022, n3024, n3025, n3026, n3027, n3028, n3029,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3080, n3081, n3082, n3083, n3084, n3086, n3087, n3088,
    n3089, n3091, n3092, n3093, n3094, n3096, n3097, n3098, n3100, n3101,
    n3102, n3104, n3105, n3107, n3109, n3110, n3111, n3112, n3113, n3114,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3125, n3126,
    n3127, n3130, n3131, n3132, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157;
  assign n482 = \V149(3)  & \V149(2) ;
  assign n483 = \V149(1)  & n482;
  assign n484 = ~\V149(0)  & n483;
  assign n485 = ~\V149(4)  & ~\V149(0) ;
  assign n486 = \V149(1)  & n485;
  assign n487 = \V149(2)  & n486;
  assign n488 = ~\V149(3)  & n487;
  assign n489 = \V165(7)  & \V165(6) ;
  assign n490 = \V165(5)  & n489;
  assign n491 = \V165(3)  & n490;
  assign n492 = \V165(4)  & n491;
  assign n493 = \V261(0)  & n492;
  assign n494 = ~\V204(0)  & n493;
  assign n495 = \V165(0)  & n494;
  assign n496 = \V165(1)  & n495;
  assign n497 = \V165(2)  & n496;
  assign n498 = ~\V165(5)  & \V70(0) ;
  assign n499 = \V165(3)  & n498;
  assign n500 = ~\V165(4)  & n499;
  assign n501 = ~\V165(6)  & n500;
  assign \V802(0)  = \V52(0)  | \V51(0) ;
  assign n503 = ~\V149(2)  & \V149(1) ;
  assign n504 = ~\V149(0)  & n503;
  assign n505 = \V149(5)  & ~\V149(7) ;
  assign n506 = ~\V149(3)  & n505;
  assign n507 = n504 & n506;
  assign n508 = \V149(4)  & n507;
  assign n509 = \V149(6)  & n508;
  assign n510 = \V149(5)  & \V149(7) ;
  assign n511 = ~\V149(3)  & n510;
  assign n512 = n504 & n511;
  assign n513 = \V149(4)  & n512;
  assign n514 = \V149(6)  & n513;
  assign n515 = ~n509 & ~n514;
  assign n516 = ~\V55(0)  & ~n515;
  assign n517 = ~\V802(0)  & n516;
  assign n518 = ~\V149(2)  & ~\V149(0) ;
  assign n519 = ~\V149(1)  & n518;
  assign n520 = \V149(4)  & ~\V149(0) ;
  assign n521 = \V149(1)  & n520;
  assign n522 = \V149(2)  & n521;
  assign n523 = ~\V149(3)  & n522;
  assign n524 = ~n519 & ~n523;
  assign n525 = ~n517 & n524;
  assign n526 = \V169(0)  & ~n525;
  assign n527 = ~\V291(0)  & n526;
  assign n528 = ~n501 & n527;
  assign V763 = ~\V292(0)  & n528;
  assign n530 = \V165(7)  & \V70(0) ;
  assign n531 = \V261(0)  & n530;
  assign n532 = \V165(5)  & n531;
  assign n533 = \V165(3)  & n532;
  assign n534 = \V165(4)  & n533;
  assign n535 = \V165(6)  & n534;
  assign n536 = \V165(0)  & n535;
  assign n537 = \V165(1)  & n536;
  assign n538 = \V165(2)  & n537;
  assign n539 = V763 & n538;
  assign n540 = ~n497 & ~n539;
  assign n541 = ~\V262(0)  & n540;
  assign n542 = ~n488 & n541;
  assign n543 = ~n484 & n542;
  assign n544 = \V53(0)  & n543;
  assign n545 = ~\V56(0)  & n544;
  assign n546 = ~\V56(0)  & ~\V53(0) ;
  assign n547 = ~\V57(0)  & n546;
  assign n548 = \V149(2)  & ~\V149(1) ;
  assign n549 = ~\V149(0)  & n548;
  assign n550 = \V149(3)  & n549;
  assign n551 = ~\V174(0)  & n519;
  assign n552 = ~\V149(3)  & ~\V149(4) ;
  assign n553 = n551 & n552;
  assign n554 = \V149(5)  & n553;
  assign n555 = ~\V88(2)  & n554;
  assign n556 = \V88(3)  & n555;
  assign V707 = ~\V149(3)  & n551;
  assign n558 = ~\V149(5)  & ~\V149(4) ;
  assign n559 = V707 & n558;
  assign n560 = \V88(2)  & n559;
  assign n561 = \V88(3)  & n560;
  assign n562 = ~\V88(2)  & n559;
  assign n563 = \V88(3)  & n562;
  assign n564 = ~\V149(5)  & V707;
  assign n565 = \V149(4)  & n564;
  assign n566 = \V149(5)  & V707;
  assign n567 = \V149(4)  & n566;
  assign n568 = ~\V88(3)  & n560;
  assign n569 = ~\V88(3)  & n555;
  assign n570 = \V88(2)  & n554;
  assign n571 = ~\V88(3)  & n570;
  assign n572 = ~n569 & ~n571;
  assign n573 = ~n568 & n572;
  assign n574 = ~n567 & n573;
  assign n575 = ~n565 & n574;
  assign n576 = ~n563 & n575;
  assign n577 = ~n561 & n576;
  assign n578 = ~n556 & n577;
  assign n579 = \V149(3)  & n551;
  assign n580 = ~\V149(3)  & \V149(5) ;
  assign n581 = n549 & n580;
  assign n582 = ~\V149(4)  & n581;
  assign n583 = ~\V149(3)  & ~\V149(5) ;
  assign n584 = n549 & n583;
  assign n585 = ~\V149(4)  & n584;
  assign n586 = \V149(4)  & n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n582 & n587;
  assign n589 = ~\V174(0)  & n523;
  assign n590 = \V277(0)  & n589;
  assign n591 = \V278(0)  & ~n590;
  assign n592 = n589 & ~n591;
  assign n593 = n588 & ~n592;
  assign n594 = ~n579 & n593;
  assign n595 = n578 & n594;
  assign n596 = ~n550 & n595;
  assign n597 = ~n519 & ~n549;
  assign n598 = \V169(1)  & ~n597;
  assign n599 = ~n578 & n598;
  assign n600 = \V56(0)  & n599;
  assign n601 = n579 & n598;
  assign n602 = \V56(0)  & n601;
  assign n603 = \V60(0)  & n601;
  assign n604 = \V60(0)  & n599;
  assign n605 = ~n603 & ~n604;
  assign n606 = ~n602 & n605;
  assign n607 = ~n600 & n606;
  assign n608 = ~n596 & n607;
  assign n609 = ~n547 & n608;
  assign n610 = ~\V149(5)  & \V149(7) ;
  assign n611 = ~\V149(3)  & n610;
  assign n612 = n504 & n611;
  assign n613 = \V149(4)  & n612;
  assign n614 = \V149(6)  & n613;
  assign n615 = ~n609 & ~n614;
  assign n616 = ~n545 & n615;
  assign n617 = ~n550 & ~n589;
  assign n618 = \V60(0)  & ~n617;
  assign n619 = ~n616 & ~n618;
  assign n620 = \V84(5)  & n619;
  assign n621 = ~n616 & n620;
  assign n622 = V763 & n541;
  assign n623 = ~\V59(0)  & ~\V56(0) ;
  assign n624 = ~\V60(0)  & n623;
  assign n625 = V763 & ~n624;
  assign n626 = \V32(9)  & n625;
  assign n627 = n622 & n626;
  assign n628 = n622 & n627;
  assign n629 = n484 & ~n591;
  assign n630 = ~\V59(0)  & n629;
  assign n631 = ~n484 & ~n589;
  assign n632 = ~n488 & n631;
  assign n633 = \V199(2)  & n597;
  assign n634 = ~n632 & n633;
  assign n635 = \V239(2)  & ~n597;
  assign n636 = n632 & n635;
  assign n637 = ~n634 & ~n636;
  assign n638 = ~\V60(0)  & ~\V59(0) ;
  assign n639 = n629 & ~n638;
  assign n640 = n484 & n591;
  assign n641 = ~n589 & n597;
  assign n642 = ~n488 & n641;
  assign n643 = ~\V174(0)  & ~n642;
  assign n644 = ~n640 & ~n643;
  assign n645 = ~n639 & n644;
  assign n646 = ~n637 & ~n645;
  assign n647 = n541 & n646;
  assign n648 = ~n630 & n647;
  assign n649 = ~n622 & n648;
  assign n650 = ~n622 & n649;
  assign n651 = ~n628 & ~n650;
  assign n652 = ~n619 & ~n651;
  assign n653 = n616 & n652;
  assign \V1243(7)  = n621 | n653;
  assign \V500(0)  = \V271(0)  | ~\V14(0) ;
  assign n656 = \V84(4)  & n619;
  assign n657 = ~n616 & n656;
  assign n658 = \V32(11)  & ~n625;
  assign n659 = ~n625 & n658;
  assign n660 = \V32(8)  & n625;
  assign n661 = ~n659 & ~n660;
  assign n662 = n622 & ~n661;
  assign n663 = n622 & n662;
  assign n664 = \V199(1)  & n597;
  assign n665 = ~n632 & n664;
  assign n666 = \V239(1)  & ~n597;
  assign n667 = n632 & n666;
  assign n668 = ~n665 & ~n667;
  assign n669 = ~n645 & ~n668;
  assign n670 = n541 & n669;
  assign n671 = ~n630 & n670;
  assign n672 = ~n622 & n671;
  assign n673 = ~n622 & n672;
  assign n674 = ~n663 & ~n673;
  assign n675 = ~n619 & ~n674;
  assign n676 = n616 & n675;
  assign \V1243(6)  = n657 | n676;
  assign n678 = \V88(1)  & n619;
  assign n679 = ~n616 & n678;
  assign n680 = \V32(11)  & n625;
  assign n681 = n622 & n680;
  assign n682 = n622 & n681;
  assign n683 = \V199(4)  & n597;
  assign n684 = ~n632 & n683;
  assign n685 = \V239(4)  & ~n597;
  assign n686 = n632 & n685;
  assign n687 = ~n684 & ~n686;
  assign n688 = ~n645 & ~n687;
  assign n689 = n541 & n688;
  assign n690 = ~n630 & n689;
  assign n691 = ~n622 & n690;
  assign n692 = ~n622 & n691;
  assign n693 = ~n682 & ~n692;
  assign n694 = ~n619 & ~n693;
  assign n695 = n616 & n694;
  assign \V1243(9)  = n679 | n695;
  assign n697 = \V88(0)  & n619;
  assign n698 = ~n616 & n697;
  assign n699 = \V32(10)  & n625;
  assign n700 = n622 & n699;
  assign n701 = n622 & n700;
  assign n702 = \V199(3)  & n597;
  assign n703 = ~n632 & n702;
  assign n704 = \V239(3)  & ~n597;
  assign n705 = n632 & n704;
  assign n706 = ~n703 & ~n705;
  assign n707 = ~n645 & ~n706;
  assign n708 = n541 & n707;
  assign n709 = ~n630 & n708;
  assign n710 = ~n622 & n709;
  assign n711 = ~n622 & n710;
  assign n712 = ~n701 & ~n711;
  assign n713 = ~n619 & ~n712;
  assign n714 = n616 & n713;
  assign \V1243(8)  = n698 | n714;
  assign n716 = \V78(5)  & n619;
  assign n717 = ~n616 & n716;
  assign n718 = \V32(6)  & ~n625;
  assign n719 = ~n625 & n718;
  assign n720 = \V32(3)  & n625;
  assign n721 = ~n719 & ~n720;
  assign n722 = n622 & ~n721;
  assign n723 = n622 & n722;
  assign n724 = ~\V59(0)  & \V149(5) ;
  assign n725 = ~n591 & n724;
  assign n726 = n484 & n725;
  assign n727 = n541 & n726;
  assign n728 = n645 & n727;
  assign n729 = \V194(1)  & n597;
  assign n730 = ~n632 & n729;
  assign n731 = \V234(1)  & ~n597;
  assign n732 = n632 & n731;
  assign n733 = ~n730 & ~n732;
  assign n734 = n541 & ~n733;
  assign n735 = ~n630 & n734;
  assign n736 = ~n645 & n735;
  assign n737 = ~n728 & ~n736;
  assign n738 = ~n622 & ~n737;
  assign n739 = ~n622 & n738;
  assign n740 = ~n723 & ~n739;
  assign n741 = ~n619 & ~n740;
  assign n742 = n616 & n741;
  assign \V1243(1)  = n717 | n742;
  assign n744 = \V78(4)  & n619;
  assign n745 = ~n616 & n744;
  assign n746 = \V32(5)  & ~n625;
  assign n747 = ~n625 & n746;
  assign n748 = \V32(2)  & n625;
  assign n749 = ~n747 & ~n748;
  assign n750 = n622 & ~n749;
  assign n751 = n622 & n750;
  assign n752 = \V194(0)  & n597;
  assign n753 = ~n632 & n752;
  assign n754 = \V234(0)  & ~n597;
  assign n755 = n632 & n754;
  assign n756 = ~n753 & ~n755;
  assign n757 = n541 & ~n756;
  assign n758 = ~n630 & n757;
  assign n759 = ~n645 & n758;
  assign n760 = ~\V59(0)  & \V149(4) ;
  assign n761 = ~n591 & n760;
  assign n762 = n484 & n761;
  assign n763 = n541 & n762;
  assign n764 = n645 & n763;
  assign n765 = \V257(7)  & ~n541;
  assign n766 = ~n630 & n765;
  assign n767 = n645 & n766;
  assign n768 = ~n764 & ~n767;
  assign n769 = ~n759 & n768;
  assign n770 = ~n622 & ~n769;
  assign n771 = ~n622 & n770;
  assign n772 = ~n751 & ~n771;
  assign n773 = ~n619 & ~n772;
  assign n774 = n616 & n773;
  assign \V321(2)  = ~n745 & ~n774;
  assign n776 = ~n591 & ~n632;
  assign n777 = ~n550 & ~n776;
  assign n778 = \V802(0)  & ~n777;
  assign n779 = ~\V280(0)  & n550;
  assign n780 = \V134(1)  & \V134(0) ;
  assign n781 = \V242(0)  & n780;
  assign n782 = ~\V802(0)  & n781;
  assign n783 = \V272(0)  & n782;
  assign n784 = ~\V275(0)  & n783;
  assign n785 = n591 & n784;
  assign n786 = \V241(0)  & ~n631;
  assign n787 = ~n488 & ~n786;
  assign n788 = \V261(0)  & ~n591;
  assign n789 = ~n787 & n788;
  assign n790 = ~\V802(0)  & n789;
  assign n791 = \V56(0)  & ~n631;
  assign n792 = ~n591 & ~n791;
  assign n793 = \V242(0)  & n792;
  assign n794 = ~\V802(0)  & n793;
  assign n795 = ~n632 & n794;
  assign n796 = ~\V174(0)  & n514;
  assign n797 = \V56(0)  & \V172(0) ;
  assign n798 = \V207(0)  & ~n797;
  assign n799 = \V59(0)  & ~n549;
  assign n800 = n798 & n799;
  assign n801 = n796 & n800;
  assign n802 = ~\V149(4)  & n507;
  assign n803 = ~\V149(6)  & n802;
  assign n804 = ~n549 & n798;
  assign n805 = ~n796 & n804;
  assign n806 = ~n803 & n805;
  assign n807 = ~n598 & n806;
  assign n808 = \V172(0)  & \V67(0) ;
  assign n809 = \V215(0)  & n808;
  assign n810 = ~n549 & n598;
  assign n811 = n798 & n810;
  assign n812 = \V59(0)  & n811;
  assign n813 = ~n549 & n803;
  assign n814 = n798 & n813;
  assign n815 = \V62(0)  & n814;
  assign n816 = ~n812 & ~n815;
  assign n817 = ~\V214(0)  & n816;
  assign n818 = ~n809 & n817;
  assign n819 = ~n807 & n818;
  assign n820 = ~n801 & n819;
  assign n821 = \V261(0)  & ~n787;
  assign n822 = ~\V802(0)  & n821;
  assign n823 = \V272(0)  & n822;
  assign n824 = ~\V275(0)  & n823;
  assign n825 = n591 & n824;
  assign n826 = n820 & ~n825;
  assign n827 = ~n795 & n826;
  assign n828 = ~n790 & n827;
  assign n829 = ~n785 & n828;
  assign n830 = ~\V165(2)  & \V165(0) ;
  assign n831 = \V165(1)  & n830;
  assign n832 = ~\V165(7)  & n831;
  assign n833 = ~\V290(0)  & n831;
  assign n834 = \V165(7)  & n833;
  assign n835 = ~\V302(0)  & ~n834;
  assign n836 = ~n832 & n835;
  assign n837 = n829 & n836;
  assign n838 = \V203(0)  & \V165(1) ;
  assign n839 = ~\V165(0)  & n838;
  assign n840 = \V165(2)  & n839;
  assign n841 = ~n831 & ~n840;
  assign n842 = n837 & n841;
  assign n843 = ~n779 & n842;
  assign n844 = \V240(0)  & n843;
  assign n845 = ~\V172(0)  & n844;
  assign \V1717(0)  = n778 | n845;
  assign n847 = \V84(1)  & n619;
  assign n848 = ~n616 & n847;
  assign n849 = \V32(8)  & ~n625;
  assign n850 = ~n625 & n849;
  assign n851 = \V32(5)  & n625;
  assign n852 = ~n850 & ~n851;
  assign n853 = n622 & ~n852;
  assign n854 = n622 & n853;
  assign n855 = ~\V59(0)  & \V149(7) ;
  assign n856 = ~n591 & n855;
  assign n857 = n484 & n856;
  assign n858 = n541 & n857;
  assign n859 = n645 & n858;
  assign n860 = \V194(3)  & n597;
  assign n861 = ~n632 & n860;
  assign n862 = \V234(3)  & ~n597;
  assign n863 = n632 & n862;
  assign n864 = ~n861 & ~n863;
  assign n865 = n541 & ~n864;
  assign n866 = ~n630 & n865;
  assign n867 = ~n645 & n866;
  assign n868 = ~n859 & ~n867;
  assign n869 = ~n622 & ~n868;
  assign n870 = ~n622 & n869;
  assign n871 = ~n854 & ~n870;
  assign n872 = ~n619 & ~n871;
  assign n873 = n616 & n872;
  assign \V1243(3)  = n848 | n873;
  assign n875 = \V84(0)  & n619;
  assign n876 = ~n616 & n875;
  assign n877 = \V32(7)  & ~n625;
  assign n878 = ~n625 & n877;
  assign n879 = \V32(4)  & n625;
  assign n880 = ~n878 & ~n879;
  assign n881 = n622 & ~n880;
  assign n882 = n622 & n881;
  assign n883 = ~\V59(0)  & \V149(6) ;
  assign n884 = ~n591 & n883;
  assign n885 = n484 & n884;
  assign n886 = n541 & n885;
  assign n887 = n645 & n886;
  assign n888 = \V194(2)  & n597;
  assign n889 = ~n632 & n888;
  assign n890 = \V234(2)  & ~n597;
  assign n891 = n632 & n890;
  assign n892 = ~n889 & ~n891;
  assign n893 = n541 & ~n892;
  assign n894 = ~n630 & n893;
  assign n895 = ~n645 & n894;
  assign n896 = ~n887 & ~n895;
  assign n897 = ~n622 & ~n896;
  assign n898 = ~n622 & n897;
  assign n899 = ~n882 & ~n898;
  assign n900 = ~n619 & ~n899;
  assign n901 = n616 & n900;
  assign \V1243(2)  = n876 | n901;
  assign n903 = \V84(3)  & n619;
  assign n904 = ~n616 & n903;
  assign n905 = \V32(10)  & ~n625;
  assign n906 = ~n625 & n905;
  assign n907 = \V32(7)  & n625;
  assign n908 = ~n906 & ~n907;
  assign n909 = n622 & ~n908;
  assign n910 = n622 & n909;
  assign n911 = \V199(0)  & n597;
  assign n912 = ~n632 & n911;
  assign n913 = \V239(0)  & ~n597;
  assign n914 = n632 & n913;
  assign n915 = ~n912 & ~n914;
  assign n916 = ~n645 & ~n915;
  assign n917 = n541 & n916;
  assign n918 = ~n630 & n917;
  assign n919 = ~n622 & n918;
  assign n920 = ~n622 & n919;
  assign n921 = ~n910 & ~n920;
  assign n922 = ~n619 & ~n921;
  assign n923 = n616 & n922;
  assign \V1243(5)  = n904 | n923;
  assign n925 = \V84(2)  & n619;
  assign n926 = ~n616 & n925;
  assign n927 = \V32(9)  & ~n625;
  assign n928 = ~n625 & n927;
  assign n929 = \V32(6)  & n625;
  assign n930 = ~n928 & ~n929;
  assign n931 = n622 & ~n930;
  assign n932 = n622 & n931;
  assign n933 = \V194(4)  & n597;
  assign n934 = ~n632 & n933;
  assign n935 = \V234(4)  & ~n597;
  assign n936 = n632 & n935;
  assign n937 = ~n934 & ~n936;
  assign n938 = ~n645 & ~n937;
  assign n939 = n541 & n938;
  assign n940 = ~n630 & n939;
  assign n941 = ~n622 & n940;
  assign n942 = ~n622 & n941;
  assign n943 = ~n932 & ~n942;
  assign n944 = ~n619 & ~n943;
  assign n945 = n616 & n944;
  assign \V1243(4)  = n926 | n945;
  assign n947 = \V802(0)  & ~n632;
  assign n948 = \V244(0)  & \V243(0) ;
  assign n949 = ~\V245(0)  & n948;
  assign n950 = ~n947 & n949;
  assign n951 = \V245(0)  & ~n948;
  assign n952 = ~n947 & n951;
  assign \V597(0)  = n950 | n952;
  assign n954 = ~\V259(0)  & ~\V59(0) ;
  assign n955 = ~\V260(0)  & n954;
  assign n956 = \V258(0)  & n955;
  assign n957 = \V262(0)  & \V14(0) ;
  assign n958 = ~n956 & n957;
  assign \V1679(0)  = ~n540 | n958;
  assign n960 = \V15(0)  & ~\V16(0) ;
  assign n961 = ~\V15(0)  & \V16(0) ;
  assign \V1758(0)  = n960 | n961;
  assign n963 = ~\V102(0)  & ~\V1758(0) ;
  assign n964 = ~\V110(0)  & ~n963;
  assign n965 = n519 & n964;
  assign n966 = ~\V149(6)  & n613;
  assign n967 = \V56(0)  & n966;
  assign n968 = ~\V108(4)  & n960;
  assign n969 = \V101(0)  & n968;
  assign n970 = \V110(0)  & ~n969;
  assign n971 = ~n967 & n970;
  assign n972 = \V14(0)  & n971;
  assign \V1968(0)  = n965 | n972;
  assign n974 = ~\V134(1)  & ~n614;
  assign n975 = ~n614 & n974;
  assign n976 = ~\V88(3)  & n614;
  assign n977 = n614 & n976;
  assign \V1771(1)  = n975 | n977;
  assign n979 = ~\V134(0)  & ~n614;
  assign n980 = ~n614 & n979;
  assign n981 = ~\V88(2)  & n614;
  assign n982 = n614 & n981;
  assign \V1771(0)  = n980 | n982;
  assign n984 = \V274(0)  & ~\V202(0) ;
  assign n985 = ~\V271(0)  & n984;
  assign \V640(0)  = \V271(0)  | n985;
  assign V1423 = \V1(0)  & \V9(0) ;
  assign V1258 = \V9(0)  & \V2(0) ;
  assign n989 = \V109(0)  & ~\V13(0) ;
  assign V1431 = V1423 & ~n989;
  assign V787 = \V7(0)  & \V9(0) ;
  assign V778 = \V5(0)  & \V9(0) ;
  assign V780 = \V9(0)  & \V6(0) ;
  assign V1387 = \V8(0)  & \V9(0) ;
  assign V1259 = \V9(0)  & \V3(0) ;
  assign V1263 = \V4(0)  & \V9(0) ;
  assign n997 = \V71(0)  & \V202(0) ;
  assign n998 = ~\V13(0)  & n997;
  assign n999 = \V9(0)  & ~n998;
  assign V789 = \V4(0)  & n999;
  assign n1001 = ~V1263 & ~V789;
  assign n1002 = ~V1259 & n1001;
  assign n1003 = ~V1387 & n1002;
  assign n1004 = ~V780 & n1003;
  assign n1005 = ~V778 & n1004;
  assign n1006 = ~V787 & n1005;
  assign n1007 = ~V1431 & n1006;
  assign n1008 = ~V1258 & n1007;
  assign n1009 = ~V1423 & n1008;
  assign \V375(0)  = V1423 | ~n1009;
  assign n1011 = \V245(0)  & n948;
  assign n1012 = ~\V246(0)  & n1011;
  assign n1013 = ~n947 & n1012;
  assign n1014 = \V246(0)  & ~n1011;
  assign n1015 = ~n947 & n1014;
  assign \V603(0)  = n1013 | n1015;
  assign n1017 = \V149(3)  & n610;
  assign n1018 = n504 & n1017;
  assign n1019 = ~\V149(4)  & n1018;
  assign n1020 = ~\V149(6)  & n1019;
  assign n1021 = \V56(0)  & n1020;
  assign n1022 = \V108(4)  & ~n1021;
  assign \V1900(0)  = n960 | n1022;
  assign n1024 = ~n504 & ~n519;
  assign n1025 = n831 & ~n1024;
  assign n1026 = \V290(0)  & n1025;
  assign n1027 = \V165(4)  & n1026;
  assign n1028 = n1026 & n1027;
  assign n1029 = ~\V149(5)  & ~\V149(7) ;
  assign n1030 = ~\V149(3)  & n1029;
  assign n1031 = n504 & n1030;
  assign n1032 = ~\V149(4)  & n1031;
  assign n1033 = \V149(6)  & n1032;
  assign n1034 = \V56(0)  & n1033;
  assign n1035 = \V14(0)  & ~n1034;
  assign n1036 = \V100(2)  & n1035;
  assign n1037 = ~n1026 & n1036;
  assign n1038 = ~n1026 & n1037;
  assign \V1709(1)  = n1028 | n1038;
  assign n1040 = \V165(3)  & n1026;
  assign n1041 = n1026 & n1040;
  assign n1042 = \V100(1)  & n1035;
  assign n1043 = ~n1026 & n1042;
  assign n1044 = ~n1026 & n1043;
  assign \V1709(0)  = n1041 | n1044;
  assign n1046 = \V165(6)  & n1026;
  assign n1047 = n1026 & n1046;
  assign n1048 = \V100(4)  & n1035;
  assign n1049 = ~n1026 & n1048;
  assign n1050 = ~n1026 & n1049;
  assign \V1709(3)  = n1047 | n1050;
  assign n1052 = \V165(5)  & n1026;
  assign n1053 = n1026 & n1052;
  assign n1054 = \V100(3)  & n1035;
  assign n1055 = ~n1026 & n1054;
  assign n1056 = ~n1026 & n1055;
  assign \V1709(2)  = n1053 | n1056;
  assign n1058 = \V165(7)  & n1026;
  assign n1059 = n1026 & n1058;
  assign n1060 = \V100(5)  & n1035;
  assign n1061 = ~n1026 & n1060;
  assign n1062 = ~n1026 & n1061;
  assign \V1709(4)  = n1059 | n1062;
  assign n1064 = \V288(1)  & \V288(0) ;
  assign n1065 = \V32(2)  & n619;
  assign n1066 = ~n616 & n1065;
  assign n1067 = \V183(2)  & n597;
  assign n1068 = ~n632 & n1067;
  assign n1069 = \V223(2)  & ~n597;
  assign n1070 = n632 & n1069;
  assign n1071 = ~n1068 & ~n1070;
  assign n1072 = ~n622 & ~n645;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = n541 & n1073;
  assign n1075 = ~n630 & n1074;
  assign n1076 = ~n622 & n1075;
  assign n1077 = ~n619 & n1076;
  assign n1078 = n616 & n1077;
  assign \V1213(2)  = n1066 | n1078;
  assign n1080 = \V288(7)  & ~\V288(6) ;
  assign n1081 = \V288(5)  & ~\V288(4) ;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n1080 & n1081;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = \V288(3)  & ~\V288(2) ;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = n1084 & n1085;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = \V288(1)  & ~\V288(0) ;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n1088 & n1089;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~n1088 & n1089;
  assign n1094 = ~n1084 & n1085;
  assign n1095 = ~n1080 & n1081;
  assign n1096 = ~\V288(7)  & \V288(6) ;
  assign n1097 = ~n1080 & ~n1096;
  assign n1098 = ~\V288(5)  & \V288(4) ;
  assign n1099 = n1097 & ~n1098;
  assign n1100 = ~n1097 & n1098;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n1095 & n1101;
  assign n1103 = ~n1095 & ~n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~\V288(3)  & \V288(2) ;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = n1104 & n1105;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = n1094 & n1108;
  assign n1110 = ~n1094 & ~n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~\V288(1)  & \V288(0) ;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n1111 & n1112;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = n1093 & n1115;
  assign n1117 = ~n1093 & ~n1115;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = n1092 & n1118;
  assign n1120 = ~n1092 & ~n1118;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = \V1213(2)  & n1121;
  assign n1123 = ~\V1213(2)  & ~n1121;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = \V32(0)  & n619;
  assign n1126 = ~n616 & n1125;
  assign n1127 = \V183(0)  & n597;
  assign n1128 = ~n632 & n1127;
  assign n1129 = \V223(0)  & ~n597;
  assign n1130 = n632 & n1129;
  assign n1131 = ~n1128 & ~n1130;
  assign n1132 = n1072 & ~n1131;
  assign n1133 = n541 & n1132;
  assign n1134 = ~n630 & n1133;
  assign n1135 = ~n622 & n1134;
  assign n1136 = ~n619 & n1135;
  assign n1137 = n616 & n1136;
  assign \V1213(0)  = n1126 | n1137;
  assign n1139 = ~\V288(7)  & ~\V288(6) ;
  assign n1140 = \V288(5)  & \V288(4) ;
  assign n1141 = n1139 & ~n1140;
  assign n1142 = ~n1139 & n1140;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = n1095 & n1097;
  assign n1145 = n1095 & n1098;
  assign n1146 = n1097 & n1098;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = ~n1144 & n1147;
  assign n1149 = ~n1143 & n1148;
  assign n1150 = n1143 & ~n1148;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = \V288(3)  & \V288(2) ;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1151 & n1152;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = n1094 & ~n1104;
  assign n1157 = n1094 & n1105;
  assign n1158 = ~n1104 & n1105;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n1156 & n1159;
  assign n1161 = ~n1155 & n1160;
  assign n1162 = n1155 & ~n1160;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1064 & ~n1163;
  assign n1165 = n1064 & n1163;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = n1093 & ~n1111;
  assign n1168 = n1093 & n1112;
  assign n1169 = ~n1111 & n1112;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1167 & n1170;
  assign n1172 = ~n1166 & n1171;
  assign n1173 = n1166 & ~n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n1119 & n1174;
  assign n1176 = ~n1163 & ~n1171;
  assign n1177 = n1064 & ~n1171;
  assign n1178 = n1064 & ~n1163;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~n1176 & n1179;
  assign n1181 = ~n1151 & ~n1160;
  assign n1182 = n1152 & ~n1160;
  assign n1183 = ~n1151 & n1152;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1181 & n1184;
  assign n1186 = n1139 & ~n1148;
  assign n1187 = n1140 & ~n1148;
  assign n1188 = n1139 & n1140;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1186 & n1189;
  assign n1191 = ~n1139 & ~n1190;
  assign n1192 = n1139 & n1190;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1185 & n1193;
  assign n1195 = n1185 & ~n1193;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1180 & n1196;
  assign n1198 = n1180 & ~n1196;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n1175 & n1199;
  assign n1201 = ~n1175 & ~n1199;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = \V1213(0)  & n1202;
  assign n1204 = ~\V1213(0)  & ~n1202;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = \V32(1)  & n619;
  assign n1207 = ~n616 & n1206;
  assign n1208 = \V183(1)  & n597;
  assign n1209 = ~n632 & n1208;
  assign n1210 = \V223(1)  & ~n597;
  assign n1211 = n632 & n1210;
  assign n1212 = ~n1209 & ~n1211;
  assign n1213 = n1072 & ~n1212;
  assign n1214 = n541 & n1213;
  assign n1215 = ~n630 & n1214;
  assign n1216 = ~n622 & n1215;
  assign n1217 = ~n619 & n1216;
  assign n1218 = n616 & n1217;
  assign \V1213(1)  = n1207 | n1218;
  assign n1220 = ~n1119 & ~n1174;
  assign n1221 = ~n1175 & ~n1220;
  assign n1222 = \V1213(1)  & n1221;
  assign n1223 = ~\V1213(1)  & ~n1221;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = \V32(3)  & n619;
  assign n1226 = ~n616 & n1225;
  assign n1227 = \V183(3)  & n597;
  assign n1228 = ~n632 & n1227;
  assign n1229 = \V223(3)  & ~n597;
  assign n1230 = n632 & n1229;
  assign n1231 = ~n1228 & ~n1230;
  assign n1232 = n1072 & ~n1231;
  assign n1233 = n541 & n1232;
  assign n1234 = ~n630 & n1233;
  assign n1235 = ~n622 & n1234;
  assign n1236 = ~n619 & n1235;
  assign n1237 = n616 & n1236;
  assign \V1213(3)  = n1226 | n1237;
  assign n1239 = ~n1092 & \V1213(3) ;
  assign n1240 = n1092 & ~\V1213(3) ;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = \V149(3)  & n1029;
  assign n1243 = n504 & n1242;
  assign n1244 = ~\V149(4)  & n1243;
  assign n1245 = ~\V149(6)  & n1244;
  assign n1246 = ~\V802(0)  & n1245;
  assign n1247 = n1241 & ~n1246;
  assign n1248 = n1224 & n1247;
  assign n1249 = n1205 & n1248;
  assign n1250 = n1124 & n1249;
  assign n1251 = n1064 & n1250;
  assign n1252 = ~\V288(1)  & ~\V288(0) ;
  assign n1253 = ~n1092 & ~n1112;
  assign n1254 = ~n1112 & n1253;
  assign n1255 = ~n1092 & n1112;
  assign n1256 = n1112 & n1255;
  assign n1257 = ~n1254 & ~n1256;
  assign n1258 = ~n1092 & n1121;
  assign n1259 = n1092 & ~n1121;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1112 & ~n1260;
  assign n1262 = ~n1112 & n1261;
  assign n1263 = n1112 & ~n1118;
  assign n1264 = n1112 & n1263;
  assign n1265 = ~n1262 & ~n1264;
  assign n1266 = n1257 & n1265;
  assign n1267 = ~n1257 & ~n1265;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~n1089 & ~n1268;
  assign n1270 = ~n1089 & n1269;
  assign n1271 = n1089 & ~n1118;
  assign n1272 = n1089 & n1271;
  assign n1273 = ~n1270 & ~n1272;
  assign n1274 = \V1213(2)  & n1273;
  assign n1275 = ~\V1213(2)  & ~n1273;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1221 & n1258;
  assign n1278 = ~n1221 & ~n1258;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1112 & ~n1279;
  assign n1281 = ~n1112 & n1280;
  assign n1282 = n1112 & ~n1174;
  assign n1283 = n1112 & n1282;
  assign n1284 = ~n1281 & ~n1283;
  assign n1285 = n1266 & n1284;
  assign n1286 = n1202 & n1277;
  assign n1287 = ~n1202 & ~n1277;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = ~n1112 & ~n1288;
  assign n1290 = ~n1112 & n1289;
  assign n1291 = n1112 & ~n1199;
  assign n1292 = n1112 & n1291;
  assign n1293 = ~n1290 & ~n1292;
  assign n1294 = n1285 & n1293;
  assign n1295 = ~n1285 & ~n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1089 & ~n1296;
  assign n1298 = ~n1089 & n1297;
  assign n1299 = n1089 & ~n1199;
  assign n1300 = n1089 & n1299;
  assign n1301 = ~n1298 & ~n1300;
  assign n1302 = \V1213(0)  & n1301;
  assign n1303 = ~\V1213(0)  & ~n1301;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = ~n1266 & ~n1284;
  assign n1306 = ~n1285 & ~n1305;
  assign n1307 = ~n1089 & ~n1306;
  assign n1308 = ~n1089 & n1307;
  assign n1309 = n1089 & ~n1174;
  assign n1310 = n1089 & n1309;
  assign n1311 = ~n1308 & ~n1310;
  assign n1312 = \V1213(1)  & n1311;
  assign n1313 = ~\V1213(1)  & ~n1311;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1089 & n1257;
  assign n1316 = ~n1089 & n1315;
  assign n1317 = n1089 & ~n1092;
  assign n1318 = n1089 & n1317;
  assign n1319 = ~n1316 & ~n1318;
  assign n1320 = \V1213(3)  & n1319;
  assign n1321 = ~\V1213(3)  & ~n1319;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1246 & n1322;
  assign n1324 = n1314 & n1323;
  assign n1325 = n1304 & n1324;
  assign n1326 = n1276 & n1325;
  assign n1327 = ~n1252 & n1326;
  assign n1328 = n1088 & n1111;
  assign n1329 = ~n1088 & ~n1111;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = \V1213(2)  & n1330;
  assign n1332 = ~\V1213(2)  & ~n1330;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = n1163 & n1328;
  assign n1335 = n1196 & n1334;
  assign n1336 = ~n1196 & ~n1334;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = \V1213(0)  & n1337;
  assign n1339 = ~\V1213(0)  & ~n1337;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = ~n1163 & ~n1328;
  assign n1342 = ~n1334 & ~n1341;
  assign n1343 = \V1213(1)  & n1342;
  assign n1344 = ~\V1213(1)  & ~n1342;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1088 & \V1213(3) ;
  assign n1347 = n1088 & ~\V1213(3) ;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1246 & n1348;
  assign n1350 = n1345 & n1349;
  assign n1351 = n1340 & n1350;
  assign n1352 = n1333 & n1351;
  assign n1353 = n1152 & n1352;
  assign n1354 = ~\V288(3)  & ~\V288(2) ;
  assign n1355 = ~n1088 & ~n1105;
  assign n1356 = ~n1105 & n1355;
  assign n1357 = ~n1088 & n1105;
  assign n1358 = n1105 & n1357;
  assign n1359 = ~n1356 & ~n1358;
  assign n1360 = ~n1088 & n1330;
  assign n1361 = n1088 & ~n1330;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1105 & ~n1362;
  assign n1364 = ~n1105 & n1363;
  assign n1365 = n1105 & ~n1111;
  assign n1366 = n1105 & n1365;
  assign n1367 = ~n1364 & ~n1366;
  assign n1368 = n1359 & n1367;
  assign n1369 = ~n1359 & ~n1367;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1085 & ~n1370;
  assign n1372 = ~n1085 & n1371;
  assign n1373 = n1085 & ~n1111;
  assign n1374 = n1085 & n1373;
  assign n1375 = ~n1372 & ~n1374;
  assign n1376 = \V1213(2)  & n1375;
  assign n1377 = ~\V1213(2)  & ~n1375;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = n1342 & n1360;
  assign n1380 = ~n1342 & ~n1360;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = ~n1105 & ~n1381;
  assign n1383 = ~n1105 & n1382;
  assign n1384 = n1105 & ~n1163;
  assign n1385 = n1105 & n1384;
  assign n1386 = ~n1383 & ~n1385;
  assign n1387 = n1368 & n1386;
  assign n1388 = n1337 & n1379;
  assign n1389 = ~n1337 & ~n1379;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = ~n1105 & ~n1390;
  assign n1392 = ~n1105 & n1391;
  assign n1393 = n1105 & ~n1196;
  assign n1394 = n1105 & n1393;
  assign n1395 = ~n1392 & ~n1394;
  assign n1396 = n1387 & n1395;
  assign n1397 = ~n1387 & ~n1395;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1085 & ~n1398;
  assign n1400 = ~n1085 & n1399;
  assign n1401 = n1085 & ~n1196;
  assign n1402 = n1085 & n1401;
  assign n1403 = ~n1400 & ~n1402;
  assign n1404 = \V1213(0)  & n1403;
  assign n1405 = ~\V1213(0)  & ~n1403;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1368 & ~n1386;
  assign n1408 = ~n1387 & ~n1407;
  assign n1409 = ~n1085 & ~n1408;
  assign n1410 = ~n1085 & n1409;
  assign n1411 = n1085 & ~n1163;
  assign n1412 = n1085 & n1411;
  assign n1413 = ~n1410 & ~n1412;
  assign n1414 = \V1213(1)  & n1413;
  assign n1415 = ~\V1213(1)  & ~n1413;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1085 & n1359;
  assign n1418 = ~n1085 & n1417;
  assign n1419 = n1085 & ~n1088;
  assign n1420 = n1085 & n1419;
  assign n1421 = ~n1418 & ~n1420;
  assign n1422 = \V1213(3)  & n1421;
  assign n1423 = ~\V1213(3)  & ~n1421;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1246 & n1424;
  assign n1426 = n1416 & n1425;
  assign n1427 = n1406 & n1426;
  assign n1428 = n1378 & n1427;
  assign n1429 = ~n1354 & n1428;
  assign n1430 = \V1213(2)  & n1367;
  assign n1431 = ~\V1213(2)  & ~n1367;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = \V1213(0)  & n1395;
  assign n1434 = ~\V1213(0)  & ~n1395;
  assign n1435 = ~n1433 & ~n1434;
  assign n1436 = \V1213(1)  & n1386;
  assign n1437 = ~\V1213(1)  & ~n1386;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = \V1213(3)  & n1359;
  assign n1440 = ~\V1213(3)  & ~n1359;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~n1246 & n1441;
  assign n1443 = n1438 & n1442;
  assign n1444 = n1435 & n1443;
  assign n1445 = n1432 & n1444;
  assign n1446 = \V288(2)  & n1445;
  assign n1447 = \V1213(2)  & n1111;
  assign n1448 = ~\V1213(2)  & ~n1111;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = \V1213(0)  & n1196;
  assign n1451 = ~\V1213(0)  & ~n1196;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = n1163 & \V1213(1) ;
  assign n1454 = ~n1163 & ~\V1213(1) ;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = n1088 & \V1213(3) ;
  assign n1457 = ~n1088 & ~\V1213(3) ;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1246 & n1458;
  assign n1460 = n1455 & n1459;
  assign n1461 = n1452 & n1460;
  assign n1462 = n1449 & n1461;
  assign n1463 = n1152 & n1462;
  assign n1464 = \V1213(2)  & n1265;
  assign n1465 = ~\V1213(2)  & ~n1265;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = \V1213(0)  & n1293;
  assign n1468 = ~\V1213(0)  & ~n1293;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = \V1213(1)  & n1284;
  assign n1471 = ~\V1213(1)  & ~n1284;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = \V1213(3)  & n1257;
  assign n1474 = ~\V1213(3)  & ~n1257;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n1246 & n1475;
  assign n1477 = n1472 & n1476;
  assign n1478 = n1469 & n1477;
  assign n1479 = n1466 & n1478;
  assign n1480 = \V288(0)  & n1479;
  assign n1481 = \V1213(2)  & n1118;
  assign n1482 = ~\V1213(2)  & ~n1118;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = \V1213(0)  & n1199;
  assign n1485 = ~\V1213(0)  & ~n1199;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n1174 & \V1213(1) ;
  assign n1488 = ~n1174 & ~\V1213(1) ;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = n1092 & \V1213(3) ;
  assign n1491 = ~n1092 & ~\V1213(3) ;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1246 & n1492;
  assign n1494 = n1489 & n1493;
  assign n1495 = n1486 & n1494;
  assign n1496 = n1483 & n1495;
  assign n1497 = n1064 & n1496;
  assign n1498 = ~n1480 & ~n1497;
  assign n1499 = ~n1463 & n1498;
  assign n1500 = ~n1446 & n1499;
  assign n1501 = ~n1429 & n1500;
  assign n1502 = ~n1353 & n1501;
  assign n1503 = ~n1327 & n1502;
  assign n1504 = ~n1251 & n1503;
  assign n1505 = \V56(0)  & n549;
  assign n1506 = \V149(7)  & n1505;
  assign n1507 = n549 & n798;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~\V88(3)  & n562;
  assign n1510 = \V88(3)  & n570;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n598 & ~n1511;
  assign n1513 = \V149(4)  & n581;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = \V56(0)  & ~n1514;
  assign n1516 = ~\V172(0)  & n1515;
  assign n1517 = ~\V274(0)  & ~\V271(0) ;
  assign n1518 = \V278(0)  & ~n632;
  assign n1519 = \V56(0)  & ~n597;
  assign n1520 = \V171(0)  & n1519;
  assign n1521 = ~n1518 & ~n1520;
  assign n1522 = \V177(0)  & n1521;
  assign n1523 = ~\V248(0)  & n1522;
  assign n1524 = ~n797 & n1523;
  assign n1525 = n598 & ~n1511;
  assign n1526 = \V59(0)  & n1525;
  assign n1527 = ~n1524 & ~n1526;
  assign n1528 = ~n1517 & n1527;
  assign n1529 = ~n1516 & n1528;
  assign n1530 = n829 & ~n1529;
  assign \V1536(0)  = ~n1508 | ~n1530;
  assign n1532 = ~n1504 & ~\V1536(0) ;
  assign n1533 = \V56(0)  & ~n515;
  assign n1534 = n829 & n1533;
  assign n1535 = \V1536(0)  & ~n1534;
  assign \V1512(1)  = n1532 | n1535;
  assign n1537 = n1084 & n1104;
  assign n1538 = ~n1084 & ~n1104;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = \V1213(2)  & n1539;
  assign n1541 = ~\V1213(2)  & ~n1539;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = n1151 & n1537;
  assign n1544 = n1193 & n1543;
  assign n1545 = ~n1193 & ~n1543;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = \V1213(0)  & n1546;
  assign n1548 = ~\V1213(0)  & ~n1546;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1151 & ~n1537;
  assign n1551 = ~n1543 & ~n1550;
  assign n1552 = \V1213(1)  & n1551;
  assign n1553 = ~\V1213(1)  & ~n1551;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1084 & \V1213(3) ;
  assign n1556 = n1084 & ~\V1213(3) ;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1246 & n1557;
  assign n1559 = n1554 & n1558;
  assign n1560 = n1549 & n1559;
  assign n1561 = n1542 & n1560;
  assign n1562 = n1140 & n1561;
  assign n1563 = \V1213(2)  & ~n1246;
  assign n1564 = ~\V1213(1)  & n1563;
  assign n1565 = ~\V1213(0)  & n1564;
  assign n1566 = ~\V1213(3)  & n1565;
  assign n1567 = \V288(6)  & n1566;
  assign n1568 = \V288(7)  & n1567;
  assign n1569 = ~\V1213(1)  & ~n1246;
  assign n1570 = ~\V1213(0)  & n1569;
  assign n1571 = \V1213(2)  & n1570;
  assign n1572 = \V1213(3)  & n1571;
  assign n1573 = \V288(6)  & n1572;
  assign n1574 = \V288(7)  & n1573;
  assign n1575 = \V1213(2)  & n1104;
  assign n1576 = ~\V1213(2)  & ~n1104;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = \V1213(0)  & n1193;
  assign n1579 = ~\V1213(0)  & ~n1193;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = n1151 & \V1213(1) ;
  assign n1582 = ~n1151 & ~\V1213(1) ;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = n1084 & \V1213(3) ;
  assign n1585 = ~n1084 & ~\V1213(3) ;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~n1246 & n1586;
  assign n1588 = n1583 & n1587;
  assign n1589 = n1580 & n1588;
  assign n1590 = n1577 & n1589;
  assign n1591 = n1140 & n1590;
  assign n1592 = ~n1463 & ~n1497;
  assign n1593 = ~n1591 & n1592;
  assign n1594 = ~n1574 & n1593;
  assign n1595 = ~n1568 & n1594;
  assign n1596 = ~n1562 & n1595;
  assign n1597 = ~n1353 & n1596;
  assign n1598 = ~n1251 & n1597;
  assign n1599 = ~\V1536(0)  & ~n1598;
  assign n1600 = n829 & \V1536(0) ;
  assign \V1512(3)  = n1599 | n1600;
  assign n1602 = ~\V288(5)  & ~\V288(4) ;
  assign n1603 = ~n1084 & ~n1098;
  assign n1604 = ~n1098 & n1603;
  assign n1605 = ~n1084 & n1098;
  assign n1606 = n1098 & n1605;
  assign n1607 = ~n1604 & ~n1606;
  assign n1608 = ~n1084 & n1539;
  assign n1609 = n1084 & ~n1539;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = ~n1098 & ~n1610;
  assign n1612 = ~n1098 & n1611;
  assign n1613 = n1098 & ~n1104;
  assign n1614 = n1098 & n1613;
  assign n1615 = ~n1612 & ~n1614;
  assign n1616 = n1607 & n1615;
  assign n1617 = ~n1607 & ~n1615;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = ~n1081 & ~n1618;
  assign n1620 = ~n1081 & n1619;
  assign n1621 = n1081 & ~n1104;
  assign n1622 = n1081 & n1621;
  assign n1623 = ~n1620 & ~n1622;
  assign n1624 = \V1213(2)  & n1623;
  assign n1625 = ~\V1213(2)  & ~n1623;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = n1551 & n1608;
  assign n1628 = ~n1551 & ~n1608;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~n1098 & ~n1629;
  assign n1631 = ~n1098 & n1630;
  assign n1632 = n1098 & ~n1151;
  assign n1633 = n1098 & n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign n1635 = n1616 & n1634;
  assign n1636 = n1546 & n1627;
  assign n1637 = ~n1546 & ~n1627;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1098 & ~n1638;
  assign n1640 = ~n1098 & n1639;
  assign n1641 = n1098 & ~n1193;
  assign n1642 = n1098 & n1641;
  assign n1643 = ~n1640 & ~n1642;
  assign n1644 = n1635 & n1643;
  assign n1645 = ~n1635 & ~n1643;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = ~n1081 & ~n1646;
  assign n1648 = ~n1081 & n1647;
  assign n1649 = n1081 & ~n1193;
  assign n1650 = n1081 & n1649;
  assign n1651 = ~n1648 & ~n1650;
  assign n1652 = \V1213(0)  & n1651;
  assign n1653 = ~\V1213(0)  & ~n1651;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1616 & ~n1634;
  assign n1656 = ~n1635 & ~n1655;
  assign n1657 = ~n1081 & ~n1656;
  assign n1658 = ~n1081 & n1657;
  assign n1659 = n1081 & ~n1151;
  assign n1660 = n1081 & n1659;
  assign n1661 = ~n1658 & ~n1660;
  assign n1662 = \V1213(1)  & n1661;
  assign n1663 = ~\V1213(1)  & ~n1661;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1081 & n1607;
  assign n1666 = ~n1081 & n1665;
  assign n1667 = n1081 & ~n1084;
  assign n1668 = n1081 & n1667;
  assign n1669 = ~n1666 & ~n1668;
  assign n1670 = \V1213(3)  & n1669;
  assign n1671 = ~\V1213(3)  & ~n1669;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~n1246 & n1672;
  assign n1674 = n1664 & n1673;
  assign n1675 = n1654 & n1674;
  assign n1676 = n1626 & n1675;
  assign n1677 = ~n1602 & n1676;
  assign n1678 = \V1213(2)  & n1615;
  assign n1679 = ~\V1213(2)  & ~n1615;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = \V1213(0)  & n1643;
  assign n1682 = ~\V1213(0)  & ~n1643;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = \V1213(1)  & n1634;
  assign n1685 = ~\V1213(1)  & ~n1634;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = \V1213(3)  & n1607;
  assign n1688 = ~\V1213(3)  & ~n1607;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1246 & n1689;
  assign n1691 = n1686 & n1690;
  assign n1692 = n1683 & n1691;
  assign n1693 = n1680 & n1692;
  assign n1694 = \V288(4)  & n1693;
  assign n1695 = n1498 & ~n1591;
  assign n1696 = ~n1694 & n1695;
  assign n1697 = ~n1677 & n1696;
  assign n1698 = ~n1562 & n1697;
  assign n1699 = ~n1327 & n1698;
  assign n1700 = ~n1251 & n1699;
  assign n1701 = ~\V1536(0)  & ~n1700;
  assign n1702 = n829 & ~n1533;
  assign n1703 = ~n1508 & n1702;
  assign n1704 = \V1536(0)  & ~n1703;
  assign \V1512(2)  = n1701 | n1704;
  assign n1706 = \V108(2)  & ~n1021;
  assign n1707 = n523 & n809;
  assign \V1898(0)  = n1706 | n1707;
  assign n1709 = ~n488 & ~n589;
  assign n1710 = ~n484 & n1709;
  assign n1711 = n591 & ~n1710;
  assign n1712 = ~\V289(0)  & n541;
  assign n1713 = ~\V249(0)  & n1712;
  assign n1714 = ~n1711 & n1713;
  assign n1715 = \V295(0)  & n1714;
  assign \V1652(0)  = \V290(0)  | ~n1715;
  assign n1717 = \V199(2)  & \V199(4) ;
  assign n1718 = \V199(0)  & n1717;
  assign n1719 = \V194(3)  & n1718;
  assign n1720 = \V194(1)  & n1719;
  assign n1721 = \V194(2)  & n1720;
  assign n1722 = \V194(4)  & n1721;
  assign n1723 = \V199(1)  & n1722;
  assign n1724 = \V199(3)  & n1723;
  assign n1725 = \V194(0)  & n1724;
  assign n1726 = ~n632 & n1725;
  assign n1727 = ~\V1536(0)  & n1726;
  assign n1728 = \V242(0)  & \V14(0) ;
  assign n1729 = n631 & n1728;
  assign \V1726(0)  = n1727 | n1729;
  assign n1731 = \V149(6)  & n1244;
  assign n1732 = \V149(4)  & n1031;
  assign n1733 = ~\V149(6)  & n1732;
  assign n1734 = \V118(5)  & ~n1733;
  assign n1735 = n966 & n1734;
  assign n1736 = ~n1731 & n1735;
  assign n1737 = \V132(7)  & n1733;
  assign n1738 = ~n966 & n1737;
  assign n1739 = ~n1731 & n1738;
  assign \V1953(7)  = n1736 | n1739;
  assign n1741 = \V118(4)  & ~n1733;
  assign n1742 = n966 & n1741;
  assign n1743 = ~n1731 & n1742;
  assign n1744 = \V132(6)  & n1733;
  assign n1745 = ~n966 & n1744;
  assign n1746 = ~n1731 & n1745;
  assign \V1953(6)  = n1743 | n1746;
  assign n1748 = \V15(0)  & \V16(0) ;
  assign \V1757(0)  = n960 | n1748;
  assign n1750 = ~n578 & ~n598;
  assign n1751 = n588 & ~n1525;
  assign n1752 = ~n1750 & n1751;
  assign n1753 = \V59(0)  & ~n1752;
  assign n1754 = \V62(0)  & n599;
  assign n1755 = ~n1515 & ~n1754;
  assign n1756 = ~n1753 & n1755;
  assign n1757 = ~n831 & ~n1756;
  assign \V410(0)  = \V1757(0)  | ~n1757;
  assign n1759 = \V132(1)  & n1733;
  assign n1760 = ~n966 & n1759;
  assign \V1953(1)  = ~n1731 & n1760;
  assign n1762 = \V108(5)  & ~n1733;
  assign n1763 = ~n966 & n1762;
  assign n1764 = n1731 & n1763;
  assign n1765 = \V132(0)  & n1733;
  assign n1766 = ~n966 & n1765;
  assign n1767 = ~n1731 & n1766;
  assign \V1953(0)  = n1764 | n1767;
  assign n1769 = \V118(1)  & ~n1733;
  assign n1770 = n966 & n1769;
  assign n1771 = ~n1731 & n1770;
  assign n1772 = \V132(3)  & n1733;
  assign n1773 = ~n966 & n1772;
  assign n1774 = ~n1731 & n1773;
  assign \V1953(3)  = n1771 | n1774;
  assign n1776 = \V118(0)  & ~n1733;
  assign n1777 = n966 & n1776;
  assign n1778 = ~n1731 & n1777;
  assign n1779 = \V132(2)  & n1733;
  assign n1780 = ~n966 & n1779;
  assign n1781 = ~n1731 & n1780;
  assign \V1953(2)  = n1778 | n1781;
  assign n1783 = \V118(3)  & ~n1733;
  assign n1784 = n966 & n1783;
  assign n1785 = ~n1731 & n1784;
  assign n1786 = \V132(5)  & n1733;
  assign n1787 = ~n966 & n1786;
  assign n1788 = ~n1731 & n1787;
  assign \V1953(5)  = n1785 | n1788;
  assign n1790 = \V118(2)  & ~n1733;
  assign n1791 = n966 & n1790;
  assign n1792 = ~n1731 & n1791;
  assign n1793 = \V132(4)  & n1733;
  assign n1794 = ~n966 & n1793;
  assign n1795 = ~n1731 & n1794;
  assign \V1953(4)  = n1792 | n1795;
  assign n1797 = \V149(6)  & n802;
  assign n1798 = ~\V149(4)  & n512;
  assign n1799 = \V149(6)  & n1798;
  assign n1800 = ~n1797 & ~n1799;
  assign n1801 = \V56(0)  & ~n1800;
  assign n1802 = \V62(0)  & n1799;
  assign n1803 = n579 & ~n598;
  assign n1804 = ~\V149(6)  & n1798;
  assign n1805 = ~n549 & ~n551;
  assign n1806 = ~n589 & n1805;
  assign n1807 = \V802(0)  & ~n1806;
  assign n1808 = \V149(6)  & n1732;
  assign n1809 = ~n614 & ~n1804;
  assign n1810 = ~n1808 & n1809;
  assign n1811 = \V56(0)  & ~n1810;
  assign n1812 = ~n1807 & ~n1811;
  assign n1813 = \V78(0)  & ~\V78(1) ;
  assign n1814 = ~\V78(0)  & \V78(1) ;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = \V78(2)  & ~\V78(3) ;
  assign n1817 = ~\V78(2)  & \V78(3) ;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1815 & n1818;
  assign n1820 = n1815 & ~n1818;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = \V78(4)  & ~\V78(5) ;
  assign n1823 = ~\V78(4)  & \V78(5) ;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = \V84(0)  & ~\V84(1) ;
  assign n1826 = ~\V84(0)  & \V84(1) ;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = ~n1824 & n1827;
  assign n1829 = n1824 & ~n1827;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~n1821 & n1830;
  assign n1832 = n1821 & ~n1830;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~\V94(0)  & ~n1833;
  assign n1835 = \V94(0)  & n1833;
  assign n1836 = ~n1834 & ~n1835;
  assign n1837 = \V84(2)  & ~\V84(3) ;
  assign n1838 = ~\V84(2)  & \V84(3) ;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = \V84(4)  & ~\V84(5) ;
  assign n1841 = ~\V84(4)  & \V84(5) ;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1839 & n1842;
  assign n1844 = n1839 & ~n1842;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = \V88(0)  & ~\V88(1) ;
  assign n1847 = ~\V88(0)  & \V88(1) ;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = \V88(2)  & ~\V88(3) ;
  assign n1850 = ~\V88(2)  & \V88(3) ;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = ~n1848 & n1851;
  assign n1853 = n1848 & ~n1851;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1845 & n1854;
  assign n1856 = n1845 & ~n1854;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~\V94(1)  & ~n1857;
  assign n1859 = \V94(1)  & n1857;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1836 & ~n1860;
  assign n1862 = ~n1812 & ~n1861;
  assign n1863 = n1804 & ~n1862;
  assign n1864 = ~n589 & ~n1863;
  assign n1865 = ~n1803 & n1864;
  assign n1866 = ~n550 & n1865;
  assign n1867 = ~n484 & n1866;
  assign n1868 = \V56(0)  & ~n1867;
  assign n1869 = \V59(0)  & n601;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = ~n1802 & n1870;
  assign \V508(0)  = n1801 | ~n1871;
  assign n1873 = \V14(0)  & n837;
  assign n1874 = ~n1799 & n1873;
  assign n1875 = \V65(0)  & n1874;
  assign n1876 = ~n599 & n1875;
  assign n1877 = V763 & n1873;
  assign n1878 = ~\V165(5)  & n1877;
  assign n1879 = \V165(3)  & n1878;
  assign n1880 = ~\V165(4)  & n1879;
  assign n1881 = \V165(6)  & n1880;
  assign n1882 = \V70(0)  & n1881;
  assign \V1392(0)  = n1876 | n1882;
  assign n1884 = \V32(10)  & n619;
  assign n1885 = ~n616 & n1884;
  assign n1886 = \V32(3)  & ~n625;
  assign n1887 = ~n625 & n1886;
  assign n1888 = \V32(0)  & n625;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = n622 & ~n1889;
  assign n1891 = n622 & n1890;
  assign n1892 = \V189(4)  & n597;
  assign n1893 = ~n632 & n1892;
  assign n1894 = \V229(4)  & ~n597;
  assign n1895 = n632 & n1894;
  assign n1896 = ~n1893 & ~n1895;
  assign n1897 = n541 & ~n1896;
  assign n1898 = ~n630 & n1897;
  assign n1899 = ~n645 & n1898;
  assign n1900 = \V257(5)  & ~n541;
  assign n1901 = ~n630 & n1900;
  assign n1902 = n645 & n1901;
  assign n1903 = ~n1899 & ~n1902;
  assign n1904 = ~n622 & ~n1903;
  assign n1905 = ~n622 & n1904;
  assign n1906 = ~n1891 & ~n1905;
  assign n1907 = ~n619 & ~n1906;
  assign n1908 = n616 & n1907;
  assign \V1213(10)  = n1885 | n1908;
  assign n1910 = ~\V37(0)  & ~\V1213(10) ;
  assign n1911 = ~\V37(0)  & n1910;
  assign n1912 = \V37(0)  & ~\V1243(7) ;
  assign n1913 = \V37(0)  & n1912;
  assign \V1829(7)  = n1911 | n1913;
  assign n1915 = \V32(9)  & n619;
  assign n1916 = ~n616 & n1915;
  assign n1917 = \V32(2)  & ~n625;
  assign n1918 = ~n625 & n1917;
  assign n1919 = ~n625 & ~n1918;
  assign n1920 = n622 & ~n1919;
  assign n1921 = n622 & n1920;
  assign n1922 = \V189(3)  & n597;
  assign n1923 = ~n632 & n1922;
  assign n1924 = \V229(3)  & ~n597;
  assign n1925 = n632 & n1924;
  assign n1926 = ~n1923 & ~n1925;
  assign n1927 = n541 & ~n1926;
  assign n1928 = ~n630 & n1927;
  assign n1929 = ~n645 & n1928;
  assign n1930 = \V257(4)  & ~n541;
  assign n1931 = ~n630 & n1930;
  assign n1932 = n645 & n1931;
  assign n1933 = ~n1929 & ~n1932;
  assign n1934 = ~n622 & ~n1933;
  assign n1935 = ~n622 & n1934;
  assign n1936 = ~n1921 & ~n1935;
  assign n1937 = ~n619 & ~n1936;
  assign n1938 = n616 & n1937;
  assign \V1213(9)  = n1916 | n1938;
  assign n1940 = ~\V37(0)  & ~\V1213(9) ;
  assign n1941 = ~\V37(0)  & n1940;
  assign n1942 = \V37(0)  & ~\V1243(6) ;
  assign n1943 = \V37(0)  & n1942;
  assign \V1829(6)  = n1941 | n1943;
  assign n1945 = ~\V37(0)  & \V321(2) ;
  assign n1946 = ~\V37(0)  & n1945;
  assign n1947 = \V37(0)  & ~\V1243(9) ;
  assign n1948 = \V37(0)  & n1947;
  assign \V1829(9)  = n1946 | n1948;
  assign n1950 = \V32(11)  & n619;
  assign n1951 = ~n616 & n1950;
  assign n1952 = \V32(4)  & ~n625;
  assign n1953 = ~n625 & n1952;
  assign n1954 = \V32(1)  & n625;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = n622 & ~n1955;
  assign n1957 = n622 & n1956;
  assign n1958 = \V189(5)  & n597;
  assign n1959 = ~n632 & n1958;
  assign n1960 = \V229(5)  & ~n597;
  assign n1961 = n632 & n1960;
  assign n1962 = ~n1959 & ~n1961;
  assign n1963 = n541 & ~n1962;
  assign n1964 = ~n630 & n1963;
  assign n1965 = ~n645 & n1964;
  assign n1966 = \V257(6)  & ~n541;
  assign n1967 = ~n630 & n1966;
  assign n1968 = n645 & n1967;
  assign n1969 = ~n1965 & ~n1968;
  assign n1970 = ~n622 & ~n1969;
  assign n1971 = ~n622 & n1970;
  assign n1972 = ~n1957 & ~n1971;
  assign n1973 = ~n619 & ~n1972;
  assign n1974 = n616 & n1973;
  assign \V1213(11)  = n1951 | n1974;
  assign n1976 = ~\V37(0)  & ~\V1213(11) ;
  assign n1977 = ~\V37(0)  & n1976;
  assign n1978 = \V37(0)  & ~\V1243(8) ;
  assign n1979 = \V37(0)  & n1978;
  assign \V1829(8)  = n1977 | n1979;
  assign n1981 = \V290(0)  & n831;
  assign n1982 = n523 & n1981;
  assign n1983 = n551 & n598;
  assign n1984 = ~\V302(0)  & n549;
  assign n1985 = ~n796 & ~n1984;
  assign n1986 = ~n1983 & n1985;
  assign n1987 = ~n803 & n1986;
  assign n1988 = ~\V289(0)  & \V14(0) ;
  assign n1989 = ~n1987 & n1988;
  assign n1990 = n798 & n1989;
  assign n1991 = ~n831 & n1990;
  assign n1992 = n523 & ~n831;
  assign n1993 = n798 & n1992;
  assign n1994 = ~n1991 & n1993;
  assign n1995 = ~n509 & n1994;
  assign n1996 = ~n1982 & ~n1995;
  assign n1997 = ~\V165(5)  & ~\V165(7) ;
  assign n1998 = ~\V165(3)  & n1997;
  assign n1999 = ~\V165(4)  & n1998;
  assign n2000 = ~\V165(6)  & n1999;
  assign n2001 = ~n798 & ~n2000;
  assign n2002 = ~n1996 & ~n2001;
  assign n2003 = ~n1996 & n2002;
  assign n2004 = ~\V149(4)  & n612;
  assign n2005 = ~\V149(6)  & n2004;
  assign n2006 = \V56(0)  & n2005;
  assign n2007 = \V14(0)  & ~n2006;
  assign n2008 = \V213(0)  & n2007;
  assign n2009 = n1996 & n2008;
  assign n2010 = n1996 & n2009;
  assign \V1281(0)  = n2003 | n2010;
  assign n2012 = \V174(0)  & ~n829;
  assign n2013 = ~\V302(0)  & \V292(0) ;
  assign n2014 = \V174(0)  & n831;
  assign n2015 = ~n501 & ~n2014;
  assign n2016 = ~n2013 & n2015;
  assign \V1620(0)  = n2012 | ~n2016;
  assign n2018 = \V32(4)  & n619;
  assign n2019 = ~n616 & n2018;
  assign n2020 = \V183(4)  & n597;
  assign n2021 = ~n632 & n2020;
  assign n2022 = \V223(4)  & ~n597;
  assign n2023 = n632 & n2022;
  assign n2024 = ~n2021 & ~n2023;
  assign n2025 = n541 & ~n2024;
  assign n2026 = ~n630 & n2025;
  assign n2027 = ~n645 & n2026;
  assign n2028 = ~n1968 & ~n2027;
  assign n2029 = ~n622 & ~n2028;
  assign n2030 = ~n622 & n2029;
  assign n2031 = ~n619 & n2030;
  assign n2032 = n616 & n2031;
  assign \V1213(4)  = n2019 | n2032;
  assign n2034 = ~\V37(0)  & ~\V1213(4) ;
  assign n2035 = ~\V37(0)  & n2034;
  assign n2036 = \V37(0)  & ~\V1243(1) ;
  assign n2037 = \V37(0)  & n2036;
  assign \V1829(1)  = n2035 | n2037;
  assign n2039 = \V37(0)  & ~\V1213(2) ;
  assign n2040 = \V37(0)  & n2039;
  assign \V1829(0)  = n1946 | n2040;
  assign n2042 = \V32(6)  & n619;
  assign n2043 = ~n616 & n2042;
  assign n2044 = n622 & n625;
  assign n2045 = n622 & n2044;
  assign n2046 = \V189(0)  & n597;
  assign n2047 = ~n632 & n2046;
  assign n2048 = \V229(0)  & ~n597;
  assign n2049 = n632 & n2048;
  assign n2050 = ~n2047 & ~n2049;
  assign n2051 = n541 & ~n2050;
  assign n2052 = ~n630 & n2051;
  assign n2053 = ~n645 & n2052;
  assign n2054 = \V257(1)  & ~n541;
  assign n2055 = ~n630 & n2054;
  assign n2056 = n645 & n2055;
  assign n2057 = ~n2053 & ~n2056;
  assign n2058 = ~n622 & ~n2057;
  assign n2059 = ~n622 & n2058;
  assign n2060 = ~n2045 & ~n2059;
  assign n2061 = ~n619 & ~n2060;
  assign n2062 = n616 & n2061;
  assign \V1213(6)  = n2043 | n2062;
  assign n2064 = ~\V37(0)  & ~\V1213(6) ;
  assign n2065 = ~\V37(0)  & n2064;
  assign n2066 = \V37(0)  & ~\V1243(3) ;
  assign n2067 = \V37(0)  & n2066;
  assign \V1829(3)  = n2065 | n2067;
  assign n2069 = \V32(5)  & n619;
  assign n2070 = ~n616 & n2069;
  assign n2071 = n622 & ~n625;
  assign n2072 = n622 & n2071;
  assign n2073 = \V183(5)  & n597;
  assign n2074 = ~n632 & n2073;
  assign n2075 = \V223(5)  & ~n597;
  assign n2076 = n632 & n2075;
  assign n2077 = ~n2074 & ~n2076;
  assign n2078 = n541 & ~n2077;
  assign n2079 = ~n630 & n2078;
  assign n2080 = ~n645 & n2079;
  assign n2081 = \V257(0)  & ~n541;
  assign n2082 = ~n630 & n2081;
  assign n2083 = n645 & n2082;
  assign n2084 = ~n2080 & ~n2083;
  assign n2085 = ~n622 & ~n2084;
  assign n2086 = ~n622 & n2085;
  assign n2087 = ~n2072 & ~n2086;
  assign n2088 = ~n619 & ~n2087;
  assign n2089 = n616 & n2088;
  assign \V1213(5)  = n2070 | n2089;
  assign n2091 = ~\V37(0)  & ~\V1213(5) ;
  assign n2092 = ~\V37(0)  & n2091;
  assign n2093 = \V37(0)  & ~\V1243(2) ;
  assign n2094 = \V37(0)  & n2093;
  assign \V1829(2)  = n2092 | n2094;
  assign n2096 = ~n831 & ~n1024;
  assign n2097 = n798 & n2096;
  assign n2098 = ~n1991 & n2097;
  assign n2099 = ~n509 & n2098;
  assign n2100 = ~n1026 & ~n2099;
  assign n2101 = ~n2001 & ~n2100;
  assign n2102 = ~n2100 & n2101;
  assign n2103 = \V100(0)  & n1035;
  assign n2104 = n2100 & n2103;
  assign n2105 = n2100 & n2104;
  assign \V1693(0)  = n2102 | n2105;
  assign n2107 = \V32(8)  & n619;
  assign n2108 = ~n616 & n2107;
  assign n2109 = \V32(1)  & ~n625;
  assign n2110 = ~n625 & n2109;
  assign n2111 = ~n625 & ~n2110;
  assign n2112 = n622 & ~n2111;
  assign n2113 = n622 & n2112;
  assign n2114 = \V189(2)  & n597;
  assign n2115 = ~n632 & n2114;
  assign n2116 = \V229(2)  & ~n597;
  assign n2117 = n632 & n2116;
  assign n2118 = ~n2115 & ~n2117;
  assign n2119 = n541 & ~n2118;
  assign n2120 = ~n630 & n2119;
  assign n2121 = ~n645 & n2120;
  assign n2122 = \V257(3)  & ~n541;
  assign n2123 = ~n630 & n2122;
  assign n2124 = n645 & n2123;
  assign n2125 = ~n2121 & ~n2124;
  assign n2126 = ~n622 & ~n2125;
  assign n2127 = ~n622 & n2126;
  assign n2128 = ~n2113 & ~n2127;
  assign n2129 = ~n619 & ~n2128;
  assign n2130 = n616 & n2129;
  assign \V1213(8)  = n2108 | n2130;
  assign n2132 = ~\V37(0)  & ~\V1213(8) ;
  assign n2133 = ~\V37(0)  & n2132;
  assign n2134 = \V37(0)  & ~\V1243(5) ;
  assign n2135 = \V37(0)  & n2134;
  assign \V1829(5)  = n2133 | n2135;
  assign n2137 = \V32(7)  & n619;
  assign n2138 = ~n616 & n2137;
  assign n2139 = \V32(0)  & ~n625;
  assign n2140 = ~n625 & n2139;
  assign n2141 = ~n625 & ~n2140;
  assign n2142 = n622 & ~n2141;
  assign n2143 = n622 & n2142;
  assign n2144 = \V189(1)  & n597;
  assign n2145 = ~n632 & n2144;
  assign n2146 = \V229(1)  & ~n597;
  assign n2147 = n632 & n2146;
  assign n2148 = ~n2145 & ~n2147;
  assign n2149 = n541 & ~n2148;
  assign n2150 = ~n630 & n2149;
  assign n2151 = ~n645 & n2150;
  assign n2152 = \V257(2)  & ~n541;
  assign n2153 = ~n630 & n2152;
  assign n2154 = n645 & n2153;
  assign n2155 = ~n2151 & ~n2154;
  assign n2156 = ~n622 & ~n2155;
  assign n2157 = ~n622 & n2156;
  assign n2158 = ~n2143 & ~n2157;
  assign n2159 = ~n619 & ~n2158;
  assign n2160 = n616 & n2159;
  assign \V1213(7)  = n2138 | n2160;
  assign n2162 = ~\V37(0)  & ~\V1213(7) ;
  assign n2163 = ~\V37(0)  & n2162;
  assign n2164 = \V37(0)  & ~\V1243(4) ;
  assign n2165 = \V37(0)  & n2164;
  assign \V1829(4)  = n2163 | n2165;
  assign n2167 = \V108(1)  & ~n1033;
  assign n2168 = ~n2005 & n2167;
  assign n2169 = ~n1733 & n2168;
  assign n2170 = n1020 & n2169;
  assign n2171 = \V124(1)  & ~n1033;
  assign n2172 = ~n2005 & n2171;
  assign n2173 = n1733 & n2172;
  assign n2174 = ~n1020 & n2173;
  assign n2175 = \V213(1)  & ~n1033;
  assign n2176 = n2005 & n2175;
  assign n2177 = ~n1733 & n2176;
  assign n2178 = ~n1020 & n2177;
  assign n2179 = \V100(1)  & n1033;
  assign n2180 = ~n2005 & n2179;
  assign n2181 = ~n1733 & n2180;
  assign n2182 = ~n1020 & n2181;
  assign n2183 = ~n2178 & ~n2182;
  assign n2184 = ~n2174 & n2183;
  assign \V1921(1)  = n2170 | ~n2184;
  assign n2186 = \V108(0)  & ~n1033;
  assign n2187 = ~n2005 & n2186;
  assign n2188 = ~n1733 & n2187;
  assign n2189 = n1020 & n2188;
  assign n2190 = \V124(0)  & ~n1033;
  assign n2191 = ~n2005 & n2190;
  assign n2192 = n1733 & n2191;
  assign n2193 = ~n1020 & n2192;
  assign n2194 = \V213(0)  & ~n1033;
  assign n2195 = n2005 & n2194;
  assign n2196 = ~n1733 & n2195;
  assign n2197 = ~n1020 & n2196;
  assign n2198 = \V100(0)  & n1033;
  assign n2199 = ~n2005 & n2198;
  assign n2200 = ~n1733 & n2199;
  assign n2201 = ~n1020 & n2200;
  assign n2202 = ~n2197 & ~n2201;
  assign n2203 = ~n2193 & n2202;
  assign \V1921(0)  = n2189 | ~n2203;
  assign n2205 = \V108(3)  & ~n1033;
  assign n2206 = ~n2005 & n2205;
  assign n2207 = ~n1733 & n2206;
  assign n2208 = n1020 & n2207;
  assign n2209 = \V124(3)  & ~n1033;
  assign n2210 = ~n2005 & n2209;
  assign n2211 = n1733 & n2210;
  assign n2212 = ~n1020 & n2211;
  assign n2213 = \V213(3)  & ~n1033;
  assign n2214 = n2005 & n2213;
  assign n2215 = ~n1733 & n2214;
  assign n2216 = ~n1020 & n2215;
  assign n2217 = \V100(3)  & n1033;
  assign n2218 = ~n2005 & n2217;
  assign n2219 = ~n1733 & n2218;
  assign n2220 = ~n1020 & n2219;
  assign n2221 = ~n2216 & ~n2220;
  assign n2222 = ~n2212 & n2221;
  assign \V1921(3)  = n2208 | ~n2222;
  assign n2224 = \V108(2)  & ~n1033;
  assign n2225 = ~n2005 & n2224;
  assign n2226 = ~n1733 & n2225;
  assign n2227 = n1020 & n2226;
  assign n2228 = \V124(2)  & ~n1033;
  assign n2229 = ~n2005 & n2228;
  assign n2230 = n1733 & n2229;
  assign n2231 = ~n1020 & n2230;
  assign n2232 = \V213(2)  & ~n1033;
  assign n2233 = n2005 & n2232;
  assign n2234 = ~n1733 & n2233;
  assign n2235 = ~n1020 & n2234;
  assign n2236 = \V100(2)  & n1033;
  assign n2237 = ~n2005 & n2236;
  assign n2238 = ~n1733 & n2237;
  assign n2239 = ~n1020 & n2238;
  assign n2240 = ~n2235 & ~n2239;
  assign n2241 = ~n2231 & n2240;
  assign \V1921(2)  = n2227 | ~n2241;
  assign n2243 = \V124(5)  & ~n1033;
  assign n2244 = ~n2005 & n2243;
  assign n2245 = n1733 & n2244;
  assign n2246 = ~n1020 & n2245;
  assign n2247 = \V213(5)  & ~n1033;
  assign n2248 = n2005 & n2247;
  assign n2249 = ~n1733 & n2248;
  assign n2250 = ~n1020 & n2249;
  assign n2251 = \V100(5)  & n1033;
  assign n2252 = ~n2005 & n2251;
  assign n2253 = ~n1733 & n2252;
  assign n2254 = ~n1020 & n2253;
  assign n2255 = ~n2250 & ~n2254;
  assign \V1921(5)  = n2246 | ~n2255;
  assign n2257 = \V108(4)  & ~n1033;
  assign n2258 = ~n2005 & n2257;
  assign n2259 = ~n1733 & n2258;
  assign n2260 = n1020 & n2259;
  assign n2261 = \V124(4)  & ~n1033;
  assign n2262 = ~n2005 & n2261;
  assign n2263 = n1733 & n2262;
  assign n2264 = ~n1020 & n2263;
  assign n2265 = \V213(4)  & ~n1033;
  assign n2266 = n2005 & n2265;
  assign n2267 = ~n1733 & n2266;
  assign n2268 = ~n1020 & n2267;
  assign n2269 = \V100(4)  & n1033;
  assign n2270 = ~n2005 & n2269;
  assign n2271 = ~n1733 & n2270;
  assign n2272 = ~n1020 & n2271;
  assign n2273 = ~n2268 & ~n2272;
  assign n2274 = ~n2264 & n2273;
  assign \V1921(4)  = n2260 | ~n2274;
  assign n2276 = \V802(0)  & n550;
  assign n2277 = ~\V279(0)  & ~n2276;
  assign n2278 = ~\V280(0)  & n2277;
  assign n2279 = \V149(4)  & n2276;
  assign n2280 = \V280(0)  & ~n2276;
  assign n2281 = \V279(0)  & n2280;
  assign n2282 = ~n2279 & ~n2281;
  assign \V826(0)  = n2278 | ~n2282;
  assign n2284 = ~\V244(0)  & \V243(0) ;
  assign n2285 = ~n947 & n2284;
  assign n2286 = \V244(0)  & ~\V243(0) ;
  assign n2287 = ~n947 & n2286;
  assign \V591(0)  = n2285 | n2287;
  assign n2289 = \V56(0)  & n1731;
  assign n2290 = \V101(0)  & ~n2289;
  assign n2291 = \V14(0)  & n2290;
  assign n2292 = n519 & n961;
  assign n2293 = n523 & n961;
  assign n2294 = ~n2292 & ~n2293;
  assign \V1759(0)  = n2291 | ~n2294;
  assign n2296 = \V108(5)  & ~n2289;
  assign \V1901(0)  = n961 | n2296;
  assign n2298 = \V165(4)  & n1982;
  assign n2299 = n1982 & n2298;
  assign n2300 = \V213(2)  & n2007;
  assign n2301 = ~n1982 & n2300;
  assign n2302 = ~n1982 & n2301;
  assign \V1297(1)  = n2299 | n2302;
  assign n2304 = \V165(3)  & n1982;
  assign n2305 = n1982 & n2304;
  assign n2306 = \V213(1)  & n2007;
  assign n2307 = ~n1982 & n2306;
  assign n2308 = ~n1982 & n2307;
  assign \V1297(0)  = n2305 | n2308;
  assign n2310 = \V165(6)  & n1982;
  assign n2311 = n1982 & n2310;
  assign n2312 = \V213(4)  & n2007;
  assign n2313 = ~n1982 & n2312;
  assign n2314 = ~n1982 & n2313;
  assign \V1297(3)  = n2311 | n2314;
  assign n2316 = \V165(5)  & n1982;
  assign n2317 = n1982 & n2316;
  assign n2318 = \V213(3)  & n2007;
  assign n2319 = ~n1982 & n2318;
  assign n2320 = ~n1982 & n2319;
  assign \V1297(2)  = n2317 | n2320;
  assign n2322 = \V165(7)  & n1982;
  assign n2323 = n1982 & n2322;
  assign n2324 = \V213(5)  & n2007;
  assign n2325 = ~n1982 & n2324;
  assign n2326 = ~n1982 & n2325;
  assign \V1297(4)  = n2323 | n2326;
  assign n2328 = \V268(3)  & \V268(5) ;
  assign n2329 = \V268(1)  & n2328;
  assign n2330 = \V268(2)  & n2329;
  assign n2331 = \V268(4)  & n2330;
  assign n2332 = \V268(0)  & n2331;
  assign n2333 = ~\V56(0)  & ~\V50(0) ;
  assign n2334 = ~\V62(0)  & n2333;
  assign n2335 = ~n541 & ~n2334;
  assign n2336 = ~n2332 & ~n2335;
  assign n2337 = \V14(0)  & ~n2336;
  assign n2338 = ~\V258(0)  & n2337;
  assign n2339 = \V14(0)  & n2336;
  assign n2340 = \V258(0)  & n2339;
  assign \V1451(0)  = n2338 | n2340;
  assign n2342 = \V240(0)  & ~n831;
  assign V1719 = ~\V172(0)  & n2342;
  assign n2344 = ~\V248(0)  & n1724;
  assign n2345 = V1719 & n2344;
  assign n2346 = n541 & ~n1562;
  assign n2347 = ~n1591 & n2346;
  assign n2348 = n541 & ~n1677;
  assign n2349 = ~n1694 & n2348;
  assign n2350 = n2347 & n2349;
  assign n2351 = n1140 & ~n2350;
  assign n2352 = n541 & ~n1251;
  assign n2353 = ~n1497 & n2352;
  assign n2354 = n541 & ~n1327;
  assign n2355 = ~n1480 & n2354;
  assign n2356 = n2353 & n2355;
  assign n2357 = n1064 & ~n2356;
  assign n2358 = n541 & ~n1353;
  assign n2359 = ~n1463 & n2358;
  assign n2360 = n541 & ~n1429;
  assign n2361 = ~n1446 & n2360;
  assign n2362 = n2359 & n2361;
  assign n2363 = n1152 & ~n2362;
  assign n2364 = n541 & ~n1568;
  assign n2365 = ~n1574 & n2364;
  assign n2366 = \V1213(3)  & ~n1246;
  assign n2367 = ~\V1213(1)  & n2366;
  assign n2368 = ~\V1213(0)  & n2367;
  assign n2369 = ~\V1213(2)  & n2368;
  assign n2370 = \V288(6)  & n2369;
  assign n2371 = ~\V1213(3)  & ~n1246;
  assign n2372 = ~\V1213(1)  & n2371;
  assign n2373 = ~\V1213(0)  & n2372;
  assign n2374 = ~\V1213(2)  & n2373;
  assign n2375 = ~n1139 & n2374;
  assign n2376 = n541 & ~n2375;
  assign n2377 = ~n2370 & n2376;
  assign n2378 = n2365 & n2377;
  assign n2379 = \V288(6)  & ~n2378;
  assign n2380 = \V288(7)  & n2379;
  assign n2381 = ~n2363 & ~n2380;
  assign n2382 = ~n2357 & n2381;
  assign n2383 = ~n2351 & n2382;
  assign n2384 = ~\V248(0)  & ~n2383;
  assign n2385 = \V1243(8)  & n2384;
  assign n2386 = \V1243(7)  & n2385;
  assign n2387 = \V1243(9)  & n2386;
  assign n2388 = V1719 & n2387;
  assign n2389 = \V246(0)  & n1011;
  assign n2390 = ~\V248(0)  & n2389;
  assign n2391 = V1719 & n2390;
  assign n2392 = \V247(0)  & n2391;
  assign n2393 = ~n2388 & ~n2392;
  assign \V393(0)  = n2345 | ~n2393;
  assign n2395 = \V108(3)  & ~n1021;
  assign n2396 = n519 & n809;
  assign \V1899(0)  = n2395 | n2396;
  assign n2398 = ~n549 & \V1757(0) ;
  assign n2399 = \V802(0)  & \V1757(0) ;
  assign n2400 = n549 & n2399;
  assign n2401 = ~n1862 & ~n2400;
  assign \V1480(0)  = n2398 | ~n2401;
  assign n2403 = \V70(0)  & ~n541;
  assign n2404 = n541 & n1752;
  assign n2405 = \V59(0)  & ~n2404;
  assign n2406 = n541 & n588;
  assign n2407 = ~n579 & n2406;
  assign n2408 = n578 & n2407;
  assign n2409 = ~n550 & n2408;
  assign n2410 = \V802(0)  & ~n2409;
  assign n2411 = ~n599 & n1514;
  assign n2412 = ~n601 & n2411;
  assign n2413 = ~\V174(0)  & n2412;
  assign n2414 = \V56(0)  & ~n2413;
  assign n2415 = \V66(0)  & ~n831;
  assign n2416 = V763 & n2415;
  assign n2417 = ~\V215(0)  & n2416;
  assign n2418 = \V802(0)  & n776;
  assign n2419 = ~V1719 & ~n2418;
  assign n2420 = ~n2417 & n2419;
  assign n2421 = ~n2414 & n2420;
  assign n2422 = ~n2410 & n2421;
  assign n2423 = ~n2405 & n2422;
  assign n2424 = ~n1754 & n2423;
  assign \V423(0)  = n2403 | ~n2424;
  assign n2426 = ~\V68(0)  & ~\V70(0) ;
  assign n2427 = ~\V66(0)  & n2426;
  assign n2428 = ~\V69(0)  & n2427;
  assign n2429 = \V215(0)  & \V14(0) ;
  assign n2430 = ~n2428 & n2429;
  assign n2431 = n820 & n2430;
  assign n2432 = \V216(0)  & ~\V214(0) ;
  assign \V1492(0)  = n2431 | n2432;
  assign n2434 = n840 & V1719;
  assign n2435 = \V302(0)  & V1719;
  assign n2436 = n832 & V1719;
  assign n2437 = ~V763 & ~n598;
  assign n2438 = \V802(0)  & ~n2437;
  assign n2439 = ~n796 & ~n1797;
  assign n2440 = ~n1799 & n2439;
  assign n2441 = ~n1804 & n2440;
  assign n2442 = \V56(0)  & ~n2441;
  assign n2443 = \V802(0)  & n549;
  assign n2444 = ~n551 & ~n589;
  assign n2445 = \V802(0)  & ~n2444;
  assign n2446 = ~V763 & n2445;
  assign n2447 = \V149(6)  & n2004;
  assign n2448 = \V66(0)  & n2447;
  assign n2449 = \V66(0)  & V763;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = ~n2446 & n2450;
  assign n2452 = ~n2443 & n2451;
  assign n2453 = ~n2442 & n2452;
  assign n2454 = \V32(0)  & n1199;
  assign n2455 = ~\V32(0)  & ~n1199;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = \V32(1)  & n1174;
  assign n2458 = ~\V32(1)  & ~n1174;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = n1118 & n2459;
  assign n2461 = \V32(2)  & n2460;
  assign n2462 = n2456 & n2461;
  assign n2463 = \V32(1)  & n2456;
  assign n2464 = n1174 & n2463;
  assign n2465 = \V32(2)  & n1118;
  assign n2466 = ~\V32(2)  & ~n1118;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = n2456 & n2467;
  assign n2469 = \V32(3)  & n2468;
  assign n2470 = n1092 & n2469;
  assign n2471 = n2459 & n2470;
  assign n2472 = ~n2464 & ~n2471;
  assign n2473 = ~n2454 & n2472;
  assign n2474 = ~n2462 & n2473;
  assign n2475 = ~n2453 & ~n2474;
  assign n2476 = \V215(0)  & \V66(0) ;
  assign n2477 = ~\V214(0)  & ~\V43(0) ;
  assign n2478 = n541 & n2477;
  assign n2479 = ~n2476 & n2478;
  assign n2480 = ~n2475 & n2479;
  assign n2481 = ~\V1757(0)  & n2480;
  assign n2482 = ~n2438 & n2481;
  assign n2483 = ~n1862 & n2482;
  assign n2484 = ~n798 & n2483;
  assign n2485 = \V423(0)  & n2484;
  assign n2486 = ~n2436 & n2485;
  assign n2487 = ~n2435 & n2486;
  assign n2488 = ~n2345 & n2487;
  assign n2489 = ~n2388 & n2488;
  assign n2490 = ~n2434 & n2489;
  assign V432 = ~n2392 & n2490;
  assign n2492 = \V62(0)  & n614;
  assign n2493 = \V802(0)  & n1711;
  assign n2494 = \V59(0)  & n591;
  assign n2495 = ~n787 & n2494;
  assign n2496 = \V56(0)  & n614;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2493 & n2497;
  assign n2499 = ~\V270(0)  & n2498;
  assign n2500 = ~\V302(0)  & ~n2499;
  assign V630 = ~n2492 & n2500;
  assign \V435(0)  = V432 | V630;
  assign n2503 = ~\V78(3)  & n614;
  assign n2504 = n614 & n2503;
  assign n2505 = ~n614 & ~\V1213(11) ;
  assign n2506 = ~n614 & n2505;
  assign \V1781(1)  = n2504 | n2506;
  assign n2508 = ~\V78(2)  & n614;
  assign n2509 = n614 & n2508;
  assign n2510 = ~n614 & ~\V1213(10) ;
  assign n2511 = ~n614 & n2510;
  assign \V1781(0)  = n2509 | n2511;
  assign n2513 = ~\V13(0)  & \V10(0) ;
  assign V1256 = \V2(0)  & n2513;
  assign n2515 = ~\V60(0)  & ~\V63(0) ;
  assign n2516 = n614 & ~n2515;
  assign n2517 = ~n550 & n1511;
  assign n2518 = n578 & n2517;
  assign n2519 = ~n579 & n2518;
  assign n2520 = n588 & n2519;
  assign n2521 = ~n589 & n2520;
  assign n2522 = \V57(0)  & ~n2521;
  assign n2523 = ~\V57(0)  & n1804;
  assign n2524 = \V12(0)  & \V2(0) ;
  assign n2525 = ~\V174(0)  & n2524;
  assign n2526 = ~n2523 & n2525;
  assign n2527 = ~n2522 & n2526;
  assign n2528 = ~n2516 & n2527;
  assign V1257 = ~\V35(0)  & n2528;
  assign V1260 = \V11(0)  & \V3(0) ;
  assign V1261 = ~\V62(0)  & V1260;
  assign V1262 = \V4(0)  & n2513;
  assign V1264 = \V4(0)  & \V12(0) ;
  assign V1265 = \V52(0)  & V1264;
  assign V1266 = \V11(0)  & \V4(0) ;
  assign V1267 = \V11(0)  & \V2(0) ;
  assign n2537 = \V258(0)  & n2332;
  assign n2538 = \V259(0)  & n2537;
  assign n2539 = ~\V258(0)  & n2335;
  assign n2540 = ~\V259(0)  & n2539;
  assign n2541 = ~n2538 & ~n2540;
  assign n2542 = ~\V260(0)  & ~n2541;
  assign n2543 = \V14(0)  & n2542;
  assign n2544 = \V260(0)  & n2541;
  assign n2545 = \V14(0)  & n2544;
  assign \V1467(0)  = n2543 | n2545;
  assign n2547 = ~n1804 & n1873;
  assign n2548 = ~n803 & n2547;
  assign n2549 = ~n1525 & n2548;
  assign n2550 = n541 & n2549;
  assign n2551 = ~n1750 & n2550;
  assign n2552 = n588 & n2551;
  assign n2553 = ~n1797 & n2552;
  assign V1365 = \V62(0)  & n2553;
  assign n2555 = ~\V268(0)  & n2331;
  assign n2556 = \V268(0)  & ~n2331;
  assign V1370 = n2555 | n2556;
  assign n2558 = \V268(2)  & n2328;
  assign n2559 = \V268(4)  & n2558;
  assign n2560 = ~\V268(1)  & n2559;
  assign n2561 = \V268(1)  & ~n2559;
  assign V1371 = n2560 | n2561;
  assign n2563 = \V268(4)  & n2328;
  assign n2564 = ~\V268(2)  & n2563;
  assign n2565 = \V268(2)  & ~n2563;
  assign V1372 = n2564 | n2565;
  assign n2567 = \V268(5)  & \V268(4) ;
  assign n2568 = ~\V268(3)  & n2567;
  assign n2569 = \V268(3)  & ~n2567;
  assign V1373 = n2568 | n2569;
  assign n2571 = \V268(5)  & ~\V268(4) ;
  assign n2572 = ~\V268(5)  & \V268(4) ;
  assign V1374 = n2571 | n2572;
  assign n2574 = \V802(0)  & ~n631;
  assign V782 = \V7(0)  & n2513;
  assign V1378 = n2574 & V782;
  assign n2577 = \V248(0)  & ~\V802(0) ;
  assign n2578 = ~n790 & ~n2577;
  assign n2579 = ~n591 & n2578;
  assign n2580 = ~\V802(0)  & n2579;
  assign n2581 = n488 & n2580;
  assign n2582 = ~n1725 & n2581;
  assign n2583 = ~\V802(0)  & n591;
  assign n2584 = ~\V802(0)  & n1725;
  assign n2585 = ~n790 & ~n2584;
  assign n2586 = ~n631 & n2585;
  assign n2587 = ~n2583 & n2586;
  assign n2588 = ~n2577 & n2587;
  assign n2589 = \V271(0)  & ~n614;
  assign n2590 = ~\V274(0)  & n2589;
  assign n2591 = ~n1725 & n2590;
  assign n2592 = n591 & n2591;
  assign n2593 = \V134(0)  & n2592;
  assign n2594 = \V134(1)  & n2593;
  assign n2595 = ~n2588 & ~n2594;
  assign n2596 = ~n2582 & n2595;
  assign V1380 = V782 & ~n2596;
  assign n2598 = \V802(0)  & ~n1805;
  assign n2599 = ~n550 & ~n2598;
  assign n2600 = \V7(0)  & ~n2599;
  assign V1382 = n2513 & n2600;
  assign n2602 = \V56(0)  & ~n831;
  assign n2603 = n1808 & n2602;
  assign n2604 = ~n1862 & n2603;
  assign n2605 = \V7(0)  & n2604;
  assign V1384 = n2513 & n2605;
  assign n2607 = \V7(0)  & n2335;
  assign V1386 = n2513 & n2607;
  assign V1426 = \V1(0)  & n2513;
  assign V1428 = \V11(0)  & \V1(0) ;
  assign V1429 = \V12(0)  & \V1(0) ;
  assign n2612 = \V66(0)  & n837;
  assign V1432 = \V14(0)  & n2612;
  assign n2614 = \V14(0)  & ~n2447;
  assign n2615 = n837 & n2614;
  assign V1470 = \V67(0)  & n2615;
  assign n2617 = \V149(7)  & n2443;
  assign n2618 = ~n1991 & ~n2617;
  assign \V1645(0)  = n2475 | ~n2618;
  assign n2620 = \V68(0)  & n837;
  assign V1537 = \V14(0)  & n2620;
  assign n2622 = ~\V69(0)  & ~\V50(0) ;
  assign n2623 = n837 & ~n2622;
  assign V1539 = \V14(0)  & n2623;
  assign n2625 = ~\V289(0)  & n832;
  assign n2626 = ~\V802(0)  & n2625;
  assign n2627 = \V262(0)  & n958;
  assign n2628 = n540 & ~n2627;
  assign n2629 = ~\V149(6)  & n513;
  assign n2630 = ~n1808 & n2628;
  assign n2631 = ~n1733 & n2630;
  assign n2632 = ~n2005 & n2631;
  assign n2633 = ~n1033 & n2632;
  assign n2634 = ~n966 & n2633;
  assign n2635 = ~n2629 & n2634;
  assign n2636 = ~n1797 & ~n1804;
  assign n2637 = n2635 & n2636;
  assign n2638 = n2628 & n2637;
  assign n2639 = ~n1799 & n2638;
  assign n2640 = \V62(0)  & ~n2636;
  assign n2641 = \V65(0)  & n1799;
  assign n2642 = ~\V59(0)  & ~n541;
  assign n2643 = ~\V259(0)  & n2642;
  assign n2644 = ~\V260(0)  & n2643;
  assign n2645 = \V258(0)  & n2644;
  assign n2646 = ~n1808 & ~n2629;
  assign n2647 = ~n1733 & n2646;
  assign n2648 = ~n2645 & n2647;
  assign n2649 = ~n1033 & n2648;
  assign n2650 = ~n966 & n2649;
  assign n2651 = ~n2005 & n2650;
  assign n2652 = \V56(0)  & ~n2651;
  assign n2653 = ~n2641 & ~n2652;
  assign n2654 = ~n2640 & n2653;
  assign n2655 = ~\V289(0)  & n2654;
  assign n2656 = n829 & n2655;
  assign n2657 = ~n2639 & n2656;
  assign n2658 = ~n834 & n2657;
  assign n2659 = n801 & ~n831;
  assign n2660 = n807 & ~n831;
  assign n2661 = n812 & ~n831;
  assign n2662 = ~n815 & ~n2661;
  assign n2663 = ~n1981 & n2662;
  assign n2664 = ~n2660 & n2663;
  assign \V1741(0)  = n2659 | ~n2664;
  assign n2666 = ~\V289(0)  & n2635;
  assign n2667 = \V1741(0)  & n2666;
  assign n2668 = ~n2448 & ~n2667;
  assign n2669 = ~n2658 & n2668;
  assign V1669 = ~n2626 & n2669;
  assign n2671 = \V108(0)  & ~n1021;
  assign n2672 = ~n1862 & ~n2671;
  assign \V1896(0)  = n1748 | ~n2672;
  assign n2674 = n787 & n2625;
  assign n2675 = ~\V802(0)  & n2674;
  assign V1736 = ~\V290(0)  & n2675;
  assign n2677 = \V262(0)  & ~n958;
  assign n2678 = ~n2334 & n2677;
  assign n2679 = \V261(0)  & ~n2678;
  assign n2680 = ~n2332 & ~n2679;
  assign V1832 = \V14(0)  & ~n2680;
  assign n2682 = ~n2537 & ~n2539;
  assign n2683 = ~\V259(0)  & ~n2682;
  assign n2684 = \V14(0)  & n2683;
  assign n2685 = \V259(0)  & n2682;
  assign n2686 = \V14(0)  & n2685;
  assign \V1459(0)  = n2684 | n2686;
  assign n2688 = ~\V1953(3)  & \V1953(2) ;
  assign n2689 = \V1953(3)  & ~\V1953(2) ;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = ~\V1953(5)  & \V1953(4) ;
  assign n2692 = \V1953(5)  & ~\V1953(4) ;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = ~n2690 & n2693;
  assign n2695 = n2690 & ~n2693;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = ~\V1953(7)  & \V1953(6) ;
  assign n2698 = \V1953(7)  & ~\V1953(6) ;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = \V48(0)  & ~n966;
  assign n2701 = ~n1800 & n2700;
  assign n2702 = \V118(6)  & n966;
  assign n2703 = n1800 & n2702;
  assign \V1960(0)  = n2701 | n2703;
  assign n2705 = \V46(0)  & ~n966;
  assign n2706 = ~n1800 & n2705;
  assign n2707 = \V118(7)  & n966;
  assign n2708 = n1800 & n2707;
  assign \V1960(1)  = n2706 | n2708;
  assign n2710 = \V1960(0)  & ~\V1960(1) ;
  assign n2711 = ~\V1960(0)  & \V1960(1) ;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = ~n2699 & n2712;
  assign n2714 = n2699 & ~n2712;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = ~n2696 & n2715;
  assign n2717 = n2696 & ~n2715;
  assign \V1613(1)  = ~n2716 & ~n2717;
  assign n2719 = ~\V174(0)  & n509;
  assign n2720 = ~n484 & ~n1513;
  assign n2721 = ~n589 & n2720;
  assign n2722 = ~n1803 & n2721;
  assign n2723 = ~n1512 & n2722;
  assign n2724 = ~n488 & n2723;
  assign n2725 = ~n550 & n2724;
  assign n2726 = \V59(0)  & ~V1719;
  assign n2727 = ~n796 & n2726;
  assign n2728 = n2725 & n2727;
  assign n2729 = ~n2719 & n2728;
  assign n2730 = ~n1245 & n2729;
  assign n2731 = n837 & n2730;
  assign n2732 = \V14(0)  & n2731;
  assign n2733 = n601 & n1873;
  assign n2734 = \V62(0)  & n2733;
  assign \V1274(0)  = n2732 | n2734;
  assign n2736 = ~\V1921(1)  & \V1921(0) ;
  assign n2737 = \V1921(1)  & ~\V1921(0) ;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = ~\V1921(3)  & \V1921(2) ;
  assign n2740 = \V1921(3)  & ~\V1921(2) ;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = ~n2738 & n2741;
  assign n2743 = n2738 & ~n2741;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = ~\V1921(5)  & \V1921(4) ;
  assign n2746 = \V1921(5)  & ~\V1921(4) ;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = ~\V1953(1)  & \V1953(0) ;
  assign n2749 = \V1953(1)  & ~\V1953(0) ;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = ~n2747 & n2750;
  assign n2752 = n2747 & ~n2750;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2744 & n2753;
  assign n2755 = n2744 & ~n2753;
  assign \V1613(0)  = ~n2754 & ~n2755;
  assign \V1440(0)  = ~\V14(0)  | n591;
  assign n2758 = n484 & \V802(0) ;
  assign n2759 = ~\V802(0)  & ~n591;
  assign n2760 = ~n632 & n2759;
  assign n2761 = ~n2594 & ~n2760;
  assign n2762 = \V802(0)  & \V1243(3) ;
  assign n2763 = n589 & n2762;
  assign n2764 = n2761 & n2763;
  assign n2765 = ~n2758 & n2764;
  assign n2766 = \V802(0)  & n589;
  assign n2767 = \V194(4)  & n1718;
  assign n2768 = \V199(1)  & n2767;
  assign n2769 = \V199(3)  & n2768;
  assign n2770 = ~\V194(3)  & n2769;
  assign n2771 = \V194(3)  & ~n2769;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = ~n2758 & ~n2772;
  assign n2774 = ~n2761 & n2773;
  assign n2775 = ~n2766 & n2774;
  assign n2776 = \V149(7)  & \V802(0) ;
  assign n2777 = n484 & n2776;
  assign n2778 = n2761 & n2777;
  assign n2779 = ~n2766 & n2778;
  assign n2780 = ~n2775 & ~n2779;
  assign \V572(3)  = n2765 | ~n2780;
  assign n2782 = \V802(0)  & \V1243(2) ;
  assign n2783 = n589 & n2782;
  assign n2784 = n2761 & n2783;
  assign n2785 = ~n2758 & n2784;
  assign n2786 = \V194(4)  & n1719;
  assign n2787 = \V199(1)  & n2786;
  assign n2788 = \V199(3)  & n2787;
  assign n2789 = ~\V194(2)  & n2788;
  assign n2790 = \V194(2)  & ~n2788;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = ~n2758 & ~n2791;
  assign n2793 = ~n2761 & n2792;
  assign n2794 = ~n2766 & n2793;
  assign n2795 = \V149(6)  & \V802(0) ;
  assign n2796 = n484 & n2795;
  assign n2797 = n2761 & n2796;
  assign n2798 = ~n2766 & n2797;
  assign n2799 = ~n2794 & ~n2798;
  assign \V572(2)  = n2785 | ~n2799;
  assign n2801 = \V271(0)  & ~n985;
  assign n2802 = \V269(0)  & n2801;
  assign n2803 = \V274(0)  & ~\V640(0) ;
  assign \V634(0)  = ~n2802 & ~n2803;
  assign n2805 = \V199(1)  & n1717;
  assign n2806 = \V199(3)  & n2805;
  assign n2807 = ~\V199(0)  & n2806;
  assign n2808 = \V199(0)  & ~n2806;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n2758 & ~n2809;
  assign n2811 = ~n2761 & n2810;
  assign n2812 = ~n2766 & n2811;
  assign n2813 = \V802(0)  & \V1243(5) ;
  assign n2814 = n589 & n2813;
  assign n2815 = n2761 & n2814;
  assign n2816 = ~n2758 & n2815;
  assign \V572(5)  = n2812 | n2816;
  assign n2818 = \V199(1)  & n1718;
  assign n2819 = \V199(3)  & n2818;
  assign n2820 = ~\V194(4)  & n2819;
  assign n2821 = \V194(4)  & ~n2819;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = ~n2758 & ~n2822;
  assign n2824 = ~n2761 & n2823;
  assign n2825 = ~n2766 & n2824;
  assign n2826 = \V802(0)  & \V1243(4) ;
  assign n2827 = n589 & n2826;
  assign n2828 = n2761 & n2827;
  assign n2829 = ~n2758 & n2828;
  assign \V572(4)  = n2825 | n2829;
  assign n2831 = \V277(0)  & ~n589;
  assign n2832 = \V14(0)  & n2831;
  assign \V1439(0)  = n2629 | n2832;
  assign n2834 = \V802(0)  & \V1243(1) ;
  assign n2835 = n589 & n2834;
  assign n2836 = n2761 & n2835;
  assign n2837 = ~n2758 & n2836;
  assign n2838 = \V194(2)  & n1719;
  assign n2839 = \V194(4)  & n2838;
  assign n2840 = \V199(1)  & n2839;
  assign n2841 = \V199(3)  & n2840;
  assign n2842 = ~\V194(1)  & n2841;
  assign n2843 = \V194(1)  & ~n2841;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = ~n2758 & ~n2844;
  assign n2846 = ~n2761 & n2845;
  assign n2847 = ~n2766 & n2846;
  assign n2848 = \V149(5)  & \V802(0) ;
  assign n2849 = n484 & n2848;
  assign n2850 = n2761 & n2849;
  assign n2851 = ~n2766 & n2850;
  assign n2852 = ~n2847 & ~n2851;
  assign \V572(1)  = n2837 | ~n2852;
  assign n2854 = \V802(0)  & ~\V321(2) ;
  assign n2855 = n589 & n2854;
  assign n2856 = n2761 & n2855;
  assign n2857 = ~n2758 & n2856;
  assign n2858 = ~\V194(0)  & n1724;
  assign n2859 = \V194(0)  & ~n1724;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = ~n2758 & ~n2860;
  assign n2862 = ~n2761 & n2861;
  assign n2863 = ~n2766 & n2862;
  assign n2864 = \V149(4)  & \V802(0) ;
  assign n2865 = n484 & n2864;
  assign n2866 = n2761 & n2865;
  assign n2867 = ~n2766 & n2866;
  assign n2868 = ~n2863 & ~n2867;
  assign \V572(0)  = n2857 | ~n2868;
  assign n2870 = \V45(0)  & ~\V43(0) ;
  assign \V511(0)  = \V40(0)  | n2870;
  assign n2872 = \V199(3)  & \V199(4) ;
  assign n2873 = ~\V199(2)  & n2872;
  assign n2874 = \V199(2)  & ~n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = ~n2758 & ~n2875;
  assign n2877 = ~n2761 & n2876;
  assign n2878 = ~n2766 & n2877;
  assign n2879 = \V802(0)  & \V1243(7) ;
  assign n2880 = n589 & n2879;
  assign n2881 = n2761 & n2880;
  assign n2882 = ~n2758 & n2881;
  assign \V572(7)  = n2878 | n2882;
  assign n2884 = \V199(3)  & n1717;
  assign n2885 = ~\V199(1)  & n2884;
  assign n2886 = \V199(1)  & ~n2884;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = ~n2758 & ~n2887;
  assign n2889 = ~n2761 & n2888;
  assign n2890 = ~n2766 & n2889;
  assign n2891 = \V802(0)  & \V1243(6) ;
  assign n2892 = n589 & n2891;
  assign n2893 = n2761 & n2892;
  assign n2894 = ~n2758 & n2893;
  assign \V572(6)  = n2890 | n2894;
  assign n2896 = ~\V199(4)  & ~n2758;
  assign n2897 = ~n2761 & n2896;
  assign n2898 = ~n2766 & n2897;
  assign n2899 = \V802(0)  & \V1243(9) ;
  assign n2900 = n589 & n2899;
  assign n2901 = n2761 & n2900;
  assign n2902 = ~n2758 & n2901;
  assign \V572(9)  = n2898 | n2902;
  assign n2904 = ~\V199(3)  & \V199(4) ;
  assign n2905 = \V199(3)  & ~\V199(4) ;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~n2758 & ~n2906;
  assign n2908 = ~n2761 & n2907;
  assign n2909 = ~n2766 & n2908;
  assign n2910 = \V802(0)  & \V1243(8) ;
  assign n2911 = n589 & n2910;
  assign n2912 = n2761 & n2911;
  assign n2913 = ~n2758 & n2912;
  assign \V572(8)  = n2909 | n2913;
  assign n2915 = ~n2574 & n2590;
  assign n2916 = \V134(1)  & ~n2590;
  assign n2917 = ~n2574 & n2916;
  assign n2918 = ~n2915 & n2917;
  assign n2919 = ~n2574 & ~n2590;
  assign n2920 = ~\V134(1)  & ~n2574;
  assign n2921 = n2590 & n2920;
  assign n2922 = ~n2919 & n2921;
  assign \V1992(1)  = n2918 | n2922;
  assign n2924 = \V134(0)  & ~n2590;
  assign n2925 = ~n2574 & n2924;
  assign n2926 = ~n2915 & n2925;
  assign n2927 = ~\V134(1)  & \V134(0) ;
  assign n2928 = \V134(1)  & ~\V134(0) ;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = ~n2574 & ~n2929;
  assign n2931 = n2590 & n2930;
  assign n2932 = ~n2919 & n2931;
  assign \V1992(0)  = n2926 | n2932;
  assign n2934 = ~\V247(0)  & n2389;
  assign n2935 = ~n947 & n2934;
  assign n2936 = \V247(0)  & ~n2389;
  assign n2937 = ~n947 & n2936;
  assign \V609(0)  = n2935 | n2937;
  assign n2939 = ~\V294(0)  & ~n1799;
  assign n2940 = ~n1863 & n2939;
  assign n2941 = \V59(0)  & \V91(0) ;
  assign n2942 = \V62(0)  & \V91(1) ;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n1804 & ~n2943;
  assign n2945 = ~\V41(0)  & \V45(0) ;
  assign n2946 = \V41(0)  & ~\V45(0) ;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2944 & n2947;
  assign \V1629(0)  = n2940 | ~n2948;
  assign n2950 = n837 & ~n840;
  assign n2951 = ~n787 & ~n2950;
  assign n2952 = ~n832 & ~n2654;
  assign n2953 = ~\V1741(0)  & n2952;
  assign n2954 = \V290(0)  & ~n831;
  assign n2955 = ~\V302(0)  & ~n2954;
  assign n2956 = ~\V289(0)  & n2955;
  assign n2957 = ~n2953 & n2956;
  assign n2958 = ~n2951 & n2957;
  assign n2959 = ~\V214(0)  & n2958;
  assign n2960 = ~n834 & n2959;
  assign n2961 = ~\V149(2)  & \V149(0) ;
  assign n2962 = \V149(1)  & n2961;
  assign n2963 = ~\V149(6)  & n1032;
  assign n2964 = ~n1020 & ~n1245;
  assign n2965 = n504 & n2964;
  assign n2966 = \V149(3)  & n2965;
  assign n2967 = ~n1731 & n2966;
  assign n2968 = ~\V149(3)  & ~\V149(7) ;
  assign n2969 = \V149(4)  & n2968;
  assign n2970 = n504 & n2969;
  assign n2971 = \V149(5)  & n2970;
  assign n2972 = ~\V149(6)  & n2971;
  assign n2973 = ~n2967 & ~n2972;
  assign n2974 = ~n2963 & n2973;
  assign n2975 = ~\V149(1)  & \V149(0) ;
  assign n2976 = \V149(2)  & n2975;
  assign n2977 = \V149(2)  & \V149(0) ;
  assign n2978 = \V149(1)  & n2977;
  assign n2979 = ~n2976 & ~n2978;
  assign n2980 = n2974 & n2979;
  assign n2981 = ~n2962 & n2980;
  assign n2982 = ~\V302(0)  & ~n2974;
  assign n2983 = n541 & ~n2982;
  assign n2984 = ~n2981 & n2983;
  assign n2985 = \V14(0)  & ~n2984;
  assign \V798(0)  = ~n2960 | ~n2985;
  assign n2987 = \V248(0)  & V1719;
  assign n2988 = ~\V423(0)  & ~n2987;
  assign n2989 = ~\V214(0)  & ~n2438;
  assign n2990 = ~n2988 & n2989;
  assign n2991 = ~\V43(0)  & n2990;
  assign n2992 = ~n2436 & n2991;
  assign n2993 = ~n2435 & n2992;
  assign n2994 = ~n2345 & n2993;
  assign n2995 = ~n2388 & n2994;
  assign n2996 = ~n2434 & n2995;
  assign \V398(0)  = n2392 | ~n2996;
  assign n2998 = \V33(0)  & ~n509;
  assign n2999 = \V289(0)  & n2998;
  assign \V1745(0)  = n523 | ~n2999;
  assign n3001 = n541 & ~n1246;
  assign n3002 = ~n1327 & n3001;
  assign n3003 = ~n1429 & n3002;
  assign n3004 = ~n1677 & n3003;
  assign n3005 = ~n2375 & n3004;
  assign n3006 = ~n1568 & n3005;
  assign n3007 = ~n1562 & n3006;
  assign n3008 = ~n1353 & n3007;
  assign V356 = ~n1251 & n3008;
  assign n3010 = n541 & ~n1480;
  assign n3011 = ~n1446 & n3010;
  assign n3012 = ~n1694 & n3011;
  assign n3013 = ~n2370 & n3012;
  assign n3014 = ~n1574 & n3013;
  assign n3015 = ~n1591 & n3014;
  assign n3016 = ~n1463 & n3015;
  assign V357 = ~n1497 & n3016;
  assign V373 = \V13(0)  & \V10(0) ;
  assign n3019 = ~\V35(0)  & ~n840;
  assign V377 = \V203(0)  & ~n3019;
  assign n3021 = \V108(1)  & ~n1021;
  assign n3022 = n589 & n1862;
  assign \V1897(0)  = n3021 | n3022;
  assign n3024 = ~\V39(0)  & \V38(0) ;
  assign n3025 = \V39(0)  & ~\V38(0) ;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = \V44(0)  & ~\V42(0) ;
  assign n3028 = ~\V44(0)  & \V42(0) ;
  assign n3029 = ~n3027 & ~n3028;
  assign V512 = n3026 & n3029;
  assign n3031 = \V59(0)  & ~n588;
  assign n3032 = \V56(0)  & n1512;
  assign n3033 = \V56(0)  & n1513;
  assign n3034 = \V59(0)  & ~n598;
  assign n3035 = ~n578 & n3034;
  assign n3036 = ~n1754 & ~n3035;
  assign n3037 = ~n3033 & n3036;
  assign n3038 = ~n3032 & n3037;
  assign n3039 = ~n1526 & n3038;
  assign n3040 = ~n3031 & n3039;
  assign n3041 = ~\V214(0)  & ~n798;
  assign n3042 = ~n3040 & n3041;
  assign n3043 = ~n831 & n3042;
  assign V527 = ~\V43(0)  & n3043;
  assign V537 = n589 & \V1213(0) ;
  assign V538 = n589 & \V1213(1) ;
  assign V539 = n589 & \V1213(2) ;
  assign V540 = n589 & \V1213(3) ;
  assign V541 = n589 & \V1213(4) ;
  assign V542 = n589 & \V1213(5) ;
  assign V543 = n589 & \V1213(6) ;
  assign V544 = n589 & \V1213(7) ;
  assign V545 = n589 & \V1213(8) ;
  assign V546 = n589 & \V1213(9) ;
  assign V547 = n589 & \V1213(10) ;
  assign V548 = n589 & \V1213(11) ;
  assign V587 = ~\V243(0)  & ~n947;
  assign n3058 = ~n601 & ~n1863;
  assign n3059 = \V59(0)  & ~\V214(0) ;
  assign n3060 = ~n3058 & n3059;
  assign n3061 = ~n831 & n3060;
  assign n3062 = ~n798 & ~n831;
  assign n3063 = n1868 & n3062;
  assign n3064 = ~\V214(0)  & n3063;
  assign n3065 = \V62(0)  & ~\V214(0) ;
  assign n3066 = n1799 & n3065;
  assign n3067 = ~n831 & n3066;
  assign n3068 = ~n3064 & ~n3067;
  assign V620 = ~n3061 & n3068;
  assign V621 = \V293(0)  & n2947;
  assign n3071 = \V257(5)  & \V257(7) ;
  assign n3072 = \V257(3)  & n3071;
  assign n3073 = \V257(1)  & n3072;
  assign n3074 = \V257(2)  & n3073;
  assign n3075 = \V257(4)  & n3074;
  assign n3076 = \V257(6)  & n3075;
  assign n3077 = ~\V257(0)  & n3076;
  assign n3078 = \V257(0)  & ~n3076;
  assign V650 = n3077 | n3078;
  assign n3080 = \V257(2)  & n3072;
  assign n3081 = \V257(4)  & n3080;
  assign n3082 = \V257(6)  & n3081;
  assign n3083 = ~\V257(1)  & n3082;
  assign n3084 = \V257(1)  & ~n3082;
  assign V651 = n3083 | n3084;
  assign n3086 = \V257(4)  & n3072;
  assign n3087 = \V257(6)  & n3086;
  assign n3088 = ~\V257(2)  & n3087;
  assign n3089 = \V257(2)  & ~n3087;
  assign V652 = n3088 | n3089;
  assign n3091 = \V257(4)  & n3071;
  assign n3092 = \V257(6)  & n3091;
  assign n3093 = ~\V257(3)  & n3092;
  assign n3094 = \V257(3)  & ~n3092;
  assign V653 = n3093 | n3094;
  assign n3096 = \V257(6)  & n3071;
  assign n3097 = ~\V257(4)  & n3096;
  assign n3098 = \V257(4)  & ~n3096;
  assign V654 = n3097 | n3098;
  assign n3100 = \V257(7)  & \V257(6) ;
  assign n3101 = ~\V257(5)  & n3100;
  assign n3102 = \V257(5)  & ~n3100;
  assign V655 = n3101 | n3102;
  assign n3104 = \V257(7)  & ~\V257(6) ;
  assign n3105 = ~\V257(7)  & \V257(6) ;
  assign V656 = n3104 | n3105;
  assign n3107 = \V149(5)  & n2276;
  assign \V821(0)  = n2277 | n3107;
  assign n3109 = ~\V802(0)  & n550;
  assign n3110 = \V1243(9)  & ~n3109;
  assign n3111 = n2598 & n3110;
  assign n3112 = ~\V239(4)  & ~\V802(0) ;
  assign n3113 = n550 & n3112;
  assign n3114 = ~n2598 & n3113;
  assign \V1552(1)  = n3111 | n3114;
  assign n3116 = \V1243(8)  & ~n3109;
  assign n3117 = n2598 & n3116;
  assign n3118 = \V239(3)  & ~\V239(4) ;
  assign n3119 = ~\V239(3)  & \V239(4) ;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = ~\V802(0)  & ~n3120;
  assign n3122 = n550 & n3121;
  assign n3123 = ~n2598 & n3122;
  assign \V1552(0)  = n3117 | n3123;
  assign n3125 = \V70(0)  & ~n540;
  assign n3126 = V763 & n3125;
  assign n3127 = n837 & n3126;
  assign V775 = \V14(0)  & n3127;
  assign V779 = \V6(0)  & n2513;
  assign n3130 = ~\V174(0)  & n1533;
  assign n3131 = ~\V52(0)  & ~n3130;
  assign n3132 = \V12(0)  & ~n3131;
  assign V781 = \V6(0)  & n3132;
  assign V783 = \V11(0)  & \V5(0) ;
  assign V784 = \V7(0)  & \V11(0) ;
  assign V801 = n501 & n515;
  assign n3137 = \V56(0)  & ~n2974;
  assign n3138 = \V802(0)  & ~n2984;
  assign n3139 = \V56(0)  & V763;
  assign n3140 = ~n515 & n3139;
  assign n3141 = ~n3131 & n3140;
  assign n3142 = n501 & ~n515;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = ~n3138 & n3143;
  assign n3145 = ~n3137 & n3144;
  assign n3146 = n837 & ~n3145;
  assign V966 = \V14(0)  & n3146;
  assign n3148 = ~n550 & n632;
  assign n3149 = ~n1803 & n3148;
  assign n3150 = \V59(0)  & ~n3149;
  assign n3151 = \V56(0)  & n2974;
  assign n3152 = n2651 & n3151;
  assign n3153 = ~n3141 & n3152;
  assign n3154 = \V62(0)  & ~n541;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3150 & n3155;
  assign n3157 = n837 & ~n3156;
  assign V986 = \V14(0)  & n3157;
  assign \V1243(0)  = ~\V321(2) ;
  assign \V585(0)  = ~\V34(0) ;
  assign \V1833(0)  = ~\V261(0) ;
  assign \V1760(0)  = ~\V101(0) ;
  assign \V1495(0)  = ~\V175(0) ;
  assign \V1863(0)  = ~\V301(0) ;
  assign V1375 = ~\V268(5) ;
  assign \V1864(0)  = ~\V302(0) ;
  assign \V1481(0)  = ~\V214(0) ;
  assign \V1671(0)  = ~\V205(0) ;
  assign V657 = ~\V257(7) ;
endmodule


