// Benchmark "i10" written by ABC on Tue May 16 16:07:49 2017

module i10 ( 
    \V223(1) , \V223(0) , \V100(3) , \V100(2) , \V100(5) , \V100(4) ,
    \V100(1) , \V100(0) , \V60(0) , \V247(0) , \V7(0) , \V124(3) ,
    \V124(2) , \V124(5) , \V124(4) , \V11(0) , \V124(1) , \V124(0) ,
    \V259(0) , \V84(0) , \V84(1) , \V84(2) , \V84(3) , \V84(4) , \V84(5) ,
    \V35(0) , \V302(0) , \V59(0) , \V240(0) , \V203(0) , \V288(3) ,
    \V215(0) , \V288(2) , \V288(5) , \V288(4) , \V40(0) , \V288(1) ,
    \V288(0) , \V165(3) , \V165(2) , \V165(5) , \V165(4) , \V239(3) ,
    \V288(7) , \V239(2) , \V288(6) , \V52(0) , \V165(1) , \V239(4) ,
    \V165(0) , \V239(1) , \V239(0) , \V165(7) , \V165(6) , \V177(0) ,
    \V189(3) , \V189(2) , \V189(5) , \V189(4) , \V189(1) , \V189(0) ,
    \V15(0) , \V88(0) , \V88(1) , \V88(2) , \V88(3) , \V39(0) , \V293(0) ,
    \V244(0) , \V4(0) , \V194(3) , \V194(2) , \V194(4) , \V268(3) ,
    \V268(2) , \V268(5) , \V194(1) , \V268(4) , \V194(0) , \V268(1) ,
    \V268(0) , \V207(0) , \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V32(4) ,
    \V32(5) , \V32(6) , \V32(7) , \V32(8) , \V44(0) , \V32(9) , \V108(3) ,
    \V108(2) , \V56(0) , \V108(5) , \V108(4) , \V169(1) , \V169(0) ,
    \V108(1) , \V108(0) , \V68(0) , \V261(0) , \V101(0) , \V174(0) ,
    \V248(0) , \V8(0) , \V12(0) , \V149(3) , \V149(2) , \V149(5) ,
    \V149(4) , \V149(1) , \V149(0) , \V149(7) , \V149(6) , \V48(0) ,
    \V290(0) , \V32(11) , \V32(10) , \V241(0) , \V1(0) , \V204(0) ,
    \V277(0) , \V216(0) , \V41(0) , \V289(0) , \V53(0) , \V65(0) ,
    \V16(0) , \V270(0) , \V294(0) , \V171(0) , \V183(3) , \V110(0) ,
    \V183(2) , \V245(0) , \V183(5) , \V5(0) , \V183(4) , \V257(3) ,
    \V257(2) , \V70(0) , \V257(5) , \V183(1) , \V257(4) , \V183(0) ,
    \V257(1) , \V257(0) , \V257(7) , \V257(6) , \V134(1) , \V134(0) ,
    \V269(0) , \V94(0) , \V94(1) , \V33(0) , \V45(0) , \V57(0) , \V109(0) ,
    \V69(0) , \V262(0) , \V213(3) , \V213(2) , \V213(5) , \V213(4) ,
    \V274(0) , \V213(1) , \V213(0) , \V50(0) , \V102(0) , \V62(0) ,
    \V175(0) , \V249(0) , \V9(0) , \V13(0) , \V199(3) , \V199(2) ,
    \V199(4) , \V199(1) , \V199(0) , \V37(0) , \V291(0) , \V242(0) ,
    \V2(0) , \V205(0) , \V91(0) , \V91(1) , \V278(0) , \V229(3) ,
    \V229(2) , \V42(0) , \V229(5) , \V229(4) , \V229(1) , \V229(0) ,
    \V118(3) , \V118(2) , \V66(0) , \V118(5) , \V118(4) , \V118(1) ,
    \V118(0) , \V78(0) , \V78(1) , \V118(7) , \V78(2) , \V118(6) ,
    \V78(3) , \V78(4) , \V78(5) , \V271(0) , \V234(3) , \V234(2) ,
    \V234(4) , \V295(0) , \V234(1) , \V234(0) , \V172(0) , \V246(0) ,
    \V6(0) , \V71(0) , \V10(0) , \V258(0) , \V34(0) , \V46(0) , \V301(0) ,
    \V202(0) , \V275(0) , \V214(0) , \V51(0) , \V63(0) , \V14(0) ,
    \V38(0) , \V280(0) , \V292(0) , \V243(0) , \V3(0) , \V132(3) ,
    \V132(2) , \V132(5) , \V132(4) , \V132(1) , \V132(0) , \V132(7) ,
    \V132(6) , \V279(0) , \V43(0) , \V55(0) , \V67(0) , \V260(0) ,
    \V272(0) , \V223(3) , \V223(2) , \V223(5) , \V223(4) ,
    \V1243(7) , \V500(0) , \V1243(6) , \V1243(9) , \V1243(8) , \V1243(1) ,
    \V1243(0) , \V1717(0) , \V1243(3) , \V1243(2) , \V1243(5) , \V1243(4) ,
    \V585(0) , \V597(0) , \V1679(0) , \V1833(0) , \V1968(0) , \V1771(1) ,
    \V1771(0) , \V640(0) , \V375(0) , \V603(0) , \V1758(0) , \V1900(0) ,
    \V1709(1) , \V1709(0) , \V1709(3) , \V1709(2) , \V1709(4) , \V1512(1) ,
    \V1512(3) , \V1512(2) , \V1536(0) , \V1898(0) , \V1652(0) , \V1726(0) ,
    \V1953(7) , \V1953(6) , \V410(0) , \V1953(1) , \V1953(0) , \V1953(3) ,
    \V1953(2) , \V1953(5) , \V1953(4) , \V508(0) , \V1392(0) , \V1829(7) ,
    \V1829(6) , \V1829(9) , \V1829(8) , \V1281(0) , \V1620(0) , \V1829(1) ,
    \V1829(0) , \V1829(3) , \V1829(2) , \V1693(0) , \V1829(5) , \V1829(4) ,
    \V1921(1) , \V1921(0) , \V1921(3) , \V1921(2) , \V1921(5) , \V1921(4) ,
    \V802(0) , \V826(0) , \V1213(10) , \V1213(11) , \V1760(0) , \V1495(0) ,
    \V591(0) , \V1759(0) , \V1901(0) , \V1297(1) , \V1297(0) , \V1297(3) ,
    \V1297(2) , \V1297(4) , \V1451(0) , \V1863(0) , \V393(0) , \V1899(0) ,
    \V1480(0) , \V423(0) , \V1492(0) , \V435(0) , \V1781(1) , \V1781(0) ,
    V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265,
    V1266, V1267, \V1467(0) , V1365, V1370, V1371, V1372, V1373, V1374,
    V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1423, V1426, V1428,
    V1429, V1431, V1432, V1470, \V1645(0) , V1537, V1539, V1669, V1719,
    \V1896(0) , V1736, V1832, \V1459(0) , \V1213(7) , \V1213(6) ,
    \V1213(9) , \V1213(8) , \V1613(1) , \V1274(0) , \V1613(0) , \V1213(1) ,
    \V1213(0) , \V1213(3) , \V1213(2) , \V1213(5) , \V1213(4) , \V1440(0) ,
    \V321(2) , \V1864(0) , \V1741(0) , \V572(3) , \V572(2) , \V634(0) ,
    \V572(5) , \V572(4) , \V1439(0) , \V572(1) , \V572(0) , \V511(0) ,
    \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) , \V1992(0) ,
    \V609(0) , \V1481(0) , \V1629(0) , \V798(0) , \V398(0) , \V1671(0) ,
    \V1745(0) , \V1757(0) , \V1960(1) , \V1960(0) , V356, V357, V373, V377,
    \V1897(0) , V432, V512, V527, V537, V538, V539, V540, V541, V542, V543,
    V544, V545, V546, V547, V548, V587, V620, V621, V630, V650, V651, V652,
    V653, V654, V655, V656, V657, \V821(0) , \V1552(1) , \V1552(0) , V707,
    V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V801,
    V966, V986  );
  input  \V223(1) , \V223(0) , \V100(3) , \V100(2) , \V100(5) ,
    \V100(4) , \V100(1) , \V100(0) , \V60(0) , \V247(0) , \V7(0) ,
    \V124(3) , \V124(2) , \V124(5) , \V124(4) , \V11(0) , \V124(1) ,
    \V124(0) , \V259(0) , \V84(0) , \V84(1) , \V84(2) , \V84(3) , \V84(4) ,
    \V84(5) , \V35(0) , \V302(0) , \V59(0) , \V240(0) , \V203(0) ,
    \V288(3) , \V215(0) , \V288(2) , \V288(5) , \V288(4) , \V40(0) ,
    \V288(1) , \V288(0) , \V165(3) , \V165(2) , \V165(5) , \V165(4) ,
    \V239(3) , \V288(7) , \V239(2) , \V288(6) , \V52(0) , \V165(1) ,
    \V239(4) , \V165(0) , \V239(1) , \V239(0) , \V165(7) , \V165(6) ,
    \V177(0) , \V189(3) , \V189(2) , \V189(5) , \V189(4) , \V189(1) ,
    \V189(0) , \V15(0) , \V88(0) , \V88(1) , \V88(2) , \V88(3) , \V39(0) ,
    \V293(0) , \V244(0) , \V4(0) , \V194(3) , \V194(2) , \V194(4) ,
    \V268(3) , \V268(2) , \V268(5) , \V194(1) , \V268(4) , \V194(0) ,
    \V268(1) , \V268(0) , \V207(0) , \V32(0) , \V32(1) , \V32(2) ,
    \V32(3) , \V32(4) , \V32(5) , \V32(6) , \V32(7) , \V32(8) , \V44(0) ,
    \V32(9) , \V108(3) , \V108(2) , \V56(0) , \V108(5) , \V108(4) ,
    \V169(1) , \V169(0) , \V108(1) , \V108(0) , \V68(0) , \V261(0) ,
    \V101(0) , \V174(0) , \V248(0) , \V8(0) , \V12(0) , \V149(3) ,
    \V149(2) , \V149(5) , \V149(4) , \V149(1) , \V149(0) , \V149(7) ,
    \V149(6) , \V48(0) , \V290(0) , \V32(11) , \V32(10) , \V241(0) ,
    \V1(0) , \V204(0) , \V277(0) , \V216(0) , \V41(0) , \V289(0) ,
    \V53(0) , \V65(0) , \V16(0) , \V270(0) , \V294(0) , \V171(0) ,
    \V183(3) , \V110(0) , \V183(2) , \V245(0) , \V183(5) , \V5(0) ,
    \V183(4) , \V257(3) , \V257(2) , \V70(0) , \V257(5) , \V183(1) ,
    \V257(4) , \V183(0) , \V257(1) , \V257(0) , \V257(7) , \V257(6) ,
    \V134(1) , \V134(0) , \V269(0) , \V94(0) , \V94(1) , \V33(0) ,
    \V45(0) , \V57(0) , \V109(0) , \V69(0) , \V262(0) , \V213(3) ,
    \V213(2) , \V213(5) , \V213(4) , \V274(0) , \V213(1) , \V213(0) ,
    \V50(0) , \V102(0) , \V62(0) , \V175(0) , \V249(0) , \V9(0) , \V13(0) ,
    \V199(3) , \V199(2) , \V199(4) , \V199(1) , \V199(0) , \V37(0) ,
    \V291(0) , \V242(0) , \V2(0) , \V205(0) , \V91(0) , \V91(1) ,
    \V278(0) , \V229(3) , \V229(2) , \V42(0) , \V229(5) , \V229(4) ,
    \V229(1) , \V229(0) , \V118(3) , \V118(2) , \V66(0) , \V118(5) ,
    \V118(4) , \V118(1) , \V118(0) , \V78(0) , \V78(1) , \V118(7) ,
    \V78(2) , \V118(6) , \V78(3) , \V78(4) , \V78(5) , \V271(0) ,
    \V234(3) , \V234(2) , \V234(4) , \V295(0) , \V234(1) , \V234(0) ,
    \V172(0) , \V246(0) , \V6(0) , \V71(0) , \V10(0) , \V258(0) , \V34(0) ,
    \V46(0) , \V301(0) , \V202(0) , \V275(0) , \V214(0) , \V51(0) ,
    \V63(0) , \V14(0) , \V38(0) , \V280(0) , \V292(0) , \V243(0) , \V3(0) ,
    \V132(3) , \V132(2) , \V132(5) , \V132(4) , \V132(1) , \V132(0) ,
    \V132(7) , \V132(6) , \V279(0) , \V43(0) , \V55(0) , \V67(0) ,
    \V260(0) , \V272(0) , \V223(3) , \V223(2) , \V223(5) , \V223(4) ;
  output \V1243(7) , \V500(0) , \V1243(6) , \V1243(9) , \V1243(8) ,
    \V1243(1) , \V1243(0) , \V1717(0) , \V1243(3) , \V1243(2) , \V1243(5) ,
    \V1243(4) , \V585(0) , \V597(0) , \V1679(0) , \V1833(0) , \V1968(0) ,
    \V1771(1) , \V1771(0) , \V640(0) , \V375(0) , \V603(0) , \V1758(0) ,
    \V1900(0) , \V1709(1) , \V1709(0) , \V1709(3) , \V1709(2) , \V1709(4) ,
    \V1512(1) , \V1512(3) , \V1512(2) , \V1536(0) , \V1898(0) , \V1652(0) ,
    \V1726(0) , \V1953(7) , \V1953(6) , \V410(0) , \V1953(1) , \V1953(0) ,
    \V1953(3) , \V1953(2) , \V1953(5) , \V1953(4) , \V508(0) , \V1392(0) ,
    \V1829(7) , \V1829(6) , \V1829(9) , \V1829(8) , \V1281(0) , \V1620(0) ,
    \V1829(1) , \V1829(0) , \V1829(3) , \V1829(2) , \V1693(0) , \V1829(5) ,
    \V1829(4) , \V1921(1) , \V1921(0) , \V1921(3) , \V1921(2) , \V1921(5) ,
    \V1921(4) , \V802(0) , \V826(0) , \V1213(10) , \V1213(11) , \V1760(0) ,
    \V1495(0) , \V591(0) , \V1759(0) , \V1901(0) , \V1297(1) , \V1297(0) ,
    \V1297(3) , \V1297(2) , \V1297(4) , \V1451(0) , \V1863(0) , \V393(0) ,
    \V1899(0) , \V1480(0) , \V423(0) , \V1492(0) , \V435(0) , \V1781(1) ,
    \V1781(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1467(0) , V1365, V1370, V1371, V1372,
    V1373, V1374, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1423,
    V1426, V1428, V1429, V1431, V1432, V1470, \V1645(0) , V1537, V1539,
    V1669, V1719, \V1896(0) , V1736, V1832, \V1459(0) , \V1213(7) ,
    \V1213(6) , \V1213(9) , \V1213(8) , \V1613(1) , \V1274(0) , \V1613(0) ,
    \V1213(1) , \V1213(0) , \V1213(3) , \V1213(2) , \V1213(5) , \V1213(4) ,
    \V1440(0) , \V321(2) , \V1864(0) , \V1741(0) , \V572(3) , \V572(2) ,
    \V634(0) , \V572(5) , \V572(4) , \V1439(0) , \V572(1) , \V572(0) ,
    \V511(0) , \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) ,
    \V1992(0) , \V609(0) , \V1481(0) , \V1629(0) , \V798(0) , \V398(0) ,
    \V1671(0) , \V1745(0) , \V1757(0) , \V1960(1) , \V1960(0) , V356, V357,
    V373, V377, \V1897(0) , V432, V512, V527, V537, V538, V539, V540, V541,
    V542, V543, V544, V545, V546, V547, V548, V587, V620, V621, V630, V650,
    V651, V652, V653, V654, V655, V656, V657, \V821(0) , \V1552(1) ,
    \V1552(0) , V707, V763, V775, V778, V779, V780, V781, V782, V783, V784,
    V787, V789, V801, V966, V986;
  wire n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n830, n831, n832, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n922, n923, n924, n925, n926, n927, n929,
    n930, n931, n932, n933, n935, n936, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n953, n954, n956, n957,
    n959, n960, n964, n972, n973, n974, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n986, n987, n988, n989, n990, n992, n993, n994, n995,
    n996, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1011, n1012, n1013, n1014, n1016, n1017, n1018,
    n1019, n1021, n1022, n1023, n1024, n1026, n1027, n1028, n1029, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1621, n1622, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1658, n1659, n1660, n1661, n1662, n1663,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1674, n1676,
    n1677, n1679, n1680, n1681, n1682, n1683, n1684, n1686, n1687, n1688,
    n1689, n1690, n1691, n1693, n1694, n1695, n1696, n1697, n1698, n1700,
    n1701, n1702, n1703, n1704, n1705, n1707, n1708, n1709, n1710, n1711,
    n1712, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1831, n1832, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1856, n1857,
    n1859, n1860, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1885, n1886, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1917, n1918, n1919, n1920, n1921, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1938, n1939, n1941, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1963, n1964, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1986, n1987, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2020, n2021, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2045, n2046, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2165, n2166, n2167, n2168, n2170, n2171, n2172, n2173,
    n2174, n2175, n2177, n2179, n2180, n2181, n2182, n2184, n2185, n2186,
    n2187, n2189, n2190, n2191, n2192, n2194, n2195, n2196, n2197, n2199,
    n2200, n2201, n2202, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2269, n2270, n2272, n2273,
    n2274, n2275, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2378, n2379,
    n2381, n2382, n2384, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2427, n2428, n2430, n2431, n2432, n2433,
    n2435, n2436, n2437, n2439, n2440, n2441, n2443, n2444, n2446, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2470,
    n2471, n2473, n2474, n2475, n2476, n2482, n2484, n2485, n2487, n2488,
    n2490, n2492, n2493, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2540, n2541, n2543, n2544,
    n2545, n2547, n2548, n2549, n2550, n2552, n2553, n2554, n2555, n2556,
    n2558, n2559, n2560, n2561, n2563, n2564, n2565, n2566, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2671, n2672, n2673, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2701, n2702, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2740, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2804, n2805, n2806, n2807, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2866, n2867, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2887, n2889, n2890, n2892, n2893, n2894, n2895, n2896, n2897, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2947, n2948, n2949, n2950, n2951, n2953, n2954, n2955, n2956, n2958,
    n2959, n2960, n2961, n2963, n2964, n2965, n2967, n2968, n2969, n2971,
    n2972, n2974, n2976, n2977, n2978, n2979, n2980, n2981, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2991, n2992, n2993, n2996, n2997,
    n2998, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021;
  assign n482 = ~\V149(4)  & ~\V149(0) ;
  assign n483 = \V149(1)  & n482;
  assign n484 = \V149(2)  & n483;
  assign n485 = ~\V149(3)  & n484;
  assign n486 = \V149(1)  & ~\V149(0) ;
  assign n487 = \V149(2)  & n486;
  assign n488 = \V149(3)  & n487;
  assign n489 = \V165(2)  & \V165(0) ;
  assign n490 = \V165(4)  & n489;
  assign n491 = \V165(5)  & n490;
  assign n492 = \V165(6)  & n491;
  assign n493 = \V165(7)  & n492;
  assign n494 = \V165(1)  & n493;
  assign n495 = \V165(3)  & n494;
  assign n496 = ~\V204(0)  & n495;
  assign n497 = \V261(0)  & n496;
  assign n498 = ~\V165(4)  & \V70(0) ;
  assign n499 = ~\V165(5)  & n498;
  assign n500 = ~\V165(6)  & n499;
  assign n501 = \V165(3)  & n500;
  assign n502 = ~\V149(2)  & n486;
  assign n503 = ~\V149(7)  & \V149(6) ;
  assign n504 = \V149(5)  & n503;
  assign n505 = \V149(4)  & n504;
  assign n506 = ~\V149(3)  & n505;
  assign n507 = n502 & n506;
  assign n508 = \V149(7)  & \V149(6) ;
  assign n509 = \V149(5)  & n508;
  assign n510 = \V149(4)  & n509;
  assign n511 = ~\V149(3)  & n510;
  assign n512 = n502 & n511;
  assign n513 = ~n507 & ~n512;
  assign \V802(0)  = \V52(0)  | \V51(0) ;
  assign n515 = ~\V55(0)  & ~\V802(0) ;
  assign n516 = ~n513 & n515;
  assign n517 = ~\V149(1)  & ~\V149(0) ;
  assign n518 = ~\V149(2)  & n517;
  assign n519 = \V149(4)  & ~\V149(0) ;
  assign n520 = \V149(1)  & n519;
  assign n521 = \V149(2)  & n520;
  assign n522 = ~\V149(3)  & n521;
  assign n523 = ~n518 & ~n522;
  assign n524 = ~n516 & n523;
  assign n525 = \V169(0)  & ~\V292(0) ;
  assign n526 = ~\V291(0)  & n525;
  assign n527 = ~n524 & n526;
  assign V763 = ~n501 & n527;
  assign n529 = \V165(7)  & \V70(0) ;
  assign n530 = \V261(0)  & n529;
  assign n531 = \V165(5)  & n530;
  assign n532 = \V165(3)  & n531;
  assign n533 = \V165(4)  & n532;
  assign n534 = \V165(6)  & n533;
  assign n535 = \V165(0)  & n534;
  assign n536 = \V165(1)  & n535;
  assign n537 = \V165(2)  & n536;
  assign n538 = V763 & n537;
  assign n539 = ~n497 & ~n538;
  assign n540 = ~\V262(0)  & n539;
  assign n541 = ~\V56(0)  & \V53(0) ;
  assign n542 = n540 & n541;
  assign n543 = ~n488 & n542;
  assign n544 = ~n485 & n543;
  assign n545 = \V149(2)  & n517;
  assign n546 = ~n518 & ~n545;
  assign n547 = \V169(1)  & ~n546;
  assign n548 = ~\V174(0)  & n518;
  assign n549 = \V149(5)  & ~\V149(4) ;
  assign n550 = ~\V149(3)  & n549;
  assign n551 = ~\V88(2)  & n550;
  assign n552 = \V88(3)  & n551;
  assign n553 = n548 & n552;
  assign V707 = ~\V149(3)  & n548;
  assign n555 = ~\V149(5)  & ~\V149(4) ;
  assign n556 = \V88(2)  & n555;
  assign n557 = \V88(3)  & n556;
  assign n558 = V707 & n557;
  assign n559 = ~\V88(2)  & n555;
  assign n560 = \V88(3)  & n559;
  assign n561 = V707 & n560;
  assign n562 = ~\V149(5)  & \V149(4) ;
  assign n563 = V707 & n562;
  assign n564 = \V149(5)  & V707;
  assign n565 = \V149(4)  & n564;
  assign n566 = ~\V88(3)  & n556;
  assign n567 = V707 & n566;
  assign n568 = ~\V88(3)  & n551;
  assign n569 = n548 & n568;
  assign n570 = \V88(2)  & n550;
  assign n571 = ~\V88(3)  & n570;
  assign n572 = n548 & n571;
  assign n573 = ~n569 & ~n572;
  assign n574 = ~n567 & n573;
  assign n575 = ~n565 & n574;
  assign n576 = ~n563 & n575;
  assign n577 = ~n561 & n576;
  assign n578 = ~n558 & n577;
  assign n579 = ~n553 & n578;
  assign n580 = n547 & ~n579;
  assign n581 = \V56(0)  & n580;
  assign n582 = \V149(3)  & n548;
  assign n583 = n547 & n582;
  assign n584 = \V56(0)  & n583;
  assign n585 = \V60(0)  & n583;
  assign n586 = \V60(0)  & n580;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n584 & n587;
  assign n589 = ~n581 & n588;
  assign n590 = ~\V56(0)  & ~\V53(0) ;
  assign n591 = ~\V57(0)  & n590;
  assign n592 = \V149(3)  & n545;
  assign n593 = n545 & n550;
  assign n594 = ~\V149(3)  & n555;
  assign n595 = n545 & n594;
  assign n596 = ~\V149(3)  & n562;
  assign n597 = n545 & n596;
  assign n598 = ~n595 & ~n597;
  assign n599 = ~n593 & n598;
  assign n600 = ~\V174(0)  & n522;
  assign n601 = \V277(0)  & n600;
  assign n602 = \V278(0)  & ~n601;
  assign n603 = n600 & ~n602;
  assign n604 = n599 & ~n603;
  assign n605 = ~n582 & n604;
  assign n606 = n579 & n605;
  assign n607 = ~n592 & n606;
  assign n608 = ~n591 & ~n607;
  assign n609 = n589 & n608;
  assign n610 = ~\V149(5)  & n508;
  assign n611 = \V149(4)  & n610;
  assign n612 = ~\V149(3)  & n611;
  assign n613 = n502 & n612;
  assign n614 = ~n609 & ~n613;
  assign n615 = ~n544 & n614;
  assign n616 = ~n592 & ~n600;
  assign n617 = \V60(0)  & ~n616;
  assign n618 = ~n615 & ~n617;
  assign n619 = \V84(5)  & n618;
  assign n620 = ~n615 & n619;
  assign n621 = ~\V59(0)  & ~\V56(0) ;
  assign n622 = ~\V60(0)  & n621;
  assign n623 = V763 & ~n622;
  assign n624 = V763 & n540;
  assign n625 = \V32(9)  & n624;
  assign n626 = n623 & n625;
  assign n627 = ~\V59(0)  & n488;
  assign n628 = ~n602 & n627;
  assign n629 = ~\V60(0)  & ~\V59(0) ;
  assign n630 = n488 & ~n602;
  assign n631 = ~n629 & n630;
  assign n632 = n488 & n602;
  assign n633 = n546 & ~n600;
  assign n634 = ~n485 & n633;
  assign n635 = ~\V174(0)  & ~n634;
  assign n636 = ~n632 & ~n635;
  assign n637 = ~n631 & n636;
  assign n638 = ~n488 & ~n600;
  assign n639 = ~n485 & n638;
  assign n640 = \V199(2)  & ~n639;
  assign n641 = n546 & n640;
  assign n642 = \V239(2)  & n639;
  assign n643 = ~n546 & n642;
  assign n644 = ~n641 & ~n643;
  assign n645 = n540 & ~n644;
  assign n646 = ~n637 & n645;
  assign n647 = ~n628 & n646;
  assign n648 = ~n624 & n647;
  assign n649 = ~n626 & ~n648;
  assign n650 = ~n618 & ~n649;
  assign n651 = n615 & n650;
  assign \V1243(7)  = n620 | n651;
  assign \V500(0)  = \V271(0)  | ~\V14(0) ;
  assign n654 = \V84(4)  & n618;
  assign n655 = ~n615 & n654;
  assign n656 = \V32(11)  & ~n623;
  assign n657 = \V32(8)  & n623;
  assign n658 = ~n656 & ~n657;
  assign n659 = n624 & ~n658;
  assign n660 = \V199(1)  & ~n639;
  assign n661 = n546 & n660;
  assign n662 = \V239(1)  & n639;
  assign n663 = ~n546 & n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = n540 & ~n664;
  assign n666 = ~n637 & n665;
  assign n667 = ~n628 & n666;
  assign n668 = ~n624 & n667;
  assign n669 = ~n659 & ~n668;
  assign n670 = ~n618 & ~n669;
  assign n671 = n615 & n670;
  assign \V1243(6)  = n655 | n671;
  assign n673 = \V88(1)  & n618;
  assign n674 = ~n615 & n673;
  assign n675 = \V32(11)  & n624;
  assign n676 = n623 & n675;
  assign n677 = \V199(4)  & ~n639;
  assign n678 = n546 & n677;
  assign n679 = \V239(4)  & n639;
  assign n680 = ~n546 & n679;
  assign n681 = ~n678 & ~n680;
  assign n682 = n540 & ~n681;
  assign n683 = ~n637 & n682;
  assign n684 = ~n628 & n683;
  assign n685 = ~n624 & n684;
  assign n686 = ~n676 & ~n685;
  assign n687 = ~n618 & ~n686;
  assign n688 = n615 & n687;
  assign \V1243(9)  = n674 | n688;
  assign n690 = \V88(0)  & n618;
  assign n691 = ~n615 & n690;
  assign n692 = \V32(10)  & n624;
  assign n693 = n623 & n692;
  assign n694 = \V199(3)  & ~n639;
  assign n695 = n546 & n694;
  assign n696 = \V239(3)  & n639;
  assign n697 = ~n546 & n696;
  assign n698 = ~n695 & ~n697;
  assign n699 = n540 & ~n698;
  assign n700 = ~n637 & n699;
  assign n701 = ~n628 & n700;
  assign n702 = ~n624 & n701;
  assign n703 = ~n693 & ~n702;
  assign n704 = ~n618 & ~n703;
  assign n705 = n615 & n704;
  assign \V1243(8)  = n691 | n705;
  assign n707 = \V78(5)  & n618;
  assign n708 = ~n615 & n707;
  assign n709 = \V32(6)  & ~n623;
  assign n710 = \V32(3)  & n623;
  assign n711 = ~n709 & ~n710;
  assign n712 = n624 & ~n711;
  assign n713 = ~\V59(0)  & \V149(5) ;
  assign n714 = n540 & n713;
  assign n715 = n488 & n714;
  assign n716 = ~n602 & n715;
  assign n717 = n637 & n716;
  assign n718 = \V194(1)  & ~n639;
  assign n719 = n546 & n718;
  assign n720 = \V234(1)  & n639;
  assign n721 = ~n546 & n720;
  assign n722 = ~n719 & ~n721;
  assign n723 = n540 & ~n722;
  assign n724 = ~n637 & n723;
  assign n725 = ~n628 & n724;
  assign n726 = ~n717 & ~n725;
  assign n727 = ~n624 & ~n726;
  assign n728 = ~n712 & ~n727;
  assign n729 = ~n618 & ~n728;
  assign n730 = n615 & n729;
  assign \V1243(1)  = n708 | n730;
  assign n732 = \V78(4)  & n618;
  assign n733 = ~n615 & n732;
  assign n734 = \V32(5)  & ~n623;
  assign n735 = \V32(2)  & n623;
  assign n736 = ~n734 & ~n735;
  assign n737 = n624 & ~n736;
  assign n738 = \V194(0)  & ~n639;
  assign n739 = n546 & n738;
  assign n740 = \V234(0)  & n639;
  assign n741 = ~n546 & n740;
  assign n742 = ~n739 & ~n741;
  assign n743 = n540 & ~n742;
  assign n744 = ~n637 & n743;
  assign n745 = ~n628 & n744;
  assign n746 = ~\V59(0)  & \V149(4) ;
  assign n747 = n540 & n746;
  assign n748 = n488 & n747;
  assign n749 = ~n602 & n748;
  assign n750 = n637 & n749;
  assign n751 = \V257(7)  & ~n540;
  assign n752 = n637 & n751;
  assign n753 = ~n628 & n752;
  assign n754 = ~n750 & ~n753;
  assign n755 = ~n745 & n754;
  assign n756 = ~n624 & ~n755;
  assign n757 = ~n737 & ~n756;
  assign n758 = ~n618 & ~n757;
  assign n759 = n615 & n758;
  assign \V321(2)  = ~n733 & ~n759;
  assign n761 = ~n602 & ~n639;
  assign n762 = ~n592 & ~n761;
  assign n763 = \V802(0)  & ~n762;
  assign n764 = ~\V280(0)  & n592;
  assign n765 = \V242(0)  & ~\V275(0) ;
  assign n766 = \V134(1)  & n765;
  assign n767 = \V134(0)  & n766;
  assign n768 = \V272(0)  & n767;
  assign n769 = ~\V802(0)  & n768;
  assign n770 = n602 & n769;
  assign n771 = \V241(0)  & ~n638;
  assign n772 = ~n485 & ~n771;
  assign n773 = \V261(0)  & ~\V802(0) ;
  assign n774 = ~n602 & n773;
  assign n775 = ~n772 & n774;
  assign n776 = \V56(0)  & ~n638;
  assign n777 = \V242(0)  & ~\V802(0) ;
  assign n778 = ~n639 & n777;
  assign n779 = ~n602 & n778;
  assign n780 = ~n776 & n779;
  assign n781 = ~\V174(0)  & n512;
  assign n782 = \V56(0)  & \V172(0) ;
  assign n783 = \V207(0)  & ~n782;
  assign n784 = \V59(0)  & ~n545;
  assign n785 = n783 & n784;
  assign n786 = n781 & n785;
  assign n787 = ~\V149(7)  & ~\V149(6) ;
  assign n788 = \V149(5)  & n787;
  assign n789 = ~\V149(4)  & n788;
  assign n790 = ~\V149(3)  & n789;
  assign n791 = n502 & n790;
  assign n792 = ~n545 & ~n547;
  assign n793 = n783 & n792;
  assign n794 = ~n791 & n793;
  assign n795 = ~n781 & n794;
  assign n796 = \V172(0)  & \V67(0) ;
  assign n797 = \V215(0)  & n796;
  assign n798 = n547 & n784;
  assign n799 = n783 & n798;
  assign n800 = \V62(0)  & ~n545;
  assign n801 = n783 & n800;
  assign n802 = n791 & n801;
  assign n803 = ~n799 & ~n802;
  assign n804 = ~\V214(0)  & n803;
  assign n805 = ~n797 & n804;
  assign n806 = ~n795 & n805;
  assign n807 = ~n786 & n806;
  assign n808 = \V261(0)  & ~\V275(0) ;
  assign n809 = \V272(0)  & n808;
  assign n810 = ~\V802(0)  & n809;
  assign n811 = n602 & n810;
  assign n812 = ~n772 & n811;
  assign n813 = n807 & ~n812;
  assign n814 = ~n780 & n813;
  assign n815 = ~n775 & n814;
  assign n816 = ~n770 & n815;
  assign n817 = ~\V165(2)  & \V165(0) ;
  assign n818 = \V165(1)  & n817;
  assign n819 = ~\V165(7)  & n818;
  assign n820 = \V165(7)  & ~\V290(0) ;
  assign n821 = n818 & n820;
  assign n822 = ~\V302(0)  & ~n821;
  assign n823 = ~n819 & n822;
  assign n824 = n816 & n823;
  assign n825 = \V203(0)  & ~\V165(0) ;
  assign n826 = \V165(2)  & n825;
  assign n827 = \V165(1)  & n826;
  assign n828 = \V240(0)  & ~\V172(0) ;
  assign V1719 = ~n818 & n828;
  assign n830 = ~n827 & V1719;
  assign n831 = n824 & n830;
  assign n832 = ~n764 & n831;
  assign \V1717(0)  = n763 | n832;
  assign n834 = \V84(1)  & n618;
  assign n835 = ~n615 & n834;
  assign n836 = \V32(8)  & ~n623;
  assign n837 = \V32(5)  & n623;
  assign n838 = ~n836 & ~n837;
  assign n839 = n624 & ~n838;
  assign n840 = ~\V59(0)  & \V149(7) ;
  assign n841 = n540 & n840;
  assign n842 = n488 & n841;
  assign n843 = ~n602 & n842;
  assign n844 = n637 & n843;
  assign n845 = \V194(3)  & ~n639;
  assign n846 = n546 & n845;
  assign n847 = \V234(3)  & n639;
  assign n848 = ~n546 & n847;
  assign n849 = ~n846 & ~n848;
  assign n850 = n540 & ~n849;
  assign n851 = ~n637 & n850;
  assign n852 = ~n628 & n851;
  assign n853 = ~n844 & ~n852;
  assign n854 = ~n624 & ~n853;
  assign n855 = ~n839 & ~n854;
  assign n856 = ~n618 & ~n855;
  assign n857 = n615 & n856;
  assign \V1243(3)  = n835 | n857;
  assign n859 = \V84(0)  & n618;
  assign n860 = ~n615 & n859;
  assign n861 = \V32(7)  & ~n623;
  assign n862 = \V32(4)  & n623;
  assign n863 = ~n861 & ~n862;
  assign n864 = n624 & ~n863;
  assign n865 = ~\V59(0)  & \V149(6) ;
  assign n866 = n540 & n865;
  assign n867 = n488 & n866;
  assign n868 = ~n602 & n867;
  assign n869 = n637 & n868;
  assign n870 = \V194(2)  & ~n639;
  assign n871 = n546 & n870;
  assign n872 = \V234(2)  & n639;
  assign n873 = ~n546 & n872;
  assign n874 = ~n871 & ~n873;
  assign n875 = n540 & ~n874;
  assign n876 = ~n637 & n875;
  assign n877 = ~n628 & n876;
  assign n878 = ~n869 & ~n877;
  assign n879 = ~n624 & ~n878;
  assign n880 = ~n864 & ~n879;
  assign n881 = ~n618 & ~n880;
  assign n882 = n615 & n881;
  assign \V1243(2)  = n860 | n882;
  assign n884 = \V84(3)  & n618;
  assign n885 = ~n615 & n884;
  assign n886 = \V32(10)  & ~n623;
  assign n887 = \V32(7)  & n623;
  assign n888 = ~n886 & ~n887;
  assign n889 = n624 & ~n888;
  assign n890 = \V199(0)  & ~n639;
  assign n891 = n546 & n890;
  assign n892 = \V239(0)  & n639;
  assign n893 = ~n546 & n892;
  assign n894 = ~n891 & ~n893;
  assign n895 = n540 & ~n894;
  assign n896 = ~n637 & n895;
  assign n897 = ~n628 & n896;
  assign n898 = ~n624 & n897;
  assign n899 = ~n889 & ~n898;
  assign n900 = ~n618 & ~n899;
  assign n901 = n615 & n900;
  assign \V1243(5)  = n885 | n901;
  assign n903 = \V84(2)  & n618;
  assign n904 = ~n615 & n903;
  assign n905 = \V32(9)  & ~n623;
  assign n906 = \V32(6)  & n623;
  assign n907 = ~n905 & ~n906;
  assign n908 = n624 & ~n907;
  assign n909 = \V194(4)  & ~n639;
  assign n910 = n546 & n909;
  assign n911 = \V234(4)  & n639;
  assign n912 = ~n546 & n911;
  assign n913 = ~n910 & ~n912;
  assign n914 = n540 & ~n913;
  assign n915 = ~n637 & n914;
  assign n916 = ~n628 & n915;
  assign n917 = ~n624 & n916;
  assign n918 = ~n908 & ~n917;
  assign n919 = ~n618 & ~n918;
  assign n920 = n615 & n919;
  assign \V1243(4)  = n904 | n920;
  assign n922 = \V244(0)  & \V243(0) ;
  assign n923 = \V802(0)  & ~n639;
  assign n924 = ~\V245(0)  & ~n923;
  assign n925 = n922 & n924;
  assign n926 = \V245(0)  & ~n923;
  assign n927 = ~n922 & n926;
  assign \V597(0)  = n925 | n927;
  assign n929 = ~\V59(0)  & \V258(0) ;
  assign n930 = ~\V259(0)  & n929;
  assign n931 = ~\V260(0)  & n930;
  assign n932 = \V262(0)  & \V14(0) ;
  assign n933 = ~n931 & n932;
  assign \V1679(0)  = ~n539 | n933;
  assign n935 = \V15(0)  & ~\V16(0) ;
  assign n936 = ~\V15(0)  & \V16(0) ;
  assign \V1758(0)  = n935 | n936;
  assign n938 = ~\V102(0)  & ~\V1758(0) ;
  assign n939 = ~\V110(0)  & n518;
  assign n940 = ~n938 & n939;
  assign n941 = ~\V108(4)  & \V101(0) ;
  assign n942 = n935 & n941;
  assign n943 = \V149(7)  & ~\V149(6) ;
  assign n944 = ~\V149(5)  & n943;
  assign n945 = \V149(4)  & n944;
  assign n946 = ~\V149(3)  & n945;
  assign n947 = n502 & n946;
  assign n948 = \V56(0)  & n947;
  assign n949 = \V110(0)  & \V14(0) ;
  assign n950 = ~n948 & n949;
  assign n951 = ~n942 & n950;
  assign \V1968(0)  = n940 | n951;
  assign n953 = ~\V134(1)  & ~n613;
  assign n954 = ~\V88(3)  & n613;
  assign \V1771(1)  = n953 | n954;
  assign n956 = ~\V134(0)  & ~n613;
  assign n957 = ~\V88(2)  & n613;
  assign \V1771(0)  = n956 | n957;
  assign n959 = \V274(0)  & ~\V271(0) ;
  assign n960 = ~\V202(0)  & n959;
  assign \V640(0)  = \V271(0)  | n960;
  assign V1423 = \V1(0)  & \V9(0) ;
  assign V1258 = \V9(0)  & \V2(0) ;
  assign n964 = \V109(0)  & ~\V13(0) ;
  assign V1431 = V1423 & ~n964;
  assign V787 = \V7(0)  & \V9(0) ;
  assign V778 = \V5(0)  & \V9(0) ;
  assign V780 = \V9(0)  & \V6(0) ;
  assign V1387 = \V8(0)  & \V9(0) ;
  assign V1259 = \V9(0)  & \V3(0) ;
  assign V1263 = \V4(0)  & \V9(0) ;
  assign n972 = \V71(0)  & \V202(0) ;
  assign n973 = ~\V13(0)  & n972;
  assign n974 = \V9(0)  & ~n973;
  assign V789 = \V4(0)  & n974;
  assign n976 = ~V1263 & ~V789;
  assign n977 = ~V1259 & n976;
  assign n978 = ~V1387 & n977;
  assign n979 = ~V780 & n978;
  assign n980 = ~V778 & n979;
  assign n981 = ~V787 & n980;
  assign n982 = ~V1431 & n981;
  assign n983 = ~V1258 & n982;
  assign n984 = ~V1423 & n983;
  assign \V375(0)  = V1423 | ~n984;
  assign n986 = \V245(0)  & n922;
  assign n987 = ~\V246(0)  & ~n923;
  assign n988 = n986 & n987;
  assign n989 = \V246(0)  & ~n923;
  assign n990 = ~n986 & n989;
  assign \V603(0)  = n988 | n990;
  assign n992 = ~\V149(4)  & n944;
  assign n993 = \V149(3)  & n992;
  assign n994 = n502 & n993;
  assign n995 = \V56(0)  & n994;
  assign n996 = \V108(4)  & ~n995;
  assign \V1900(0)  = n935 | n996;
  assign n998 = ~n502 & ~n518;
  assign n999 = n818 & ~n998;
  assign n1000 = \V290(0)  & n999;
  assign n1001 = \V165(4)  & n1000;
  assign n1002 = ~\V149(5)  & n503;
  assign n1003 = ~\V149(4)  & n1002;
  assign n1004 = ~\V149(3)  & n1003;
  assign n1005 = n502 & n1004;
  assign n1006 = \V56(0)  & n1005;
  assign n1007 = \V100(2)  & \V14(0) ;
  assign n1008 = ~n1006 & n1007;
  assign n1009 = ~n1000 & n1008;
  assign \V1709(1)  = n1001 | n1009;
  assign n1011 = \V165(3)  & n1000;
  assign n1012 = \V100(1)  & \V14(0) ;
  assign n1013 = ~n1006 & n1012;
  assign n1014 = ~n1000 & n1013;
  assign \V1709(0)  = n1011 | n1014;
  assign n1016 = \V165(6)  & n1000;
  assign n1017 = \V100(4)  & \V14(0) ;
  assign n1018 = ~n1006 & n1017;
  assign n1019 = ~n1000 & n1018;
  assign \V1709(3)  = n1016 | n1019;
  assign n1021 = \V165(5)  & n1000;
  assign n1022 = \V100(3)  & \V14(0) ;
  assign n1023 = ~n1006 & n1022;
  assign n1024 = ~n1000 & n1023;
  assign \V1709(2)  = n1021 | n1024;
  assign n1026 = \V165(7)  & n1000;
  assign n1027 = \V100(5)  & \V14(0) ;
  assign n1028 = ~n1006 & n1027;
  assign n1029 = ~n1000 & n1028;
  assign \V1709(4)  = n1026 | n1029;
  assign n1031 = ~\V88(3)  & n559;
  assign n1032 = V707 & n1031;
  assign n1033 = \V88(3)  & n570;
  assign n1034 = n548 & n1033;
  assign n1035 = ~n1032 & ~n1034;
  assign n1036 = n547 & ~n1035;
  assign n1037 = \V59(0)  & n1036;
  assign n1038 = ~n547 & ~n1035;
  assign n1039 = \V149(5)  & \V149(4) ;
  assign n1040 = ~\V149(3)  & n1039;
  assign n1041 = n545 & n1040;
  assign n1042 = ~n1038 & ~n1041;
  assign n1043 = \V56(0)  & ~n1042;
  assign n1044 = ~\V172(0)  & n1043;
  assign n1045 = \V56(0)  & ~n546;
  assign n1046 = \V171(0)  & n1045;
  assign n1047 = \V278(0)  & ~n639;
  assign n1048 = \V177(0)  & ~\V248(0) ;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = ~n782 & n1049;
  assign n1051 = ~n1046 & n1050;
  assign n1052 = ~\V274(0)  & ~\V271(0) ;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n1044 & n1053;
  assign n1055 = ~n1037 & n1054;
  assign n1056 = \V56(0)  & n545;
  assign n1057 = \V149(7)  & n1056;
  assign n1058 = n545 & n783;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = n816 & n1059;
  assign \V1536(0)  = n1055 | ~n1060;
  assign n1062 = \V32(3)  & n618;
  assign n1063 = ~n615 & n1062;
  assign n1064 = \V183(3)  & ~n639;
  assign n1065 = n546 & n1064;
  assign n1066 = \V223(3)  & n639;
  assign n1067 = ~n546 & n1066;
  assign n1068 = ~n1065 & ~n1067;
  assign n1069 = n540 & ~n1068;
  assign n1070 = ~n628 & n1069;
  assign n1071 = ~n637 & n1070;
  assign n1072 = ~n624 & n1071;
  assign n1073 = ~n618 & n1072;
  assign n1074 = n615 & n1073;
  assign \V1213(3)  = n1063 | n1074;
  assign n1076 = \V288(7)  & ~\V288(6) ;
  assign n1077 = \V288(5)  & ~\V288(4) ;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n1076 & n1077;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = \V288(3)  & ~\V288(2) ;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n1080 & n1081;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = \V288(1)  & ~\V288(0) ;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = n1084 & n1085;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = \V1213(3)  & n1088;
  assign n1090 = ~\V1213(3)  & ~n1088;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = \V32(2)  & n618;
  assign n1093 = ~n615 & n1092;
  assign n1094 = \V183(2)  & ~n639;
  assign n1095 = n546 & n1094;
  assign n1096 = \V223(2)  & n639;
  assign n1097 = ~n546 & n1096;
  assign n1098 = ~n1095 & ~n1097;
  assign n1099 = n540 & ~n1098;
  assign n1100 = ~n628 & n1099;
  assign n1101 = ~n637 & n1100;
  assign n1102 = ~n624 & n1101;
  assign n1103 = ~n618 & n1102;
  assign n1104 = n615 & n1103;
  assign \V1213(2)  = n1093 | n1104;
  assign n1106 = ~\V288(7)  & \V288(6) ;
  assign n1107 = ~n1076 & ~n1106;
  assign n1108 = ~\V288(5)  & \V288(4) ;
  assign n1109 = n1107 & ~n1108;
  assign n1110 = ~n1107 & n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1076 & n1077;
  assign n1113 = n1111 & n1112;
  assign n1114 = ~n1111 & ~n1112;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~\V288(3)  & \V288(2) ;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = n1115 & n1116;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1080 & n1081;
  assign n1121 = n1119 & n1120;
  assign n1122 = ~n1119 & ~n1120;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~\V288(1)  & \V288(0) ;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = n1123 & n1124;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1084 & n1085;
  assign n1129 = n1127 & n1128;
  assign n1130 = ~n1127 & ~n1128;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = \V1213(2)  & n1131;
  assign n1133 = ~\V1213(2)  & ~n1131;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = \V32(1)  & n618;
  assign n1136 = ~n615 & n1135;
  assign n1137 = \V183(1)  & ~n639;
  assign n1138 = n546 & n1137;
  assign n1139 = \V223(1)  & n639;
  assign n1140 = ~n546 & n1139;
  assign n1141 = ~n1138 & ~n1140;
  assign n1142 = n540 & ~n1141;
  assign n1143 = ~n628 & n1142;
  assign n1144 = ~n637 & n1143;
  assign n1145 = ~n624 & n1144;
  assign n1146 = ~n618 & n1145;
  assign n1147 = n615 & n1146;
  assign \V1213(1)  = n1136 | n1147;
  assign n1149 = ~\V288(7)  & ~\V288(6) ;
  assign n1150 = \V288(5)  & \V288(4) ;
  assign n1151 = n1149 & ~n1150;
  assign n1152 = ~n1149 & n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1107 & n1112;
  assign n1155 = n1108 & n1112;
  assign n1156 = n1107 & n1108;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1154 & n1157;
  assign n1159 = ~n1153 & n1158;
  assign n1160 = n1153 & ~n1158;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = \V288(3)  & \V288(2) ;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = n1161 & n1162;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1115 & n1120;
  assign n1167 = n1116 & n1120;
  assign n1168 = ~n1115 & n1116;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~n1166 & n1169;
  assign n1171 = ~n1165 & n1170;
  assign n1172 = n1165 & ~n1170;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = \V288(1)  & \V288(0) ;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n1173 & n1174;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = ~n1123 & n1128;
  assign n1179 = n1124 & n1128;
  assign n1180 = ~n1123 & n1124;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1178 & n1181;
  assign n1183 = ~n1177 & n1182;
  assign n1184 = n1177 & ~n1182;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = \V1213(1)  & n1185;
  assign n1187 = ~\V1213(1)  & ~n1185;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = \V32(0)  & n618;
  assign n1190 = ~n615 & n1189;
  assign n1191 = \V183(0)  & ~n639;
  assign n1192 = n546 & n1191;
  assign n1193 = \V223(0)  & n639;
  assign n1194 = ~n546 & n1193;
  assign n1195 = ~n1192 & ~n1194;
  assign n1196 = n540 & ~n1195;
  assign n1197 = ~n628 & n1196;
  assign n1198 = ~n637 & n1197;
  assign n1199 = ~n624 & n1198;
  assign n1200 = ~n618 & n1199;
  assign n1201 = n615 & n1200;
  assign \V1213(0)  = n1190 | n1201;
  assign n1203 = n1149 & ~n1158;
  assign n1204 = n1150 & ~n1158;
  assign n1205 = n1149 & n1150;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n1203 & n1206;
  assign n1208 = ~n1149 & ~n1207;
  assign n1209 = n1149 & n1207;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~n1161 & ~n1170;
  assign n1212 = n1162 & ~n1170;
  assign n1213 = ~n1161 & n1162;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1211 & n1214;
  assign n1216 = n1210 & ~n1215;
  assign n1217 = ~n1210 & n1215;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1173 & ~n1182;
  assign n1220 = n1174 & ~n1182;
  assign n1221 = ~n1173 & n1174;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1219 & n1222;
  assign n1224 = n1218 & ~n1223;
  assign n1225 = ~n1218 & n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = \V1213(0)  & n1226;
  assign n1228 = ~\V1213(0)  & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~\V149(5)  & n787;
  assign n1231 = ~\V149(4)  & n1230;
  assign n1232 = \V149(3)  & n1231;
  assign n1233 = n502 & n1232;
  assign n1234 = ~\V802(0)  & n1233;
  assign n1235 = n1174 & ~n1234;
  assign n1236 = n1229 & n1235;
  assign n1237 = n1188 & n1236;
  assign n1238 = n1134 & n1237;
  assign n1239 = n1091 & n1238;
  assign n1240 = \V1213(3)  & ~n1088;
  assign n1241 = ~\V1213(3)  & n1088;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = n1088 & n1131;
  assign n1244 = ~n1088 & ~n1131;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = \V1213(2)  & n1245;
  assign n1247 = ~\V1213(2)  & ~n1245;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = n1185 & n1243;
  assign n1250 = ~n1185 & ~n1243;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = \V1213(1)  & n1251;
  assign n1253 = ~\V1213(1)  & ~n1251;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = n1226 & n1249;
  assign n1256 = ~n1226 & ~n1249;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = \V1213(0)  & n1257;
  assign n1259 = ~\V1213(0)  & ~n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n1235 & n1260;
  assign n1262 = n1254 & n1261;
  assign n1263 = n1248 & n1262;
  assign n1264 = n1242 & n1263;
  assign n1265 = ~n1088 & ~n1124;
  assign n1266 = ~n1088 & n1124;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = \V1213(3)  & n1267;
  assign n1269 = ~\V1213(3)  & ~n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1088 & n1245;
  assign n1272 = n1088 & ~n1245;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~n1124 & ~n1273;
  assign n1275 = n1124 & ~n1131;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = \V1213(2)  & n1276;
  assign n1278 = ~\V1213(2)  & ~n1276;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = n1251 & n1271;
  assign n1281 = ~n1251 & ~n1271;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~n1124 & ~n1282;
  assign n1284 = n1124 & ~n1185;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = \V1213(1)  & n1285;
  assign n1287 = ~\V1213(1)  & ~n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = n1257 & n1280;
  assign n1290 = ~n1257 & ~n1280;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1124 & ~n1291;
  assign n1293 = n1124 & ~n1226;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = \V1213(0)  & n1294;
  assign n1296 = ~\V1213(0)  & ~n1294;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = \V288(0)  & ~n1234;
  assign n1299 = n1297 & n1298;
  assign n1300 = n1288 & n1299;
  assign n1301 = n1279 & n1300;
  assign n1302 = n1270 & n1301;
  assign n1303 = ~\V288(1)  & ~\V288(0) ;
  assign n1304 = ~n1085 & n1267;
  assign n1305 = n1085 & ~n1088;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = \V1213(3)  & n1306;
  assign n1308 = ~\V1213(3)  & ~n1306;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = n1267 & n1276;
  assign n1311 = ~n1267 & ~n1276;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n1085 & ~n1312;
  assign n1314 = n1085 & ~n1131;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = \V1213(2)  & n1315;
  assign n1317 = ~\V1213(2)  & ~n1315;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n1285 & n1310;
  assign n1320 = ~n1285 & ~n1310;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = ~n1085 & ~n1321;
  assign n1323 = n1085 & ~n1185;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = \V1213(1)  & n1324;
  assign n1326 = ~\V1213(1)  & ~n1324;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = n1294 & n1319;
  assign n1329 = ~n1294 & ~n1319;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~n1085 & ~n1330;
  assign n1332 = n1085 & ~n1226;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = \V1213(0)  & n1333;
  assign n1335 = ~\V1213(0)  & ~n1333;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~n1234 & n1336;
  assign n1338 = n1327 & n1337;
  assign n1339 = n1318 & n1338;
  assign n1340 = n1309 & n1339;
  assign n1341 = ~n1303 & n1340;
  assign n1342 = \V1213(3)  & n1084;
  assign n1343 = ~\V1213(3)  & ~n1084;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = \V1213(2)  & n1123;
  assign n1346 = ~\V1213(2)  & ~n1123;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = \V1213(1)  & n1173;
  assign n1349 = ~\V1213(1)  & ~n1173;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = \V1213(0)  & n1218;
  assign n1352 = ~\V1213(0)  & ~n1218;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = n1162 & ~n1234;
  assign n1355 = n1353 & n1354;
  assign n1356 = n1350 & n1355;
  assign n1357 = n1347 & n1356;
  assign n1358 = n1344 & n1357;
  assign n1359 = \V1213(3)  & ~n1084;
  assign n1360 = ~\V1213(3)  & n1084;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = n1084 & n1123;
  assign n1363 = ~n1084 & ~n1123;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = \V1213(2)  & n1364;
  assign n1366 = ~\V1213(2)  & ~n1364;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n1173 & n1362;
  assign n1369 = ~n1173 & ~n1362;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = \V1213(1)  & n1370;
  assign n1372 = ~\V1213(1)  & ~n1370;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = n1218 & n1368;
  assign n1375 = ~n1218 & ~n1368;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = \V1213(0)  & n1376;
  assign n1378 = ~\V1213(0)  & ~n1376;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = n1354 & n1379;
  assign n1381 = n1373 & n1380;
  assign n1382 = n1367 & n1381;
  assign n1383 = n1361 & n1382;
  assign n1384 = ~n1084 & ~n1116;
  assign n1385 = ~n1084 & n1116;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = \V1213(3)  & n1386;
  assign n1388 = ~\V1213(3)  & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1084 & n1364;
  assign n1391 = n1084 & ~n1364;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~n1116 & ~n1392;
  assign n1394 = n1116 & ~n1123;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = \V1213(2)  & n1395;
  assign n1397 = ~\V1213(2)  & ~n1395;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = n1370 & n1390;
  assign n1400 = ~n1370 & ~n1390;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1116 & ~n1401;
  assign n1403 = n1116 & ~n1173;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = \V1213(1)  & n1404;
  assign n1406 = ~\V1213(1)  & ~n1404;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = n1376 & n1399;
  assign n1409 = ~n1376 & ~n1399;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1116 & ~n1410;
  assign n1412 = n1116 & ~n1218;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = \V1213(0)  & n1413;
  assign n1415 = ~\V1213(0)  & ~n1413;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = \V288(2)  & ~n1234;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1407 & n1418;
  assign n1420 = n1398 & n1419;
  assign n1421 = n1389 & n1420;
  assign n1422 = ~\V288(3)  & ~\V288(2) ;
  assign n1423 = ~n1081 & n1386;
  assign n1424 = n1081 & ~n1084;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = \V1213(3)  & n1425;
  assign n1427 = ~\V1213(3)  & ~n1425;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = n1386 & n1395;
  assign n1430 = ~n1386 & ~n1395;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1081 & ~n1431;
  assign n1433 = n1081 & ~n1123;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = \V1213(2)  & n1434;
  assign n1436 = ~\V1213(2)  & ~n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = n1404 & n1429;
  assign n1439 = ~n1404 & ~n1429;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1081 & ~n1440;
  assign n1442 = n1081 & ~n1173;
  assign n1443 = ~n1441 & ~n1442;
  assign n1444 = \V1213(1)  & n1443;
  assign n1445 = ~\V1213(1)  & ~n1443;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = n1413 & n1438;
  assign n1448 = ~n1413 & ~n1438;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~n1081 & ~n1449;
  assign n1451 = n1081 & ~n1218;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = \V1213(0)  & n1452;
  assign n1454 = ~\V1213(0)  & ~n1452;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n1234 & n1455;
  assign n1457 = n1446 & n1456;
  assign n1458 = n1437 & n1457;
  assign n1459 = n1428 & n1458;
  assign n1460 = ~n1422 & n1459;
  assign n1461 = ~n1421 & ~n1460;
  assign n1462 = ~n1383 & n1461;
  assign n1463 = ~n1358 & n1462;
  assign n1464 = ~n1341 & n1463;
  assign n1465 = ~n1302 & n1464;
  assign n1466 = ~n1264 & n1465;
  assign n1467 = ~n1239 & n1466;
  assign n1468 = ~\V1536(0)  & ~n1467;
  assign n1469 = \V56(0)  & ~n513;
  assign n1470 = n816 & n1469;
  assign n1471 = \V1536(0)  & ~n1470;
  assign \V1512(1)  = n1468 | n1471;
  assign n1473 = \V288(7)  & \V288(6) ;
  assign n1474 = ~n1234 & n1473;
  assign n1475 = ~\V1213(0)  & n1474;
  assign n1476 = ~\V1213(1)  & n1475;
  assign n1477 = \V1213(2)  & n1476;
  assign n1478 = \V1213(3)  & n1477;
  assign n1479 = ~\V1213(3)  & n1477;
  assign n1480 = \V1213(3)  & n1080;
  assign n1481 = ~\V1213(3)  & ~n1080;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = \V1213(2)  & n1115;
  assign n1484 = ~\V1213(2)  & ~n1115;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = \V1213(1)  & n1161;
  assign n1487 = ~\V1213(1)  & ~n1161;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = \V1213(0)  & n1210;
  assign n1490 = ~\V1213(0)  & ~n1210;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = n1150 & ~n1234;
  assign n1493 = n1491 & n1492;
  assign n1494 = n1488 & n1493;
  assign n1495 = n1485 & n1494;
  assign n1496 = n1482 & n1495;
  assign n1497 = \V1213(3)  & ~n1080;
  assign n1498 = ~\V1213(3)  & n1080;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = n1080 & n1115;
  assign n1501 = ~n1080 & ~n1115;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = \V1213(2)  & n1502;
  assign n1504 = ~\V1213(2)  & ~n1502;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = n1161 & n1500;
  assign n1507 = ~n1161 & ~n1500;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = \V1213(1)  & n1508;
  assign n1510 = ~\V1213(1)  & ~n1508;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = n1210 & n1506;
  assign n1513 = ~n1210 & ~n1506;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = \V1213(0)  & n1514;
  assign n1516 = ~\V1213(0)  & ~n1514;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = n1492 & n1517;
  assign n1519 = n1511 & n1518;
  assign n1520 = n1505 & n1519;
  assign n1521 = n1499 & n1520;
  assign n1522 = ~n1496 & ~n1521;
  assign n1523 = ~n1383 & n1522;
  assign n1524 = ~n1358 & n1523;
  assign n1525 = ~n1264 & n1524;
  assign n1526 = ~n1239 & n1525;
  assign n1527 = ~n1479 & n1526;
  assign n1528 = ~n1478 & n1527;
  assign n1529 = ~\V1536(0)  & ~n1528;
  assign n1530 = n816 & \V1536(0) ;
  assign \V1512(3)  = n1529 | n1530;
  assign n1532 = ~n1080 & ~n1108;
  assign n1533 = ~n1080 & n1108;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = \V1213(3)  & n1534;
  assign n1536 = ~\V1213(3)  & ~n1534;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1080 & n1502;
  assign n1539 = n1080 & ~n1502;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1108 & ~n1540;
  assign n1542 = n1108 & ~n1115;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = \V1213(2)  & n1543;
  assign n1545 = ~\V1213(2)  & ~n1543;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = n1508 & n1538;
  assign n1548 = ~n1508 & ~n1538;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1108 & ~n1549;
  assign n1551 = n1108 & ~n1161;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = \V1213(1)  & n1552;
  assign n1554 = ~\V1213(1)  & ~n1552;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = n1514 & n1547;
  assign n1557 = ~n1514 & ~n1547;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~n1108 & ~n1558;
  assign n1560 = n1108 & ~n1210;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = \V1213(0)  & n1561;
  assign n1563 = ~\V1213(0)  & ~n1561;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = \V288(4)  & ~n1234;
  assign n1566 = n1564 & n1565;
  assign n1567 = n1555 & n1566;
  assign n1568 = n1546 & n1567;
  assign n1569 = n1537 & n1568;
  assign n1570 = ~\V288(5)  & ~\V288(4) ;
  assign n1571 = ~n1077 & n1534;
  assign n1572 = n1077 & ~n1080;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = \V1213(3)  & n1573;
  assign n1575 = ~\V1213(3)  & ~n1573;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = n1534 & n1543;
  assign n1578 = ~n1534 & ~n1543;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1077 & ~n1579;
  assign n1581 = n1077 & ~n1115;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = \V1213(2)  & n1582;
  assign n1584 = ~\V1213(2)  & ~n1582;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = n1552 & n1577;
  assign n1587 = ~n1552 & ~n1577;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n1077 & ~n1588;
  assign n1590 = n1077 & ~n1161;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = \V1213(1)  & n1591;
  assign n1593 = ~\V1213(1)  & ~n1591;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = n1561 & n1586;
  assign n1596 = ~n1561 & ~n1586;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1077 & ~n1597;
  assign n1599 = n1077 & ~n1210;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = \V1213(0)  & n1600;
  assign n1602 = ~\V1213(0)  & ~n1600;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1234 & n1603;
  assign n1605 = n1594 & n1604;
  assign n1606 = n1585 & n1605;
  assign n1607 = n1576 & n1606;
  assign n1608 = ~n1570 & n1607;
  assign n1609 = ~n1569 & ~n1608;
  assign n1610 = ~n1521 & n1609;
  assign n1611 = ~n1496 & n1610;
  assign n1612 = ~n1341 & n1611;
  assign n1613 = ~n1302 & n1612;
  assign n1614 = ~n1264 & n1613;
  assign n1615 = ~n1239 & n1614;
  assign n1616 = ~\V1536(0)  & ~n1615;
  assign n1617 = ~n1059 & ~n1469;
  assign n1618 = n816 & n1617;
  assign n1619 = \V1536(0)  & ~n1618;
  assign \V1512(2)  = n1616 | n1619;
  assign n1621 = \V108(2)  & ~n995;
  assign n1622 = n522 & n797;
  assign \V1898(0)  = n1621 | n1622;
  assign n1624 = ~n485 & ~n600;
  assign n1625 = ~n488 & n1624;
  assign n1626 = n602 & ~n1625;
  assign n1627 = ~\V289(0)  & ~\V249(0) ;
  assign n1628 = ~\V290(0)  & n1627;
  assign n1629 = \V295(0)  & n1628;
  assign n1630 = n540 & n1629;
  assign \V1652(0)  = n1626 | ~n1630;
  assign n1632 = \V199(2)  & \V199(4) ;
  assign n1633 = \V199(0)  & n1632;
  assign n1634 = \V194(3)  & n1633;
  assign n1635 = \V194(1)  & n1634;
  assign n1636 = \V194(2)  & n1635;
  assign n1637 = \V194(4)  & n1636;
  assign n1638 = \V199(1)  & n1637;
  assign n1639 = \V199(3)  & n1638;
  assign n1640 = \V194(0)  & n1639;
  assign n1641 = ~n639 & ~\V1536(0) ;
  assign n1642 = n1640 & n1641;
  assign n1643 = \V242(0)  & \V14(0) ;
  assign n1644 = n638 & n1643;
  assign \V1726(0)  = n1642 | n1644;
  assign n1646 = \V149(3)  & n1003;
  assign n1647 = n502 & n1646;
  assign n1648 = \V149(4)  & n1230;
  assign n1649 = ~\V149(3)  & n1648;
  assign n1650 = n502 & n1649;
  assign n1651 = \V118(5)  & ~n1650;
  assign n1652 = n947 & n1651;
  assign n1653 = ~n1647 & n1652;
  assign n1654 = \V132(7)  & n1650;
  assign n1655 = ~n947 & n1654;
  assign n1656 = ~n1647 & n1655;
  assign \V1953(7)  = n1653 | n1656;
  assign n1658 = \V118(4)  & ~n1650;
  assign n1659 = n947 & n1658;
  assign n1660 = ~n1647 & n1659;
  assign n1661 = \V132(6)  & n1650;
  assign n1662 = ~n947 & n1661;
  assign n1663 = ~n1647 & n1662;
  assign \V1953(6)  = n1660 | n1663;
  assign n1665 = ~n547 & ~n579;
  assign n1666 = n599 & ~n1036;
  assign n1667 = ~n1665 & n1666;
  assign n1668 = \V59(0)  & ~n1667;
  assign n1669 = \V62(0)  & n580;
  assign n1670 = ~n1043 & ~n1669;
  assign n1671 = ~n1668 & n1670;
  assign n1672 = \V15(0)  & \V16(0) ;
  assign \V1757(0)  = n935 | n1672;
  assign n1674 = ~n818 & ~\V1757(0) ;
  assign \V410(0)  = n1671 | ~n1674;
  assign n1676 = \V132(1)  & n1650;
  assign n1677 = ~n947 & n1676;
  assign \V1953(1)  = ~n1647 & n1677;
  assign n1679 = \V108(5)  & ~n1650;
  assign n1680 = ~n947 & n1679;
  assign n1681 = n1647 & n1680;
  assign n1682 = \V132(0)  & n1650;
  assign n1683 = ~n947 & n1682;
  assign n1684 = ~n1647 & n1683;
  assign \V1953(0)  = n1681 | n1684;
  assign n1686 = \V118(1)  & ~n1650;
  assign n1687 = n947 & n1686;
  assign n1688 = ~n1647 & n1687;
  assign n1689 = \V132(3)  & n1650;
  assign n1690 = ~n947 & n1689;
  assign n1691 = ~n1647 & n1690;
  assign \V1953(3)  = n1688 | n1691;
  assign n1693 = \V118(0)  & ~n1650;
  assign n1694 = n947 & n1693;
  assign n1695 = ~n1647 & n1694;
  assign n1696 = \V132(2)  & n1650;
  assign n1697 = ~n947 & n1696;
  assign n1698 = ~n1647 & n1697;
  assign \V1953(2)  = n1695 | n1698;
  assign n1700 = \V118(3)  & ~n1650;
  assign n1701 = n947 & n1700;
  assign n1702 = ~n1647 & n1701;
  assign n1703 = \V132(5)  & n1650;
  assign n1704 = ~n947 & n1703;
  assign n1705 = ~n1647 & n1704;
  assign \V1953(5)  = n1702 | n1705;
  assign n1707 = \V118(2)  & ~n1650;
  assign n1708 = n947 & n1707;
  assign n1709 = ~n1647 & n1708;
  assign n1710 = \V132(4)  & n1650;
  assign n1711 = ~n947 & n1710;
  assign n1712 = ~n1647 & n1711;
  assign \V1953(4)  = n1709 | n1712;
  assign n1714 = ~\V149(4)  & n504;
  assign n1715 = ~\V149(3)  & n1714;
  assign n1716 = n502 & n1715;
  assign n1717 = ~\V149(4)  & n509;
  assign n1718 = ~\V149(3)  & n1717;
  assign n1719 = n502 & n1718;
  assign n1720 = ~n1716 & ~n1719;
  assign n1721 = \V56(0)  & ~n1720;
  assign n1722 = \V62(0)  & n1719;
  assign n1723 = ~n547 & n582;
  assign n1724 = \V149(5)  & n943;
  assign n1725 = ~\V149(4)  & n1724;
  assign n1726 = ~\V149(3)  & n1725;
  assign n1727 = n502 & n1726;
  assign n1728 = ~n545 & ~n548;
  assign n1729 = ~n600 & n1728;
  assign n1730 = \V802(0)  & ~n1729;
  assign n1731 = \V149(4)  & n1002;
  assign n1732 = ~\V149(3)  & n1731;
  assign n1733 = n502 & n1732;
  assign n1734 = ~n613 & ~n1727;
  assign n1735 = ~n1733 & n1734;
  assign n1736 = \V56(0)  & ~n1735;
  assign n1737 = ~n1730 & ~n1736;
  assign n1738 = \V88(2)  & ~\V88(3) ;
  assign n1739 = ~\V88(2)  & \V88(3) ;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = \V88(0)  & ~\V88(1) ;
  assign n1742 = ~\V88(0)  & \V88(1) ;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = n1740 & ~n1743;
  assign n1745 = ~n1740 & n1743;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = \V84(4)  & ~\V84(5) ;
  assign n1748 = ~\V84(4)  & \V84(5) ;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = \V84(2)  & ~\V84(3) ;
  assign n1751 = ~\V84(2)  & \V84(3) ;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = n1749 & ~n1752;
  assign n1754 = ~n1749 & n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = n1746 & ~n1755;
  assign n1757 = ~n1746 & n1755;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~\V94(1)  & ~n1758;
  assign n1760 = \V94(1)  & n1758;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = \V84(0)  & ~\V84(1) ;
  assign n1763 = ~\V84(0)  & \V84(1) ;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = \V78(4)  & ~\V78(5) ;
  assign n1766 = ~\V78(4)  & \V78(5) ;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = n1764 & ~n1767;
  assign n1769 = ~n1764 & n1767;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = \V78(2)  & ~\V78(3) ;
  assign n1772 = ~\V78(2)  & \V78(3) ;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = \V78(0)  & ~\V78(1) ;
  assign n1775 = ~\V78(0)  & \V78(1) ;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n1773 & ~n1776;
  assign n1778 = ~n1773 & n1776;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = n1770 & ~n1779;
  assign n1781 = ~n1770 & n1779;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~\V94(0)  & ~n1782;
  assign n1784 = \V94(0)  & n1782;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = ~n1761 & ~n1785;
  assign n1787 = ~n1737 & ~n1786;
  assign n1788 = n1727 & ~n1787;
  assign n1789 = ~n600 & ~n1788;
  assign n1790 = ~n1723 & n1789;
  assign n1791 = ~n592 & n1790;
  assign n1792 = ~n488 & n1791;
  assign n1793 = \V56(0)  & ~n1792;
  assign n1794 = \V59(0)  & n583;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1722 & n1795;
  assign \V508(0)  = n1721 | ~n1796;
  assign n1798 = \V65(0)  & \V14(0) ;
  assign n1799 = ~n1719 & n1798;
  assign n1800 = ~n580 & n1799;
  assign n1801 = n824 & n1800;
  assign n1802 = \V165(6)  & n499;
  assign n1803 = \V165(3)  & n1802;
  assign n1804 = \V14(0)  & n1803;
  assign n1805 = V763 & n1804;
  assign n1806 = n824 & n1805;
  assign \V1392(0)  = n1801 | n1806;
  assign n1808 = \V32(10)  & n618;
  assign n1809 = ~n615 & n1808;
  assign n1810 = \V32(3)  & ~n623;
  assign n1811 = \V32(0)  & n623;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = n624 & ~n1812;
  assign n1814 = \V189(4)  & ~n639;
  assign n1815 = n546 & n1814;
  assign n1816 = \V229(4)  & n639;
  assign n1817 = ~n546 & n1816;
  assign n1818 = ~n1815 & ~n1817;
  assign n1819 = n540 & ~n1818;
  assign n1820 = ~n628 & n1819;
  assign n1821 = ~n637 & n1820;
  assign n1822 = \V257(5)  & ~n540;
  assign n1823 = ~n628 & n1822;
  assign n1824 = n637 & n1823;
  assign n1825 = ~n1821 & ~n1824;
  assign n1826 = ~n624 & ~n1825;
  assign n1827 = ~n1813 & ~n1826;
  assign n1828 = ~n618 & ~n1827;
  assign n1829 = n615 & n1828;
  assign \V1213(10)  = n1809 | n1829;
  assign n1831 = ~\V37(0)  & ~\V1213(10) ;
  assign n1832 = \V37(0)  & ~\V1243(7) ;
  assign \V1829(7)  = n1831 | n1832;
  assign n1834 = \V32(9)  & n618;
  assign n1835 = ~n615 & n1834;
  assign n1836 = \V32(2)  & ~n623;
  assign n1837 = ~n623 & ~n1836;
  assign n1838 = n624 & ~n1837;
  assign n1839 = \V189(3)  & ~n639;
  assign n1840 = n546 & n1839;
  assign n1841 = \V229(3)  & n639;
  assign n1842 = ~n546 & n1841;
  assign n1843 = ~n1840 & ~n1842;
  assign n1844 = n540 & ~n1843;
  assign n1845 = ~n628 & n1844;
  assign n1846 = ~n637 & n1845;
  assign n1847 = \V257(4)  & ~n540;
  assign n1848 = ~n628 & n1847;
  assign n1849 = n637 & n1848;
  assign n1850 = ~n1846 & ~n1849;
  assign n1851 = ~n624 & ~n1850;
  assign n1852 = ~n1838 & ~n1851;
  assign n1853 = ~n618 & ~n1852;
  assign n1854 = n615 & n1853;
  assign \V1213(9)  = n1835 | n1854;
  assign n1856 = ~\V37(0)  & ~\V1213(9) ;
  assign n1857 = \V37(0)  & ~\V1243(6) ;
  assign \V1829(6)  = n1856 | n1857;
  assign n1859 = ~\V37(0)  & \V321(2) ;
  assign n1860 = \V37(0)  & ~\V1243(9) ;
  assign \V1829(9)  = n1859 | n1860;
  assign n1862 = \V32(11)  & n618;
  assign n1863 = ~n615 & n1862;
  assign n1864 = \V32(4)  & ~n623;
  assign n1865 = \V32(1)  & n623;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = n624 & ~n1866;
  assign n1868 = \V189(5)  & ~n639;
  assign n1869 = n546 & n1868;
  assign n1870 = \V229(5)  & n639;
  assign n1871 = ~n546 & n1870;
  assign n1872 = ~n1869 & ~n1871;
  assign n1873 = n540 & ~n1872;
  assign n1874 = ~n628 & n1873;
  assign n1875 = ~n637 & n1874;
  assign n1876 = \V257(6)  & ~n540;
  assign n1877 = ~n628 & n1876;
  assign n1878 = n637 & n1877;
  assign n1879 = ~n1875 & ~n1878;
  assign n1880 = ~n624 & ~n1879;
  assign n1881 = ~n1867 & ~n1880;
  assign n1882 = ~n618 & ~n1881;
  assign n1883 = n615 & n1882;
  assign \V1213(11)  = n1863 | n1883;
  assign n1885 = ~\V37(0)  & ~\V1213(11) ;
  assign n1886 = \V37(0)  & ~\V1243(8) ;
  assign \V1829(8)  = n1885 | n1886;
  assign n1888 = ~\V165(5)  & ~\V165(4) ;
  assign n1889 = ~\V165(6)  & n1888;
  assign n1890 = ~\V165(7)  & n1889;
  assign n1891 = ~\V165(3)  & n1890;
  assign n1892 = ~n783 & ~n1891;
  assign n1893 = \V290(0)  & n818;
  assign n1894 = n522 & n1893;
  assign n1895 = n547 & n548;
  assign n1896 = ~\V302(0)  & n545;
  assign n1897 = ~n781 & ~n1896;
  assign n1898 = ~n1895 & n1897;
  assign n1899 = ~n791 & n1898;
  assign n1900 = ~\V289(0)  & \V14(0) ;
  assign n1901 = ~n818 & n1900;
  assign n1902 = n783 & n1901;
  assign n1903 = ~n1899 & n1902;
  assign n1904 = n783 & ~n818;
  assign n1905 = n522 & n1904;
  assign n1906 = ~n507 & n1905;
  assign n1907 = ~n1903 & n1906;
  assign n1908 = ~n1894 & ~n1907;
  assign n1909 = ~n1892 & ~n1908;
  assign n1910 = ~\V149(3)  & n992;
  assign n1911 = n502 & n1910;
  assign n1912 = \V56(0)  & n1911;
  assign n1913 = \V213(0)  & \V14(0) ;
  assign n1914 = ~n1912 & n1913;
  assign n1915 = n1908 & n1914;
  assign \V1281(0)  = n1909 | n1915;
  assign n1917 = \V174(0)  & ~n816;
  assign n1918 = ~\V302(0)  & \V292(0) ;
  assign n1919 = \V174(0)  & n818;
  assign n1920 = ~n501 & ~n1919;
  assign n1921 = ~n1918 & n1920;
  assign \V1620(0)  = n1917 | ~n1921;
  assign n1923 = \V32(4)  & n618;
  assign n1924 = ~n615 & n1923;
  assign n1925 = \V183(4)  & ~n639;
  assign n1926 = n546 & n1925;
  assign n1927 = \V223(4)  & n639;
  assign n1928 = ~n546 & n1927;
  assign n1929 = ~n1926 & ~n1928;
  assign n1930 = n540 & ~n1929;
  assign n1931 = ~n628 & n1930;
  assign n1932 = ~n637 & n1931;
  assign n1933 = ~n1878 & ~n1932;
  assign n1934 = ~n624 & ~n1933;
  assign n1935 = ~n618 & n1934;
  assign n1936 = n615 & n1935;
  assign \V1213(4)  = n1924 | n1936;
  assign n1938 = ~\V37(0)  & ~\V1213(4) ;
  assign n1939 = \V37(0)  & ~\V1243(1) ;
  assign \V1829(1)  = n1938 | n1939;
  assign n1941 = \V37(0)  & ~\V1213(2) ;
  assign \V1829(0)  = n1859 | n1941;
  assign n1943 = \V32(6)  & n618;
  assign n1944 = ~n615 & n1943;
  assign n1945 = n623 & n624;
  assign n1946 = \V189(0)  & ~n639;
  assign n1947 = n546 & n1946;
  assign n1948 = \V229(0)  & n639;
  assign n1949 = ~n546 & n1948;
  assign n1950 = ~n1947 & ~n1949;
  assign n1951 = n540 & ~n1950;
  assign n1952 = ~n628 & n1951;
  assign n1953 = ~n637 & n1952;
  assign n1954 = \V257(1)  & ~n540;
  assign n1955 = ~n628 & n1954;
  assign n1956 = n637 & n1955;
  assign n1957 = ~n1953 & ~n1956;
  assign n1958 = ~n624 & ~n1957;
  assign n1959 = ~n1945 & ~n1958;
  assign n1960 = ~n618 & ~n1959;
  assign n1961 = n615 & n1960;
  assign \V1213(6)  = n1944 | n1961;
  assign n1963 = ~\V37(0)  & ~\V1213(6) ;
  assign n1964 = \V37(0)  & ~\V1243(3) ;
  assign \V1829(3)  = n1963 | n1964;
  assign n1966 = \V32(5)  & n618;
  assign n1967 = ~n615 & n1966;
  assign n1968 = ~n623 & n624;
  assign n1969 = \V183(5)  & ~n639;
  assign n1970 = n546 & n1969;
  assign n1971 = \V223(5)  & n639;
  assign n1972 = ~n546 & n1971;
  assign n1973 = ~n1970 & ~n1972;
  assign n1974 = n540 & ~n1973;
  assign n1975 = ~n628 & n1974;
  assign n1976 = ~n637 & n1975;
  assign n1977 = \V257(0)  & ~n540;
  assign n1978 = ~n628 & n1977;
  assign n1979 = n637 & n1978;
  assign n1980 = ~n1976 & ~n1979;
  assign n1981 = ~n624 & ~n1980;
  assign n1982 = ~n1968 & ~n1981;
  assign n1983 = ~n618 & ~n1982;
  assign n1984 = n615 & n1983;
  assign \V1213(5)  = n1967 | n1984;
  assign n1986 = ~\V37(0)  & ~\V1213(5) ;
  assign n1987 = \V37(0)  & ~\V1243(2) ;
  assign \V1829(2)  = n1986 | n1987;
  assign n1989 = ~n507 & n1904;
  assign n1990 = ~n1903 & n1989;
  assign n1991 = ~n998 & n1990;
  assign n1992 = ~n1000 & ~n1991;
  assign n1993 = ~n1892 & ~n1992;
  assign n1994 = \V100(0)  & \V14(0) ;
  assign n1995 = ~n1006 & n1994;
  assign n1996 = n1992 & n1995;
  assign \V1693(0)  = n1993 | n1996;
  assign n1998 = \V32(8)  & n618;
  assign n1999 = ~n615 & n1998;
  assign n2000 = \V32(1)  & ~n623;
  assign n2001 = ~n623 & ~n2000;
  assign n2002 = n624 & ~n2001;
  assign n2003 = \V189(2)  & ~n639;
  assign n2004 = n546 & n2003;
  assign n2005 = \V229(2)  & n639;
  assign n2006 = ~n546 & n2005;
  assign n2007 = ~n2004 & ~n2006;
  assign n2008 = n540 & ~n2007;
  assign n2009 = ~n628 & n2008;
  assign n2010 = ~n637 & n2009;
  assign n2011 = \V257(3)  & ~n540;
  assign n2012 = ~n628 & n2011;
  assign n2013 = n637 & n2012;
  assign n2014 = ~n2010 & ~n2013;
  assign n2015 = ~n624 & ~n2014;
  assign n2016 = ~n2002 & ~n2015;
  assign n2017 = ~n618 & ~n2016;
  assign n2018 = n615 & n2017;
  assign \V1213(8)  = n1999 | n2018;
  assign n2020 = ~\V37(0)  & ~\V1213(8) ;
  assign n2021 = \V37(0)  & ~\V1243(5) ;
  assign \V1829(5)  = n2020 | n2021;
  assign n2023 = \V32(7)  & n618;
  assign n2024 = ~n615 & n2023;
  assign n2025 = \V32(0)  & ~n623;
  assign n2026 = ~n623 & ~n2025;
  assign n2027 = n624 & ~n2026;
  assign n2028 = \V189(1)  & ~n639;
  assign n2029 = n546 & n2028;
  assign n2030 = \V229(1)  & n639;
  assign n2031 = ~n546 & n2030;
  assign n2032 = ~n2029 & ~n2031;
  assign n2033 = n540 & ~n2032;
  assign n2034 = ~n628 & n2033;
  assign n2035 = ~n637 & n2034;
  assign n2036 = \V257(2)  & ~n540;
  assign n2037 = ~n628 & n2036;
  assign n2038 = n637 & n2037;
  assign n2039 = ~n2035 & ~n2038;
  assign n2040 = ~n624 & ~n2039;
  assign n2041 = ~n2027 & ~n2040;
  assign n2042 = ~n618 & ~n2041;
  assign n2043 = n615 & n2042;
  assign \V1213(7)  = n2024 | n2043;
  assign n2045 = ~\V37(0)  & ~\V1213(7) ;
  assign n2046 = \V37(0)  & ~\V1243(4) ;
  assign \V1829(4)  = n2045 | n2046;
  assign n2048 = \V108(1)  & ~n1911;
  assign n2049 = ~n1005 & n2048;
  assign n2050 = ~n1650 & n2049;
  assign n2051 = n994 & n2050;
  assign n2052 = \V124(1)  & ~n1911;
  assign n2053 = ~n1005 & n2052;
  assign n2054 = n1650 & n2053;
  assign n2055 = ~n994 & n2054;
  assign n2056 = \V213(1)  & n1911;
  assign n2057 = ~n1005 & n2056;
  assign n2058 = ~n1650 & n2057;
  assign n2059 = ~n994 & n2058;
  assign n2060 = \V100(1)  & ~n1911;
  assign n2061 = n1005 & n2060;
  assign n2062 = ~n1650 & n2061;
  assign n2063 = ~n994 & n2062;
  assign n2064 = ~n2059 & ~n2063;
  assign n2065 = ~n2055 & n2064;
  assign \V1921(1)  = n2051 | ~n2065;
  assign n2067 = \V108(0)  & ~n1911;
  assign n2068 = ~n1005 & n2067;
  assign n2069 = ~n1650 & n2068;
  assign n2070 = n994 & n2069;
  assign n2071 = \V124(0)  & ~n1911;
  assign n2072 = ~n1005 & n2071;
  assign n2073 = n1650 & n2072;
  assign n2074 = ~n994 & n2073;
  assign n2075 = \V213(0)  & n1911;
  assign n2076 = ~n1005 & n2075;
  assign n2077 = ~n1650 & n2076;
  assign n2078 = ~n994 & n2077;
  assign n2079 = \V100(0)  & ~n1911;
  assign n2080 = n1005 & n2079;
  assign n2081 = ~n1650 & n2080;
  assign n2082 = ~n994 & n2081;
  assign n2083 = ~n2078 & ~n2082;
  assign n2084 = ~n2074 & n2083;
  assign \V1921(0)  = n2070 | ~n2084;
  assign n2086 = \V108(3)  & ~n1911;
  assign n2087 = ~n1005 & n2086;
  assign n2088 = ~n1650 & n2087;
  assign n2089 = n994 & n2088;
  assign n2090 = \V124(3)  & ~n1911;
  assign n2091 = ~n1005 & n2090;
  assign n2092 = n1650 & n2091;
  assign n2093 = ~n994 & n2092;
  assign n2094 = \V213(3)  & n1911;
  assign n2095 = ~n1005 & n2094;
  assign n2096 = ~n1650 & n2095;
  assign n2097 = ~n994 & n2096;
  assign n2098 = \V100(3)  & ~n1911;
  assign n2099 = n1005 & n2098;
  assign n2100 = ~n1650 & n2099;
  assign n2101 = ~n994 & n2100;
  assign n2102 = ~n2097 & ~n2101;
  assign n2103 = ~n2093 & n2102;
  assign \V1921(3)  = n2089 | ~n2103;
  assign n2105 = \V108(2)  & ~n1911;
  assign n2106 = ~n1005 & n2105;
  assign n2107 = ~n1650 & n2106;
  assign n2108 = n994 & n2107;
  assign n2109 = \V124(2)  & ~n1911;
  assign n2110 = ~n1005 & n2109;
  assign n2111 = n1650 & n2110;
  assign n2112 = ~n994 & n2111;
  assign n2113 = \V213(2)  & n1911;
  assign n2114 = ~n1005 & n2113;
  assign n2115 = ~n1650 & n2114;
  assign n2116 = ~n994 & n2115;
  assign n2117 = \V100(2)  & ~n1911;
  assign n2118 = n1005 & n2117;
  assign n2119 = ~n1650 & n2118;
  assign n2120 = ~n994 & n2119;
  assign n2121 = ~n2116 & ~n2120;
  assign n2122 = ~n2112 & n2121;
  assign \V1921(2)  = n2108 | ~n2122;
  assign n2124 = \V124(5)  & ~n1911;
  assign n2125 = ~n1005 & n2124;
  assign n2126 = n1650 & n2125;
  assign n2127 = ~n994 & n2126;
  assign n2128 = \V213(5)  & n1911;
  assign n2129 = ~n1005 & n2128;
  assign n2130 = ~n1650 & n2129;
  assign n2131 = ~n994 & n2130;
  assign n2132 = \V100(5)  & ~n1911;
  assign n2133 = n1005 & n2132;
  assign n2134 = ~n1650 & n2133;
  assign n2135 = ~n994 & n2134;
  assign n2136 = ~n2131 & ~n2135;
  assign \V1921(5)  = n2127 | ~n2136;
  assign n2138 = \V108(4)  & ~n1911;
  assign n2139 = ~n1005 & n2138;
  assign n2140 = ~n1650 & n2139;
  assign n2141 = n994 & n2140;
  assign n2142 = \V124(4)  & ~n1911;
  assign n2143 = ~n1005 & n2142;
  assign n2144 = n1650 & n2143;
  assign n2145 = ~n994 & n2144;
  assign n2146 = \V213(4)  & n1911;
  assign n2147 = ~n1005 & n2146;
  assign n2148 = ~n1650 & n2147;
  assign n2149 = ~n994 & n2148;
  assign n2150 = \V100(4)  & ~n1911;
  assign n2151 = n1005 & n2150;
  assign n2152 = ~n1650 & n2151;
  assign n2153 = ~n994 & n2152;
  assign n2154 = ~n2149 & ~n2153;
  assign n2155 = ~n2145 & n2154;
  assign \V1921(4)  = n2141 | ~n2155;
  assign n2157 = \V802(0)  & n592;
  assign n2158 = ~\V279(0)  & ~n2157;
  assign n2159 = ~\V280(0)  & n2158;
  assign n2160 = \V149(4)  & n2157;
  assign n2161 = \V280(0)  & \V279(0) ;
  assign n2162 = ~n2157 & n2161;
  assign n2163 = ~n2160 & ~n2162;
  assign \V826(0)  = n2159 | ~n2163;
  assign n2165 = ~\V244(0)  & \V243(0) ;
  assign n2166 = ~n923 & n2165;
  assign n2167 = \V244(0)  & ~\V243(0) ;
  assign n2168 = ~n923 & n2167;
  assign \V591(0)  = n2166 | n2168;
  assign n2170 = \V56(0)  & n1647;
  assign n2171 = \V101(0)  & \V14(0) ;
  assign n2172 = ~n2170 & n2171;
  assign n2173 = n518 & n936;
  assign n2174 = n522 & n936;
  assign n2175 = ~n2173 & ~n2174;
  assign \V1759(0)  = n2172 | ~n2175;
  assign n2177 = \V108(5)  & ~n2170;
  assign \V1901(0)  = n936 | n2177;
  assign n2179 = \V165(4)  & n1894;
  assign n2180 = \V213(2)  & \V14(0) ;
  assign n2181 = ~n1912 & n2180;
  assign n2182 = ~n1894 & n2181;
  assign \V1297(1)  = n2179 | n2182;
  assign n2184 = \V165(3)  & n1894;
  assign n2185 = \V213(1)  & \V14(0) ;
  assign n2186 = ~n1912 & n2185;
  assign n2187 = ~n1894 & n2186;
  assign \V1297(0)  = n2184 | n2187;
  assign n2189 = \V165(6)  & n1894;
  assign n2190 = \V213(4)  & \V14(0) ;
  assign n2191 = ~n1912 & n2190;
  assign n2192 = ~n1894 & n2191;
  assign \V1297(3)  = n2189 | n2192;
  assign n2194 = \V165(5)  & n1894;
  assign n2195 = \V213(3)  & \V14(0) ;
  assign n2196 = ~n1912 & n2195;
  assign n2197 = ~n1894 & n2196;
  assign \V1297(2)  = n2194 | n2197;
  assign n2199 = \V165(7)  & n1894;
  assign n2200 = \V213(5)  & \V14(0) ;
  assign n2201 = ~n1912 & n2200;
  assign n2202 = ~n1894 & n2201;
  assign \V1297(4)  = n2199 | n2202;
  assign n2204 = \V268(3)  & \V268(5) ;
  assign n2205 = \V268(1)  & n2204;
  assign n2206 = \V268(2)  & n2205;
  assign n2207 = \V268(4)  & n2206;
  assign n2208 = \V268(0)  & n2207;
  assign n2209 = ~\V56(0)  & ~\V50(0) ;
  assign n2210 = ~\V62(0)  & n2209;
  assign n2211 = ~n540 & ~n2210;
  assign n2212 = ~n2208 & ~n2211;
  assign n2213 = ~\V258(0)  & \V14(0) ;
  assign n2214 = ~n2212 & n2213;
  assign n2215 = \V258(0)  & \V14(0) ;
  assign n2216 = n2212 & n2215;
  assign \V1451(0)  = n2214 | n2216;
  assign n2218 = ~\V248(0)  & V1719;
  assign n2219 = n1639 & n2218;
  assign n2220 = n540 & ~n1608;
  assign n2221 = ~n1569 & n2220;
  assign n2222 = n540 & ~n1521;
  assign n2223 = ~n1496 & n2222;
  assign n2224 = n2221 & n2223;
  assign n2225 = n1150 & ~n2224;
  assign n2226 = n540 & ~n1341;
  assign n2227 = ~n1302 & n2226;
  assign n2228 = n540 & ~n1264;
  assign n2229 = ~n1239 & n2228;
  assign n2230 = n2227 & n2229;
  assign n2231 = n1174 & ~n2230;
  assign n2232 = n540 & ~n1460;
  assign n2233 = ~n1421 & n2232;
  assign n2234 = n540 & ~n1383;
  assign n2235 = ~n1358 & n2234;
  assign n2236 = n2233 & n2235;
  assign n2237 = n1162 & ~n2236;
  assign n2238 = \V288(6)  & ~n1234;
  assign n2239 = ~\V1213(0)  & n2238;
  assign n2240 = ~\V1213(1)  & n2239;
  assign n2241 = ~\V1213(2)  & n2240;
  assign n2242 = \V1213(3)  & n2241;
  assign n2243 = ~\V1213(0)  & ~n1234;
  assign n2244 = ~\V1213(1)  & n2243;
  assign n2245 = ~\V1213(2)  & n2244;
  assign n2246 = ~\V1213(3)  & n2245;
  assign n2247 = ~n1149 & n2246;
  assign n2248 = n540 & ~n2247;
  assign n2249 = ~n2242 & n2248;
  assign n2250 = n540 & ~n1479;
  assign n2251 = ~n1478 & n2250;
  assign n2252 = n2249 & n2251;
  assign n2253 = \V288(6)  & ~n2252;
  assign n2254 = \V288(7)  & n2253;
  assign n2255 = ~n2237 & ~n2254;
  assign n2256 = ~n2231 & n2255;
  assign n2257 = ~n2225 & n2256;
  assign n2258 = ~\V248(0)  & \V1243(9) ;
  assign n2259 = \V1243(8)  & n2258;
  assign n2260 = \V1243(7)  & n2259;
  assign n2261 = V1719 & n2260;
  assign n2262 = ~n2257 & n2261;
  assign n2263 = \V246(0)  & n986;
  assign n2264 = \V247(0)  & ~\V248(0) ;
  assign n2265 = V1719 & n2264;
  assign n2266 = n2263 & n2265;
  assign n2267 = ~n2262 & ~n2266;
  assign \V393(0)  = n2219 | ~n2267;
  assign n2269 = \V108(3)  & ~n995;
  assign n2270 = n518 & n797;
  assign \V1899(0)  = n2269 | n2270;
  assign n2272 = ~n545 & \V1757(0) ;
  assign n2273 = \V802(0)  & \V1757(0) ;
  assign n2274 = n545 & n2273;
  assign n2275 = ~n1787 & ~n2274;
  assign \V1480(0)  = n2272 | ~n2275;
  assign n2277 = \V70(0)  & ~n540;
  assign n2278 = n540 & n1667;
  assign n2279 = \V59(0)  & ~n2278;
  assign n2280 = n540 & n599;
  assign n2281 = ~n582 & n2280;
  assign n2282 = n579 & n2281;
  assign n2283 = ~n592 & n2282;
  assign n2284 = \V802(0)  & ~n2283;
  assign n2285 = ~n580 & n1042;
  assign n2286 = ~n583 & n2285;
  assign n2287 = ~\V174(0)  & n2286;
  assign n2288 = \V56(0)  & ~n2287;
  assign n2289 = ~\V215(0)  & \V66(0) ;
  assign n2290 = V763 & n2289;
  assign n2291 = ~n818 & n2290;
  assign n2292 = \V802(0)  & n761;
  assign n2293 = ~V1719 & ~n2292;
  assign n2294 = ~n2291 & n2293;
  assign n2295 = ~n2288 & n2294;
  assign n2296 = ~n2284 & n2295;
  assign n2297 = ~n2279 & n2296;
  assign n2298 = ~n1669 & n2297;
  assign \V423(0)  = n2277 | ~n2298;
  assign n2300 = ~\V70(0)  & ~\V66(0) ;
  assign n2301 = ~\V68(0)  & n2300;
  assign n2302 = ~\V69(0)  & n2301;
  assign n2303 = \V215(0)  & \V14(0) ;
  assign n2304 = ~n2302 & n2303;
  assign n2305 = n807 & n2304;
  assign n2306 = \V216(0)  & ~\V214(0) ;
  assign \V1492(0)  = n2305 | n2306;
  assign n2308 = n819 & V1719;
  assign n2309 = n827 & V1719;
  assign n2310 = \V302(0)  & V1719;
  assign n2311 = \V215(0)  & \V66(0) ;
  assign n2312 = ~n781 & ~n1716;
  assign n2313 = ~n1719 & n2312;
  assign n2314 = ~n1727 & n2313;
  assign n2315 = \V56(0)  & ~n2314;
  assign n2316 = \V802(0)  & n545;
  assign n2317 = ~n548 & ~n600;
  assign n2318 = \V802(0)  & ~V763;
  assign n2319 = ~n2317 & n2318;
  assign n2320 = ~\V149(4)  & n610;
  assign n2321 = ~\V149(3)  & n2320;
  assign n2322 = n502 & n2321;
  assign n2323 = \V66(0)  & n2322;
  assign n2324 = \V66(0)  & V763;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n2319 & n2325;
  assign n2327 = ~n2316 & n2326;
  assign n2328 = ~n2315 & n2327;
  assign n2329 = \V32(1)  & n1185;
  assign n2330 = ~\V32(1)  & ~n1185;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = \V32(0)  & n1226;
  assign n2333 = ~\V32(0)  & ~n1226;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = \V32(2)  & n2334;
  assign n2336 = n1131 & n2335;
  assign n2337 = n2331 & n2336;
  assign n2338 = n2329 & n2334;
  assign n2339 = \V32(2)  & n1131;
  assign n2340 = ~\V32(2)  & ~n1131;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = \V32(3)  & n2334;
  assign n2343 = n2331 & n2342;
  assign n2344 = n1088 & n2343;
  assign n2345 = n2341 & n2344;
  assign n2346 = ~n2338 & ~n2345;
  assign n2347 = ~n2332 & n2346;
  assign n2348 = ~n2337 & n2347;
  assign n2349 = ~n2328 & ~n2348;
  assign n2350 = ~V763 & ~n547;
  assign n2351 = \V802(0)  & ~n2350;
  assign n2352 = ~\V214(0)  & ~\V43(0) ;
  assign n2353 = \V423(0)  & n2352;
  assign n2354 = ~\V1757(0)  & n2353;
  assign n2355 = ~n1787 & n2354;
  assign n2356 = ~n2262 & n2355;
  assign n2357 = ~n2266 & n2356;
  assign n2358 = ~n2219 & n2357;
  assign n2359 = n540 & n2358;
  assign n2360 = ~n2351 & n2359;
  assign n2361 = ~n2349 & n2360;
  assign n2362 = ~n783 & n2361;
  assign n2363 = ~n2311 & n2362;
  assign n2364 = ~n2310 & n2363;
  assign n2365 = ~n2309 & n2364;
  assign V432 = ~n2308 & n2365;
  assign n2367 = \V802(0)  & n1626;
  assign n2368 = \V59(0)  & n602;
  assign n2369 = ~n772 & n2368;
  assign n2370 = \V56(0)  & n613;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n2367 & n2371;
  assign n2373 = ~\V270(0)  & n2372;
  assign n2374 = \V62(0)  & n613;
  assign n2375 = ~\V302(0)  & ~n2374;
  assign V630 = ~n2373 & n2375;
  assign \V435(0)  = V432 | V630;
  assign n2378 = ~\V78(3)  & n613;
  assign n2379 = ~n613 & ~\V1213(11) ;
  assign \V1781(1)  = n2378 | n2379;
  assign n2381 = ~\V78(2)  & n613;
  assign n2382 = ~n613 & ~\V1213(10) ;
  assign \V1781(0)  = n2381 | n2382;
  assign n2384 = ~\V13(0)  & \V10(0) ;
  assign V1256 = \V2(0)  & n2384;
  assign n2386 = ~\V60(0)  & ~\V63(0) ;
  assign n2387 = n613 & ~n2386;
  assign n2388 = ~\V57(0)  & n1727;
  assign n2389 = ~n592 & n1035;
  assign n2390 = n579 & n2389;
  assign n2391 = ~n582 & n2390;
  assign n2392 = n599 & n2391;
  assign n2393 = ~n600 & n2392;
  assign n2394 = \V57(0)  & ~n2393;
  assign n2395 = ~\V35(0)  & ~\V174(0) ;
  assign n2396 = \V12(0)  & n2395;
  assign n2397 = \V2(0)  & n2396;
  assign n2398 = ~n2394 & n2397;
  assign n2399 = ~n2388 & n2398;
  assign V1257 = ~n2387 & n2399;
  assign V1260 = \V11(0)  & \V3(0) ;
  assign V1261 = ~\V62(0)  & V1260;
  assign V1262 = \V4(0)  & n2384;
  assign V1264 = \V4(0)  & \V12(0) ;
  assign V1265 = \V52(0)  & V1264;
  assign V1266 = \V11(0)  & \V4(0) ;
  assign V1267 = \V11(0)  & \V2(0) ;
  assign n2408 = \V258(0)  & n2208;
  assign n2409 = \V259(0)  & n2408;
  assign n2410 = ~\V258(0)  & n2211;
  assign n2411 = ~\V259(0)  & n2410;
  assign n2412 = ~n2409 & ~n2411;
  assign n2413 = \V14(0)  & ~\V260(0) ;
  assign n2414 = ~n2412 & n2413;
  assign n2415 = \V14(0)  & \V260(0) ;
  assign n2416 = n2412 & n2415;
  assign \V1467(0)  = n2414 | n2416;
  assign n2418 = \V62(0)  & \V14(0) ;
  assign n2419 = ~n1716 & n2418;
  assign n2420 = n599 & n2419;
  assign n2421 = ~n1036 & n2420;
  assign n2422 = ~n1665 & n2421;
  assign n2423 = n540 & n2422;
  assign n2424 = ~n1727 & n2423;
  assign n2425 = ~n791 & n2424;
  assign V1365 = n824 & n2425;
  assign n2427 = ~\V268(0)  & n2207;
  assign n2428 = \V268(0)  & ~n2207;
  assign V1370 = n2427 | n2428;
  assign n2430 = \V268(2)  & n2204;
  assign n2431 = \V268(4)  & n2430;
  assign n2432 = ~\V268(1)  & n2431;
  assign n2433 = \V268(1)  & ~n2431;
  assign V1371 = n2432 | n2433;
  assign n2435 = \V268(4)  & n2204;
  assign n2436 = ~\V268(2)  & n2435;
  assign n2437 = \V268(2)  & ~n2435;
  assign V1372 = n2436 | n2437;
  assign n2439 = \V268(5)  & \V268(4) ;
  assign n2440 = ~\V268(3)  & n2439;
  assign n2441 = \V268(3)  & ~n2439;
  assign V1373 = n2440 | n2441;
  assign n2443 = \V268(5)  & ~\V268(4) ;
  assign n2444 = ~\V268(5)  & \V268(4) ;
  assign V1374 = n2443 | n2444;
  assign n2446 = \V802(0)  & ~n638;
  assign V782 = \V7(0)  & n2384;
  assign V1378 = n2446 & V782;
  assign n2449 = \V248(0)  & ~\V802(0) ;
  assign n2450 = ~\V802(0)  & ~n602;
  assign n2451 = n485 & n2450;
  assign n2452 = ~n1640 & n2451;
  assign n2453 = ~n775 & n2452;
  assign n2454 = ~n2449 & n2453;
  assign n2455 = ~\V802(0)  & n1640;
  assign n2456 = ~\V802(0)  & n602;
  assign n2457 = ~n638 & ~n775;
  assign n2458 = ~n2456 & n2457;
  assign n2459 = ~n2455 & n2458;
  assign n2460 = ~n2449 & n2459;
  assign n2461 = ~\V274(0)  & \V271(0) ;
  assign n2462 = ~n613 & n2461;
  assign n2463 = \V134(1)  & \V134(0) ;
  assign n2464 = n602 & n2463;
  assign n2465 = ~n1640 & n2464;
  assign n2466 = n2462 & n2465;
  assign n2467 = ~n2460 & ~n2466;
  assign n2468 = ~n2454 & n2467;
  assign V1380 = V782 & ~n2468;
  assign n2470 = \V802(0)  & ~n1728;
  assign n2471 = ~n592 & ~n2470;
  assign V1382 = V782 & ~n2471;
  assign n2473 = \V56(0)  & ~n1787;
  assign n2474 = ~n818 & n2473;
  assign n2475 = n1733 & n2474;
  assign n2476 = \V7(0)  & n2475;
  assign V1384 = n2384 & n2476;
  assign V1386 = n2211 & V782;
  assign V1426 = \V1(0)  & n2384;
  assign V1428 = \V11(0)  & \V1(0) ;
  assign V1429 = \V12(0)  & \V1(0) ;
  assign n2482 = \V66(0)  & \V14(0) ;
  assign V1432 = n824 & n2482;
  assign n2484 = \V14(0)  & \V67(0) ;
  assign n2485 = ~n2322 & n2484;
  assign V1470 = n824 & n2485;
  assign n2487 = \V149(7)  & n2316;
  assign n2488 = ~n1903 & ~n2487;
  assign \V1645(0)  = n2349 | ~n2488;
  assign n2490 = \V68(0)  & \V14(0) ;
  assign V1537 = n824 & n2490;
  assign n2492 = ~\V69(0)  & ~\V50(0) ;
  assign n2493 = \V14(0)  & n824;
  assign V1539 = ~n2492 & n2493;
  assign n2495 = ~\V289(0)  & ~\V802(0) ;
  assign n2496 = n819 & n2495;
  assign n2497 = \V149(4)  & n1724;
  assign n2498 = ~\V149(3)  & n2497;
  assign n2499 = n502 & n2498;
  assign n2500 = \V262(0)  & n933;
  assign n2501 = n539 & ~n2500;
  assign n2502 = ~n1733 & n2501;
  assign n2503 = ~n1650 & n2502;
  assign n2504 = ~n1911 & n2503;
  assign n2505 = ~n1005 & n2504;
  assign n2506 = ~n947 & n2505;
  assign n2507 = ~n2499 & n2506;
  assign n2508 = n786 & ~n818;
  assign n2509 = n795 & ~n818;
  assign n2510 = n799 & ~n818;
  assign n2511 = ~n802 & ~n2510;
  assign n2512 = ~n1893 & n2511;
  assign n2513 = ~n2509 & n2512;
  assign \V1741(0)  = n2508 | ~n2513;
  assign n2515 = ~\V289(0)  & \V1741(0) ;
  assign n2516 = n2507 & n2515;
  assign n2517 = n1720 & ~n1727;
  assign n2518 = n2501 & n2517;
  assign n2519 = n2507 & n2518;
  assign n2520 = ~n1716 & ~n1727;
  assign n2521 = \V62(0)  & ~n2520;
  assign n2522 = \V65(0)  & n1719;
  assign n2523 = ~n540 & n931;
  assign n2524 = ~n1733 & ~n1911;
  assign n2525 = ~n1005 & n2524;
  assign n2526 = ~n1650 & n2525;
  assign n2527 = ~n947 & n2526;
  assign n2528 = ~n2499 & n2527;
  assign n2529 = ~n2523 & n2528;
  assign n2530 = \V56(0)  & ~n2529;
  assign n2531 = ~n2522 & ~n2530;
  assign n2532 = ~n2521 & n2531;
  assign n2533 = ~\V289(0)  & ~n821;
  assign n2534 = n816 & n2533;
  assign n2535 = n2532 & n2534;
  assign n2536 = ~n2519 & n2535;
  assign n2537 = ~n2516 & ~n2536;
  assign n2538 = ~n2496 & n2537;
  assign V1669 = ~n2323 & n2538;
  assign n2540 = \V108(0)  & ~n995;
  assign n2541 = ~n1787 & ~n2540;
  assign \V1896(0)  = n1672 | ~n2541;
  assign n2543 = ~\V290(0)  & ~\V289(0) ;
  assign n2544 = ~\V802(0)  & n2543;
  assign n2545 = n819 & n2544;
  assign V1736 = n772 & n2545;
  assign n2547 = \V262(0)  & ~n933;
  assign n2548 = ~n2210 & n2547;
  assign n2549 = \V261(0)  & ~n2548;
  assign n2550 = ~n2208 & ~n2549;
  assign V1832 = \V14(0)  & ~n2550;
  assign n2552 = ~n2408 & ~n2410;
  assign n2553 = ~\V259(0)  & \V14(0) ;
  assign n2554 = ~n2552 & n2553;
  assign n2555 = \V259(0)  & \V14(0) ;
  assign n2556 = n2552 & n2555;
  assign \V1459(0)  = n2554 | n2556;
  assign n2558 = \V48(0)  & ~n1720;
  assign n2559 = ~n947 & n2558;
  assign n2560 = \V118(6)  & n1720;
  assign n2561 = n947 & n2560;
  assign \V1960(0)  = n2559 | n2561;
  assign n2563 = \V46(0)  & ~n1720;
  assign n2564 = ~n947 & n2563;
  assign n2565 = \V118(7)  & n1720;
  assign n2566 = n947 & n2565;
  assign \V1960(1)  = n2564 | n2566;
  assign n2568 = \V1960(0)  & ~\V1960(1) ;
  assign n2569 = ~\V1960(0)  & \V1960(1) ;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~\V1953(7)  & \V1953(6) ;
  assign n2572 = \V1953(7)  & ~\V1953(6) ;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = n2570 & ~n2573;
  assign n2575 = ~n2570 & n2573;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = ~\V1953(5)  & \V1953(4) ;
  assign n2578 = \V1953(5)  & ~\V1953(4) ;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = ~\V1953(3)  & \V1953(2) ;
  assign n2581 = \V1953(3)  & ~\V1953(2) ;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n2579 & ~n2582;
  assign n2584 = ~n2579 & n2582;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = n2576 & ~n2585;
  assign n2587 = ~n2576 & n2585;
  assign \V1613(1)  = ~n2586 & ~n2587;
  assign n2589 = ~n488 & ~n1041;
  assign n2590 = ~n600 & n2589;
  assign n2591 = ~n1723 & n2590;
  assign n2592 = ~n1038 & n2591;
  assign n2593 = ~n485 & n2592;
  assign n2594 = ~n592 & n2593;
  assign n2595 = ~\V174(0)  & n507;
  assign n2596 = \V59(0)  & \V14(0) ;
  assign n2597 = ~V1719 & n2596;
  assign n2598 = ~n1233 & n2597;
  assign n2599 = ~n2595 & n2598;
  assign n2600 = ~n781 & n2599;
  assign n2601 = n824 & n2600;
  assign n2602 = n2594 & n2601;
  assign n2603 = n583 & n2418;
  assign n2604 = n824 & n2603;
  assign \V1274(0)  = n2602 | n2604;
  assign n2606 = ~\V1953(1)  & \V1953(0) ;
  assign n2607 = \V1953(1)  & ~\V1953(0) ;
  assign n2608 = ~n2606 & ~n2607;
  assign n2609 = ~\V1921(5)  & \V1921(4) ;
  assign n2610 = \V1921(5)  & ~\V1921(4) ;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = n2608 & ~n2611;
  assign n2613 = ~n2608 & n2611;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = ~\V1921(3)  & \V1921(2) ;
  assign n2616 = \V1921(3)  & ~\V1921(2) ;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = ~\V1921(1)  & \V1921(0) ;
  assign n2619 = \V1921(1)  & ~\V1921(0) ;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = n2617 & ~n2620;
  assign n2622 = ~n2617 & n2620;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = n2614 & ~n2623;
  assign n2625 = ~n2614 & n2623;
  assign \V1613(0)  = ~n2624 & ~n2625;
  assign \V1440(0)  = ~\V14(0)  | n602;
  assign n2628 = n488 & \V802(0) ;
  assign n2629 = ~\V802(0)  & ~n639;
  assign n2630 = ~n602 & n2629;
  assign n2631 = ~n2466 & ~n2630;
  assign n2632 = \V802(0)  & \V1243(3) ;
  assign n2633 = n600 & n2632;
  assign n2634 = n2631 & n2633;
  assign n2635 = ~n2628 & n2634;
  assign n2636 = \V802(0)  & n600;
  assign n2637 = \V194(4)  & n1633;
  assign n2638 = \V199(1)  & n2637;
  assign n2639 = \V199(3)  & n2638;
  assign n2640 = ~\V194(3)  & n2639;
  assign n2641 = \V194(3)  & ~n2639;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = ~n2628 & ~n2642;
  assign n2644 = ~n2631 & n2643;
  assign n2645 = ~n2636 & n2644;
  assign n2646 = \V149(7)  & \V802(0) ;
  assign n2647 = n488 & n2646;
  assign n2648 = ~n2636 & n2647;
  assign n2649 = n2631 & n2648;
  assign n2650 = ~n2645 & ~n2649;
  assign \V572(3)  = n2635 | ~n2650;
  assign n2652 = \V802(0)  & \V1243(2) ;
  assign n2653 = n600 & n2652;
  assign n2654 = n2631 & n2653;
  assign n2655 = ~n2628 & n2654;
  assign n2656 = \V194(4)  & n1634;
  assign n2657 = \V199(1)  & n2656;
  assign n2658 = \V199(3)  & n2657;
  assign n2659 = ~\V194(2)  & n2658;
  assign n2660 = \V194(2)  & ~n2658;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2628 & ~n2661;
  assign n2663 = ~n2631 & n2662;
  assign n2664 = ~n2636 & n2663;
  assign n2665 = \V149(6)  & \V802(0) ;
  assign n2666 = n488 & n2665;
  assign n2667 = ~n2636 & n2666;
  assign n2668 = n2631 & n2667;
  assign n2669 = ~n2664 & ~n2668;
  assign \V572(2)  = n2655 | ~n2669;
  assign n2671 = \V269(0)  & \V271(0) ;
  assign n2672 = ~n960 & n2671;
  assign n2673 = n959 & ~n960;
  assign \V634(0)  = ~n2672 & ~n2673;
  assign n2675 = \V199(1)  & n1632;
  assign n2676 = \V199(3)  & n2675;
  assign n2677 = ~\V199(0)  & n2676;
  assign n2678 = \V199(0)  & ~n2676;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2628 & ~n2679;
  assign n2681 = ~n2631 & n2680;
  assign n2682 = ~n2636 & n2681;
  assign n2683 = \V802(0)  & \V1243(5) ;
  assign n2684 = n600 & n2683;
  assign n2685 = n2631 & n2684;
  assign n2686 = ~n2628 & n2685;
  assign \V572(5)  = n2682 | n2686;
  assign n2688 = \V199(1)  & n1633;
  assign n2689 = \V199(3)  & n2688;
  assign n2690 = ~\V194(4)  & n2689;
  assign n2691 = \V194(4)  & ~n2689;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~n2628 & ~n2692;
  assign n2694 = ~n2631 & n2693;
  assign n2695 = ~n2636 & n2694;
  assign n2696 = \V802(0)  & \V1243(4) ;
  assign n2697 = n600 & n2696;
  assign n2698 = n2631 & n2697;
  assign n2699 = ~n2628 & n2698;
  assign \V572(4)  = n2695 | n2699;
  assign n2701 = \V277(0)  & \V14(0) ;
  assign n2702 = ~n600 & n2701;
  assign \V1439(0)  = n2499 | n2702;
  assign n2704 = \V802(0)  & \V1243(1) ;
  assign n2705 = n600 & n2704;
  assign n2706 = n2631 & n2705;
  assign n2707 = ~n2628 & n2706;
  assign n2708 = \V194(2)  & n1634;
  assign n2709 = \V194(4)  & n2708;
  assign n2710 = \V199(1)  & n2709;
  assign n2711 = \V199(3)  & n2710;
  assign n2712 = ~\V194(1)  & n2711;
  assign n2713 = \V194(1)  & ~n2711;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = ~n2628 & ~n2714;
  assign n2716 = ~n2631 & n2715;
  assign n2717 = ~n2636 & n2716;
  assign n2718 = \V149(5)  & \V802(0) ;
  assign n2719 = n488 & n2718;
  assign n2720 = ~n2636 & n2719;
  assign n2721 = n2631 & n2720;
  assign n2722 = ~n2717 & ~n2721;
  assign \V572(1)  = n2707 | ~n2722;
  assign n2724 = \V802(0)  & ~\V321(2) ;
  assign n2725 = n600 & n2724;
  assign n2726 = n2631 & n2725;
  assign n2727 = ~n2628 & n2726;
  assign n2728 = ~\V194(0)  & n1639;
  assign n2729 = \V194(0)  & ~n1639;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2628 & ~n2730;
  assign n2732 = ~n2631 & n2731;
  assign n2733 = ~n2636 & n2732;
  assign n2734 = \V149(4)  & \V802(0) ;
  assign n2735 = n488 & n2734;
  assign n2736 = ~n2636 & n2735;
  assign n2737 = n2631 & n2736;
  assign n2738 = ~n2733 & ~n2737;
  assign \V572(0)  = n2727 | ~n2738;
  assign n2740 = \V45(0)  & ~\V43(0) ;
  assign \V511(0)  = \V40(0)  | n2740;
  assign n2742 = \V199(3)  & \V199(4) ;
  assign n2743 = ~\V199(2)  & n2742;
  assign n2744 = \V199(2)  & ~n2742;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~n2628 & ~n2745;
  assign n2747 = ~n2631 & n2746;
  assign n2748 = ~n2636 & n2747;
  assign n2749 = \V802(0)  & \V1243(7) ;
  assign n2750 = n600 & n2749;
  assign n2751 = n2631 & n2750;
  assign n2752 = ~n2628 & n2751;
  assign \V572(7)  = n2748 | n2752;
  assign n2754 = \V199(3)  & n1632;
  assign n2755 = ~\V199(1)  & n2754;
  assign n2756 = \V199(1)  & ~n2754;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = ~n2628 & ~n2757;
  assign n2759 = ~n2631 & n2758;
  assign n2760 = ~n2636 & n2759;
  assign n2761 = \V802(0)  & \V1243(6) ;
  assign n2762 = n600 & n2761;
  assign n2763 = n2631 & n2762;
  assign n2764 = ~n2628 & n2763;
  assign \V572(6)  = n2760 | n2764;
  assign n2766 = ~\V199(4)  & ~n2628;
  assign n2767 = ~n2631 & n2766;
  assign n2768 = ~n2636 & n2767;
  assign n2769 = \V802(0)  & \V1243(9) ;
  assign n2770 = n600 & n2769;
  assign n2771 = n2631 & n2770;
  assign n2772 = ~n2628 & n2771;
  assign \V572(9)  = n2768 | n2772;
  assign n2774 = ~\V199(3)  & \V199(4) ;
  assign n2775 = \V199(3)  & ~\V199(4) ;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = ~n2628 & ~n2776;
  assign n2778 = ~n2631 & n2777;
  assign n2779 = ~n2636 & n2778;
  assign n2780 = \V802(0)  & \V1243(8) ;
  assign n2781 = n600 & n2780;
  assign n2782 = n2631 & n2781;
  assign n2783 = ~n2628 & n2782;
  assign \V572(8)  = n2779 | n2783;
  assign n2785 = ~n2446 & n2462;
  assign n2786 = \V134(1)  & ~n2462;
  assign n2787 = ~n2785 & n2786;
  assign n2788 = ~n2446 & n2787;
  assign n2789 = ~n2446 & ~n2462;
  assign n2790 = ~\V134(1)  & n2462;
  assign n2791 = ~n2789 & n2790;
  assign n2792 = ~n2446 & n2791;
  assign \V1992(1)  = n2788 | n2792;
  assign n2794 = \V134(0)  & ~n2462;
  assign n2795 = ~n2785 & n2794;
  assign n2796 = ~n2446 & n2795;
  assign n2797 = ~\V134(1)  & \V134(0) ;
  assign n2798 = \V134(1)  & ~\V134(0) ;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = n2462 & ~n2789;
  assign n2801 = ~n2799 & n2800;
  assign n2802 = ~n2446 & n2801;
  assign \V1992(0)  = n2796 | n2802;
  assign n2804 = ~\V247(0)  & ~n923;
  assign n2805 = n2263 & n2804;
  assign n2806 = \V247(0)  & ~n923;
  assign n2807 = ~n2263 & n2806;
  assign \V609(0)  = n2805 | n2807;
  assign n2809 = ~\V294(0)  & ~n1719;
  assign n2810 = ~n1788 & n2809;
  assign n2811 = \V59(0)  & \V91(0) ;
  assign n2812 = \V62(0)  & \V91(1) ;
  assign n2813 = ~n2811 & ~n2812;
  assign n2814 = n1727 & ~n2813;
  assign n2815 = ~\V41(0)  & \V45(0) ;
  assign n2816 = \V41(0)  & ~\V45(0) ;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n2814 & n2817;
  assign \V1629(0)  = n2810 | ~n2818;
  assign n2820 = n824 & ~n827;
  assign n2821 = ~n772 & ~n2820;
  assign n2822 = ~n819 & ~\V1741(0) ;
  assign n2823 = ~n2532 & n2822;
  assign n2824 = \V290(0)  & ~n818;
  assign n2825 = ~\V302(0)  & ~n2824;
  assign n2826 = ~\V289(0)  & n2825;
  assign n2827 = ~n2823 & n2826;
  assign n2828 = ~n2821 & n2827;
  assign n2829 = ~\V214(0)  & n2828;
  assign n2830 = ~n821 & n2829;
  assign n2831 = ~\V149(3)  & n1231;
  assign n2832 = n502 & n2831;
  assign n2833 = \V149(3)  & ~n1233;
  assign n2834 = n502 & n2833;
  assign n2835 = ~n994 & n2834;
  assign n2836 = ~n1647 & n2835;
  assign n2837 = \V149(4)  & n788;
  assign n2838 = ~\V149(3)  & n2837;
  assign n2839 = n502 & n2838;
  assign n2840 = ~n2836 & ~n2839;
  assign n2841 = ~n2832 & n2840;
  assign n2842 = ~\V302(0)  & ~n2841;
  assign n2843 = \V149(1)  & \V149(0) ;
  assign n2844 = ~\V149(2)  & n2843;
  assign n2845 = \V149(2)  & \V149(0) ;
  assign n2846 = \V149(1)  & n2845;
  assign n2847 = ~\V149(1)  & \V149(0) ;
  assign n2848 = \V149(2)  & n2847;
  assign n2849 = ~n2846 & ~n2848;
  assign n2850 = ~n2844 & n2849;
  assign n2851 = n2841 & n2850;
  assign n2852 = n540 & ~n2851;
  assign n2853 = ~n2842 & n2852;
  assign n2854 = \V14(0)  & ~n2853;
  assign \V798(0)  = ~n2830 | ~n2854;
  assign n2856 = \V248(0)  & V1719;
  assign n2857 = ~\V423(0)  & ~n2856;
  assign n2858 = ~n2262 & n2352;
  assign n2859 = ~n2266 & n2858;
  assign n2860 = ~n2219 & n2859;
  assign n2861 = ~n2857 & n2860;
  assign n2862 = ~n2351 & n2861;
  assign n2863 = ~n2310 & n2862;
  assign n2864 = ~n2309 & n2863;
  assign \V398(0)  = n2308 | ~n2864;
  assign n2866 = \V289(0)  & \V33(0) ;
  assign n2867 = ~n522 & n2866;
  assign \V1745(0)  = n507 | ~n2867;
  assign n2869 = n540 & ~n1234;
  assign n2870 = ~n1608 & n2869;
  assign n2871 = ~n1521 & n2870;
  assign n2872 = ~n1460 & n2871;
  assign n2873 = ~n1383 & n2872;
  assign n2874 = ~n1341 & n2873;
  assign n2875 = ~n1264 & n2874;
  assign n2876 = ~n2247 & n2875;
  assign V356 = ~n1479 & n2876;
  assign n2878 = n540 & ~n1569;
  assign n2879 = ~n1496 & n2878;
  assign n2880 = ~n1421 & n2879;
  assign n2881 = ~n1358 & n2880;
  assign n2882 = ~n1302 & n2881;
  assign n2883 = ~n1239 & n2882;
  assign n2884 = ~n2242 & n2883;
  assign V357 = ~n1478 & n2884;
  assign V373 = \V13(0)  & \V10(0) ;
  assign n2887 = ~\V35(0)  & ~n827;
  assign V377 = \V203(0)  & ~n2887;
  assign n2889 = \V108(1)  & ~n995;
  assign n2890 = n600 & n1787;
  assign \V1897(0)  = n2889 | n2890;
  assign n2892 = \V44(0)  & ~\V42(0) ;
  assign n2893 = ~\V44(0)  & \V42(0) ;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = ~\V39(0)  & \V38(0) ;
  assign n2896 = \V39(0)  & ~\V38(0) ;
  assign n2897 = ~n2895 & ~n2896;
  assign V512 = n2894 & n2897;
  assign n2899 = \V59(0)  & ~n599;
  assign n2900 = \V59(0)  & ~n547;
  assign n2901 = ~n579 & n2900;
  assign n2902 = \V56(0)  & n1041;
  assign n2903 = \V56(0)  & n1038;
  assign n2904 = ~n1669 & ~n2903;
  assign n2905 = ~n2902 & n2904;
  assign n2906 = ~n1037 & n2905;
  assign n2907 = ~n2901 & n2906;
  assign n2908 = ~n2899 & n2907;
  assign n2909 = ~n818 & n2352;
  assign n2910 = ~n783 & n2909;
  assign V527 = ~n2908 & n2910;
  assign V537 = n600 & \V1213(0) ;
  assign V538 = n600 & \V1213(1) ;
  assign V539 = n600 & \V1213(2) ;
  assign V540 = n600 & \V1213(3) ;
  assign V541 = n600 & \V1213(4) ;
  assign V542 = n600 & \V1213(5) ;
  assign V543 = n600 & \V1213(6) ;
  assign V544 = n600 & \V1213(7) ;
  assign V545 = n600 & \V1213(8) ;
  assign V546 = n600 & \V1213(9) ;
  assign V547 = n600 & \V1213(10) ;
  assign V548 = n600 & \V1213(11) ;
  assign V587 = ~\V243(0)  & ~n923;
  assign n2925 = \V62(0)  & ~\V214(0) ;
  assign n2926 = ~n818 & n2925;
  assign n2927 = n1719 & n2926;
  assign n2928 = ~n583 & ~n1788;
  assign n2929 = \V59(0)  & ~\V214(0) ;
  assign n2930 = ~n818 & n2929;
  assign n2931 = ~n2928 & n2930;
  assign n2932 = ~\V214(0)  & ~n818;
  assign n2933 = ~n783 & n2932;
  assign n2934 = n1793 & n2933;
  assign n2935 = ~n2931 & ~n2934;
  assign V620 = ~n2927 & n2935;
  assign V621 = \V293(0)  & n2817;
  assign n2938 = \V257(5)  & \V257(7) ;
  assign n2939 = \V257(3)  & n2938;
  assign n2940 = \V257(1)  & n2939;
  assign n2941 = \V257(2)  & n2940;
  assign n2942 = \V257(4)  & n2941;
  assign n2943 = \V257(6)  & n2942;
  assign n2944 = ~\V257(0)  & n2943;
  assign n2945 = \V257(0)  & ~n2943;
  assign V650 = n2944 | n2945;
  assign n2947 = \V257(2)  & n2939;
  assign n2948 = \V257(4)  & n2947;
  assign n2949 = \V257(6)  & n2948;
  assign n2950 = ~\V257(1)  & n2949;
  assign n2951 = \V257(1)  & ~n2949;
  assign V651 = n2950 | n2951;
  assign n2953 = \V257(4)  & n2939;
  assign n2954 = \V257(6)  & n2953;
  assign n2955 = ~\V257(2)  & n2954;
  assign n2956 = \V257(2)  & ~n2954;
  assign V652 = n2955 | n2956;
  assign n2958 = \V257(4)  & n2938;
  assign n2959 = \V257(6)  & n2958;
  assign n2960 = ~\V257(3)  & n2959;
  assign n2961 = \V257(3)  & ~n2959;
  assign V653 = n2960 | n2961;
  assign n2963 = \V257(6)  & n2938;
  assign n2964 = ~\V257(4)  & n2963;
  assign n2965 = \V257(4)  & ~n2963;
  assign V654 = n2964 | n2965;
  assign n2967 = \V257(7)  & \V257(6) ;
  assign n2968 = ~\V257(5)  & n2967;
  assign n2969 = \V257(5)  & ~n2967;
  assign V655 = n2968 | n2969;
  assign n2971 = \V257(7)  & ~\V257(6) ;
  assign n2972 = ~\V257(7)  & \V257(6) ;
  assign V656 = n2971 | n2972;
  assign n2974 = \V149(5)  & n2157;
  assign \V821(0)  = n2158 | n2974;
  assign n2976 = ~\V802(0)  & n592;
  assign n2977 = \V1243(9)  & ~n2976;
  assign n2978 = n2470 & n2977;
  assign n2979 = ~\V239(4)  & ~\V802(0) ;
  assign n2980 = n592 & n2979;
  assign n2981 = ~n2470 & n2980;
  assign \V1552(1)  = n2978 | n2981;
  assign n2983 = \V1243(8)  & ~n2976;
  assign n2984 = n2470 & n2983;
  assign n2985 = \V239(3)  & ~\V239(4) ;
  assign n2986 = ~\V239(3)  & \V239(4) ;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2470 & n2976;
  assign n2989 = ~n2987 & n2988;
  assign \V1552(0)  = n2984 | n2989;
  assign n2991 = \V70(0)  & \V14(0) ;
  assign n2992 = V763 & n2991;
  assign n2993 = ~n539 & n2992;
  assign V775 = n824 & n2993;
  assign V779 = \V6(0)  & n2384;
  assign n2996 = ~\V174(0)  & n1469;
  assign n2997 = ~\V52(0)  & ~n2996;
  assign n2998 = \V12(0)  & ~n2997;
  assign V781 = \V6(0)  & n2998;
  assign V783 = \V11(0)  & \V5(0) ;
  assign V784 = \V7(0)  & \V11(0) ;
  assign V801 = n501 & n513;
  assign n3003 = \V56(0)  & ~n2841;
  assign n3004 = \V802(0)  & ~n2853;
  assign n3005 = \V56(0)  & V763;
  assign n3006 = ~n513 & n3005;
  assign n3007 = ~n2997 & n3006;
  assign n3008 = n501 & ~n513;
  assign n3009 = ~n3007 & ~n3008;
  assign n3010 = ~n3004 & n3009;
  assign n3011 = ~n3003 & n3010;
  assign V966 = n2493 & ~n3011;
  assign n3013 = ~n592 & n639;
  assign n3014 = ~n1723 & n3013;
  assign n3015 = \V59(0)  & ~n3014;
  assign n3016 = \V56(0)  & n2841;
  assign n3017 = ~n3007 & n3016;
  assign n3018 = n2529 & n3017;
  assign n3019 = \V62(0)  & ~n540;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = ~n3015 & n3020;
  assign V986 = n2493 & ~n3021;
  assign \V1243(0)  = ~\V321(2) ;
  assign \V585(0)  = ~\V34(0) ;
  assign \V1833(0)  = ~\V261(0) ;
  assign \V1760(0)  = ~\V101(0) ;
  assign \V1495(0)  = ~\V175(0) ;
  assign \V1863(0)  = ~\V301(0) ;
  assign V1375 = ~\V268(5) ;
  assign \V1864(0)  = ~\V302(0) ;
  assign \V1481(0)  = ~\V214(0) ;
  assign \V1671(0)  = ~\V205(0) ;
  assign V657 = ~\V257(7) ;
endmodule


