// Benchmark "i8" written by ABC on Tue May 16 16:07:50 2017

module i8 ( 
    \V116(12) , \V133(5) , \V116(15) , \V133(4) , \V116(14) , \V133(1) ,
    \V133(0) , \V133(7) , \V133(6) , \V116(3) , \V133(9) , \V116(2) ,
    \V133(8) , \V116(5) , \V116(4) , \V116(1) , \V116(0) , \V116(7) ,
    \V116(6) , \V116(9) , \V116(8) , \V116(31) , \V116(30) , \V118(1) ,
    \V118(0) , \V84(13) , \V84(12) , \V84(15) , \V84(14) , \V15(13) ,
    \V15(12) , \V84(11) , \V84(10) , \V15(14) , \V15(11) , \V15(10) ,
    \V84(17) , \V84(16) , \V84(19) , \V84(18) , \V84(23) , \V84(22) ,
    \V84(25) , \V84(24) , \V84(21) , \V84(20) , \V84(27) , \V84(26) ,
    \V84(29) , \V84(28) , \V47(13) , \V47(12) , \V47(15) , \V47(14) ,
    \V84(31) , \V84(30) , \V47(11) , \V47(10) , \V47(17) , \V47(16) ,
    \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V47(25) , \V47(24) ,
    \V122(0) , \V47(21) , \V47(20) , \V47(27) , \V47(26) , \V47(29) ,
    \V47(28) , \V84(0) , \V84(1) , \V47(31) , \V84(2) , \V47(30) ,
    \V84(3) , \V84(4) , \V84(5) , \V84(6) , \V84(7) , \V84(8) , \V84(9) ,
    \V48(0) , \V50(0) , \V52(0) , \V133(10) , \V119(0) , \V47(0) ,
    \V47(1) , \V47(2) , \V47(3) , \V47(4) , \V47(5) , \V47(6) , \V47(7) ,
    \V47(8) , \V47(9) , \V49(0) , \V121(17) , \V121(16) , \V51(0) ,
    \V116(27) , \V116(26) , \V116(29) , \V116(28) , \V15(0) , \V15(1) ,
    \V15(2) , \V15(3) , \V15(4) , \V15(5) , \V15(6) , \V116(21) , \V15(7) ,
    \V116(20) , \V15(8) , \V116(23) , \V15(9) , \V116(22) , \V116(25) ,
    \V116(24) , \V116(17) , \V116(16) , \V116(19) , \V116(18) , \V116(11) ,
    \V116(10) , \V133(3) , \V116(13) , \V133(2) ,
    \V212(3) , \V212(2) , \V212(5) , \V212(4) , \V212(1) , \V212(0) ,
    \V212(7) , \V212(6) , \V212(9) , \V212(8) , \V214(0) , \V143(0) ,
    \V145(1) , \V145(0) , \V149(2) , \V149(1) , \V149(0) , \V134(0) ,
    \V136(1) , \V136(0) , \V165(11) , \V197(3) , \V165(10) , \V197(2) ,
    \V165(13) , \V197(5) , \V165(12) , \V197(4) , \V197(27) , \V197(26) ,
    \V165(14) , \V197(29) , \V197(1) , \V197(28) , \V197(0) , \V197(7) ,
    \V197(6) , \V197(21) , \V197(9) , \V197(20) , \V197(8) , \V197(23) ,
    \V197(22) , \V197(25) , \V197(24) , \V213(0) , \V197(17) , \V197(16) ,
    \V197(19) , \V197(18) , \V197(11) , \V197(10) , \V197(13) , \V197(12) ,
    \V197(15) , \V197(14) , \V142(3) , \V142(2) , \V142(5) , \V142(4) ,
    \V197(31) , \V142(1) , \V197(30) , \V142(0) , \V165(3) , \V212(11) ,
    \V165(2) , \V212(10) , \V165(5) , \V212(13) , \V165(4) , \V212(12) ,
    \V146(0) , \V212(14) , \V165(1) , \V165(0) , \V165(7) , \V165(6) ,
    \V165(9) , \V165(8) , \V150(0)   );
  input  \V116(12) , \V133(5) , \V116(15) , \V133(4) , \V116(14) ,
    \V133(1) , \V133(0) , \V133(7) , \V133(6) , \V116(3) , \V133(9) ,
    \V116(2) , \V133(8) , \V116(5) , \V116(4) , \V116(1) , \V116(0) ,
    \V116(7) , \V116(6) , \V116(9) , \V116(8) , \V116(31) , \V116(30) ,
    \V118(1) , \V118(0) , \V84(13) , \V84(12) , \V84(15) , \V84(14) ,
    \V15(13) , \V15(12) , \V84(11) , \V84(10) , \V15(14) , \V15(11) ,
    \V15(10) , \V84(17) , \V84(16) , \V84(19) , \V84(18) , \V84(23) ,
    \V84(22) , \V84(25) , \V84(24) , \V84(21) , \V84(20) , \V84(27) ,
    \V84(26) , \V84(29) , \V84(28) , \V47(13) , \V47(12) , \V47(15) ,
    \V47(14) , \V84(31) , \V84(30) , \V47(11) , \V47(10) , \V47(17) ,
    \V47(16) , \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V47(25) ,
    \V47(24) , \V122(0) , \V47(21) , \V47(20) , \V47(27) , \V47(26) ,
    \V47(29) , \V47(28) , \V84(0) , \V84(1) , \V47(31) , \V84(2) ,
    \V47(30) , \V84(3) , \V84(4) , \V84(5) , \V84(6) , \V84(7) , \V84(8) ,
    \V84(9) , \V48(0) , \V50(0) , \V52(0) , \V133(10) , \V119(0) ,
    \V47(0) , \V47(1) , \V47(2) , \V47(3) , \V47(4) , \V47(5) , \V47(6) ,
    \V47(7) , \V47(8) , \V47(9) , \V49(0) , \V121(17) , \V121(16) ,
    \V51(0) , \V116(27) , \V116(26) , \V116(29) , \V116(28) , \V15(0) ,
    \V15(1) , \V15(2) , \V15(3) , \V15(4) , \V15(5) , \V15(6) , \V116(21) ,
    \V15(7) , \V116(20) , \V15(8) , \V116(23) , \V15(9) , \V116(22) ,
    \V116(25) , \V116(24) , \V116(17) , \V116(16) , \V116(19) , \V116(18) ,
    \V116(11) , \V116(10) , \V133(3) , \V116(13) , \V133(2) ;
  output \V212(3) , \V212(2) , \V212(5) , \V212(4) , \V212(1) , \V212(0) ,
    \V212(7) , \V212(6) , \V212(9) , \V212(8) , \V214(0) , \V143(0) ,
    \V145(1) , \V145(0) , \V149(2) , \V149(1) , \V149(0) , \V134(0) ,
    \V136(1) , \V136(0) , \V165(11) , \V197(3) , \V165(10) , \V197(2) ,
    \V165(13) , \V197(5) , \V165(12) , \V197(4) , \V197(27) , \V197(26) ,
    \V165(14) , \V197(29) , \V197(1) , \V197(28) , \V197(0) , \V197(7) ,
    \V197(6) , \V197(21) , \V197(9) , \V197(20) , \V197(8) , \V197(23) ,
    \V197(22) , \V197(25) , \V197(24) , \V213(0) , \V197(17) , \V197(16) ,
    \V197(19) , \V197(18) , \V197(11) , \V197(10) , \V197(13) , \V197(12) ,
    \V197(15) , \V197(14) , \V142(3) , \V142(2) , \V142(5) , \V142(4) ,
    \V197(31) , \V142(1) , \V197(30) , \V142(0) , \V165(3) , \V212(11) ,
    \V165(2) , \V212(10) , \V165(5) , \V212(13) , \V165(4) , \V212(12) ,
    \V146(0) , \V212(14) , \V165(1) , \V165(0) , \V165(7) , \V165(6) ,
    \V165(9) , \V165(8) , \V150(0) ;
  wire n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
    n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909;
  assign n215 = ~\V133(1)  & ~\V133(2) ;
  assign n216 = \V133(5)  & n215;
  assign n217 = ~\V133(10)  & n216;
  assign n218 = ~\V133(7)  & n217;
  assign n219 = ~\V133(9)  & n218;
  assign n220 = ~\V118(0)  & n219;
  assign n221 = ~\V118(1)  & n220;
  assign n222 = \V133(7)  & n215;
  assign n223 = ~\V133(9)  & n222;
  assign n224 = ~\V133(5)  & n215;
  assign n225 = ~\V133(6)  & n224;
  assign n226 = ~\V133(9)  & n225;
  assign n227 = ~\V133(4)  & n226;
  assign n228 = \V133(9)  & ~\V133(10) ;
  assign n229 = \V116(3)  & n228;
  assign n230 = ~n227 & n229;
  assign n231 = ~n223 & n230;
  assign n232 = ~n221 & n231;
  assign n233 = ~\V133(10)  & ~n227;
  assign n234 = ~n223 & n233;
  assign n235 = n221 & n234;
  assign n236 = \V84(20)  & \V133(10) ;
  assign n237 = ~n227 & n236;
  assign n238 = ~n223 & n237;
  assign n239 = \V84(20)  & ~n227;
  assign n240 = n223 & n239;
  assign n241 = \V84(20)  & n227;
  assign n242 = ~n240 & ~n241;
  assign n243 = ~n238 & n242;
  assign n244 = ~n235 & n243;
  assign \V212(3)  = n232 | ~n244;
  assign n246 = \V116(2)  & ~\V133(10) ;
  assign n247 = \V133(9)  & n246;
  assign n248 = ~n227 & n247;
  assign n249 = ~n223 & n248;
  assign n250 = ~n221 & n249;
  assign n251 = \V84(19)  & \V133(10) ;
  assign n252 = ~n227 & n251;
  assign n253 = ~n223 & n252;
  assign n254 = \V84(19)  & ~n227;
  assign n255 = n223 & n254;
  assign n256 = \V84(19)  & n227;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~n253 & n257;
  assign n259 = ~n235 & n258;
  assign \V212(2)  = n250 | ~n259;
  assign n261 = \V116(5)  & n228;
  assign n262 = ~n227 & n261;
  assign n263 = ~n223 & n262;
  assign n264 = ~n221 & n263;
  assign n265 = \V84(22)  & \V133(10) ;
  assign n266 = ~n227 & n265;
  assign n267 = ~n223 & n266;
  assign n268 = \V84(22)  & ~n227;
  assign n269 = n223 & n268;
  assign n270 = \V84(22)  & n227;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~n267 & n271;
  assign n273 = ~n235 & n272;
  assign \V212(5)  = n264 | ~n273;
  assign n275 = \V116(4)  & n228;
  assign n276 = ~n227 & n275;
  assign n277 = ~n223 & n276;
  assign n278 = ~n221 & n277;
  assign n279 = \V84(21)  & \V133(10) ;
  assign n280 = ~n227 & n279;
  assign n281 = ~n223 & n280;
  assign n282 = \V84(21)  & ~n227;
  assign n283 = n223 & n282;
  assign n284 = \V84(21)  & n227;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n281 & n285;
  assign n287 = ~n235 & n286;
  assign \V212(4)  = n278 | ~n287;
  assign n289 = \V116(1)  & n228;
  assign n290 = ~n227 & n289;
  assign n291 = ~n223 & n290;
  assign n292 = ~n221 & n291;
  assign n293 = \V84(18)  & \V133(10) ;
  assign n294 = ~n227 & n293;
  assign n295 = ~n223 & n294;
  assign n296 = \V84(18)  & ~n227;
  assign n297 = n223 & n296;
  assign n298 = \V84(18)  & n227;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~n295 & n299;
  assign n301 = ~n235 & n300;
  assign \V212(1)  = n292 | ~n301;
  assign n303 = \V116(0)  & ~\V133(10) ;
  assign n304 = \V133(9)  & n303;
  assign n305 = ~n227 & n304;
  assign n306 = ~n223 & n305;
  assign n307 = ~n221 & n306;
  assign n308 = \V84(17)  & \V133(10) ;
  assign n309 = ~n227 & n308;
  assign n310 = ~n223 & n309;
  assign n311 = \V84(17)  & ~n227;
  assign n312 = n223 & n311;
  assign n313 = \V84(17)  & n227;
  assign n314 = ~n312 & ~n313;
  assign n315 = ~n310 & n314;
  assign n316 = ~n235 & n315;
  assign \V212(0)  = n307 | ~n316;
  assign n318 = \V116(7)  & n228;
  assign n319 = ~n227 & n318;
  assign n320 = ~n223 & n319;
  assign n321 = ~n221 & n320;
  assign n322 = \V84(24)  & \V133(10) ;
  assign n323 = ~n227 & n322;
  assign n324 = ~n223 & n323;
  assign n325 = \V84(24)  & ~n227;
  assign n326 = n223 & n325;
  assign n327 = \V84(24)  & n227;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n324 & n328;
  assign n330 = ~n235 & n329;
  assign \V212(7)  = n321 | ~n330;
  assign n332 = \V116(6)  & n228;
  assign n333 = ~n227 & n332;
  assign n334 = ~n223 & n333;
  assign n335 = ~n221 & n334;
  assign n336 = \V84(23)  & \V133(10) ;
  assign n337 = ~n227 & n336;
  assign n338 = ~n223 & n337;
  assign n339 = \V84(23)  & ~n227;
  assign n340 = n223 & n339;
  assign n341 = \V84(23)  & n227;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~n338 & n342;
  assign n344 = ~n235 & n343;
  assign \V212(6)  = n335 | ~n344;
  assign n346 = \V116(9)  & n228;
  assign n347 = ~n227 & n346;
  assign n348 = ~n223 & n347;
  assign n349 = ~n221 & n348;
  assign n350 = \V84(26)  & \V133(10) ;
  assign n351 = ~n227 & n350;
  assign n352 = ~n223 & n351;
  assign n353 = \V84(26)  & ~n227;
  assign n354 = n223 & n353;
  assign n355 = \V84(26)  & n227;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n352 & n356;
  assign n358 = ~n235 & n357;
  assign \V212(9)  = n349 | ~n358;
  assign n360 = \V116(8)  & n228;
  assign n361 = ~n227 & n360;
  assign n362 = ~n223 & n361;
  assign n363 = ~n221 & n362;
  assign n364 = \V84(25)  & \V133(10) ;
  assign n365 = ~n227 & n364;
  assign n366 = ~n223 & n365;
  assign n367 = \V84(25)  & ~n227;
  assign n368 = n223 & n367;
  assign n369 = \V84(25)  & n227;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~n366 & n370;
  assign n372 = ~n235 & n371;
  assign \V212(8)  = n363 | ~n372;
  assign n374 = \V133(1)  & \V133(2) ;
  assign n375 = ~\V133(10)  & n374;
  assign n376 = ~\V133(9)  & n375;
  assign n377 = \V133(7)  & ~\V133(10) ;
  assign n378 = ~\V133(9)  & n377;
  assign n379 = \V122(0)  & \V133(10) ;
  assign n380 = ~n378 & n379;
  assign n381 = ~n376 & n380;
  assign n382 = n376 & ~n378;
  assign n383 = \V121(17)  & n378;
  assign n384 = ~n382 & ~n383;
  assign \V214(0)  = n381 | ~n384;
  assign n386 = \V133(7)  & ~\V133(9) ;
  assign n387 = ~\V133(4)  & ~\V133(9) ;
  assign n388 = n346 & ~n387;
  assign n389 = ~n386 & n388;
  assign n390 = ~\V133(10)  & n224;
  assign n391 = ~\V133(6)  & n390;
  assign n392 = ~\V133(10)  & n215;
  assign n393 = \V133(7)  & n392;
  assign n394 = ~n391 & ~n393;
  assign n395 = ~\V133(1)  & \V133(2) ;
  assign n396 = \V133(0)  & n395;
  assign n397 = ~\V133(5)  & n396;
  assign n398 = ~\V133(10)  & n397;
  assign n399 = ~\V133(6)  & n398;
  assign n400 = \V133(1)  & ~\V133(3) ;
  assign n401 = \V133(2)  & n400;
  assign n402 = ~\V133(10)  & n401;
  assign n403 = ~\V133(10)  & n395;
  assign n404 = \V133(8)  & n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = ~n399 & n405;
  assign n407 = ~\V133(0)  & ~\V133(10) ;
  assign n408 = \V133(7)  & n407;
  assign n409 = ~\V133(5)  & ~\V133(0) ;
  assign n410 = ~\V133(10)  & n409;
  assign n411 = \V133(1)  & ~\V133(2) ;
  assign n412 = ~\V133(5)  & n411;
  assign n413 = ~\V133(10)  & n412;
  assign n414 = ~\V133(6)  & n413;
  assign n415 = \V133(1)  & ~\V133(10) ;
  assign n416 = \V133(8)  & n415;
  assign n417 = ~n414 & ~n416;
  assign n418 = ~n410 & n417;
  assign n419 = ~n408 & n418;
  assign n420 = \V133(1)  & \V133(3) ;
  assign n421 = \V133(2)  & n420;
  assign n422 = ~\V133(10)  & ~n421;
  assign n423 = n419 & n422;
  assign n424 = n406 & n423;
  assign n425 = n394 & n424;
  assign n426 = \V15(8)  & n422;
  assign n427 = n419 & n426;
  assign n428 = n406 & n427;
  assign n429 = ~n394 & n428;
  assign n430 = \V84(9)  & n422;
  assign n431 = n419 & n430;
  assign n432 = ~n406 & n431;
  assign n433 = \V47(1)  & n422;
  assign n434 = ~n419 & n433;
  assign n435 = \V47(9)  & ~n422;
  assign n436 = ~n434 & ~n435;
  assign n437 = ~n432 & n436;
  assign n438 = ~n429 & n437;
  assign n439 = ~n425 & n438;
  assign n440 = \V133(10)  & ~n439;
  assign n441 = ~n387 & n440;
  assign n442 = ~n386 & n441;
  assign n443 = ~n387 & ~n439;
  assign n444 = n386 & n443;
  assign n445 = n387 & ~n439;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n442 & n446;
  assign \V143(0)  = n389 | ~n447;
  assign n449 = ~\V133(6)  & ~\V133(9) ;
  assign n450 = ~\V133(4)  & n449;
  assign n451 = \V116(11)  & n228;
  assign n452 = ~n450 & n451;
  assign n453 = ~n386 & n452;
  assign n454 = \V15(10)  & n422;
  assign n455 = n419 & n454;
  assign n456 = n406 & n455;
  assign n457 = ~n394 & n456;
  assign n458 = \V84(11)  & n422;
  assign n459 = n419 & n458;
  assign n460 = ~n406 & n459;
  assign n461 = \V47(3)  & n422;
  assign n462 = ~n419 & n461;
  assign n463 = \V47(11)  & ~n422;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~n460 & n464;
  assign n466 = ~n457 & n465;
  assign n467 = ~n425 & n466;
  assign n468 = \V133(10)  & ~n467;
  assign n469 = ~n450 & n468;
  assign n470 = ~n386 & n469;
  assign n471 = ~n450 & ~n467;
  assign n472 = n386 & n471;
  assign n473 = n450 & ~n467;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n470 & n474;
  assign \V145(1)  = n453 | ~n475;
  assign n477 = \V116(10)  & n228;
  assign n478 = ~n450 & n477;
  assign n479 = ~n386 & n478;
  assign n480 = \V15(9)  & n422;
  assign n481 = n419 & n480;
  assign n482 = n406 & n481;
  assign n483 = ~n394 & n482;
  assign n484 = \V84(10)  & n422;
  assign n485 = n419 & n484;
  assign n486 = ~n406 & n485;
  assign n487 = \V47(2)  & n422;
  assign n488 = ~n419 & n487;
  assign n489 = \V47(10)  & ~n422;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n486 & n490;
  assign n492 = ~n483 & n491;
  assign n493 = ~n425 & n492;
  assign n494 = \V133(10)  & ~n493;
  assign n495 = ~n450 & n494;
  assign n496 = ~n386 & n495;
  assign n497 = ~n450 & ~n493;
  assign n498 = n386 & n497;
  assign n499 = n450 & ~n493;
  assign n500 = ~n498 & ~n499;
  assign n501 = ~n496 & n500;
  assign \V145(0)  = n479 | ~n501;
  assign n503 = ~\V133(9)  & \V133(3) ;
  assign n504 = ~\V133(4)  & n503;
  assign n505 = ~\V133(6)  & ~\V133(2) ;
  assign n506 = ~\V133(9)  & n505;
  assign n507 = ~\V133(4)  & n506;
  assign n508 = ~\V133(1)  & ~\V133(6) ;
  assign n509 = ~\V133(9)  & n508;
  assign n510 = ~\V133(4)  & n509;
  assign n511 = ~\V133(7)  & n402;
  assign n512 = \V84(15)  & n511;
  assign n513 = ~\V133(9)  & n512;
  assign n514 = ~\V133(4)  & n513;
  assign n515 = ~n510 & n514;
  assign n516 = ~n507 & n515;
  assign n517 = ~n504 & n516;
  assign n518 = ~n386 & n517;
  assign n519 = ~n228 & n518;
  assign n520 = \V116(15)  & ~\V133(10) ;
  assign n521 = ~n510 & n520;
  assign n522 = ~n507 & n521;
  assign n523 = ~n504 & n522;
  assign n524 = ~n386 & n523;
  assign n525 = n228 & n524;
  assign n526 = \V15(14)  & n422;
  assign n527 = n419 & n526;
  assign n528 = n406 & n527;
  assign n529 = ~n394 & n528;
  assign n530 = \V47(4)  & n422;
  assign n531 = n419 & n530;
  assign n532 = ~n406 & n531;
  assign n533 = \V47(7)  & n422;
  assign n534 = ~n419 & n533;
  assign n535 = \V47(15)  & ~n422;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n532 & n536;
  assign n538 = ~n529 & n537;
  assign n539 = ~n425 & n538;
  assign n540 = \V133(10)  & ~n539;
  assign n541 = ~n510 & n540;
  assign n542 = ~n507 & n541;
  assign n543 = ~n504 & n542;
  assign n544 = ~n386 & n543;
  assign n545 = ~n510 & ~n539;
  assign n546 = ~n507 & n545;
  assign n547 = ~n504 & n546;
  assign n548 = n386 & n547;
  assign n549 = n504 & n546;
  assign n550 = n507 & n545;
  assign n551 = n510 & ~n539;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n549 & n552;
  assign n554 = ~n548 & n553;
  assign n555 = ~n544 & n554;
  assign n556 = ~n525 & n555;
  assign \V149(2)  = n519 | ~n556;
  assign n558 = \V84(14)  & n511;
  assign n559 = ~\V133(9)  & n558;
  assign n560 = ~\V133(4)  & n559;
  assign n561 = ~n510 & n560;
  assign n562 = ~n507 & n561;
  assign n563 = ~n504 & n562;
  assign n564 = ~n386 & n563;
  assign n565 = ~n228 & n564;
  assign n566 = \V116(14)  & ~\V133(10) ;
  assign n567 = ~n510 & n566;
  assign n568 = ~n507 & n567;
  assign n569 = ~n504 & n568;
  assign n570 = ~n386 & n569;
  assign n571 = n228 & n570;
  assign n572 = \V15(13)  & n422;
  assign n573 = n419 & n572;
  assign n574 = n406 & n573;
  assign n575 = ~n394 & n574;
  assign n576 = n419 & n461;
  assign n577 = ~n406 & n576;
  assign n578 = \V47(6)  & n422;
  assign n579 = ~n419 & n578;
  assign n580 = \V47(14)  & ~n422;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n577 & n581;
  assign n583 = ~n575 & n582;
  assign n584 = ~n425 & n583;
  assign n585 = \V133(10)  & ~n584;
  assign n586 = ~n510 & n585;
  assign n587 = ~n507 & n586;
  assign n588 = ~n504 & n587;
  assign n589 = ~n386 & n588;
  assign n590 = ~n510 & ~n584;
  assign n591 = ~n507 & n590;
  assign n592 = ~n504 & n591;
  assign n593 = n386 & n592;
  assign n594 = n504 & n591;
  assign n595 = n507 & n590;
  assign n596 = n510 & ~n584;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n594 & n597;
  assign n599 = ~n593 & n598;
  assign n600 = ~n589 & n599;
  assign n601 = ~n571 & n600;
  assign \V149(1)  = n565 | ~n601;
  assign n603 = \V84(13)  & n511;
  assign n604 = ~\V133(9)  & n603;
  assign n605 = ~\V133(4)  & n604;
  assign n606 = ~n510 & n605;
  assign n607 = ~n507 & n606;
  assign n608 = ~n504 & n607;
  assign n609 = ~n386 & n608;
  assign n610 = ~n228 & n609;
  assign n611 = ~\V133(10)  & \V116(13) ;
  assign n612 = ~n510 & n611;
  assign n613 = ~n507 & n612;
  assign n614 = ~n504 & n613;
  assign n615 = ~n386 & n614;
  assign n616 = n228 & n615;
  assign n617 = \V15(12)  & n422;
  assign n618 = n419 & n617;
  assign n619 = n406 & n618;
  assign n620 = ~n394 & n619;
  assign n621 = n419 & n487;
  assign n622 = ~n406 & n621;
  assign n623 = \V47(5)  & n422;
  assign n624 = ~n419 & n623;
  assign n625 = \V47(13)  & ~n422;
  assign n626 = ~n624 & ~n625;
  assign n627 = ~n622 & n626;
  assign n628 = ~n620 & n627;
  assign n629 = ~n425 & n628;
  assign n630 = \V133(10)  & ~n629;
  assign n631 = ~n510 & n630;
  assign n632 = ~n507 & n631;
  assign n633 = ~n504 & n632;
  assign n634 = ~n386 & n633;
  assign n635 = ~n510 & ~n629;
  assign n636 = ~n507 & n635;
  assign n637 = ~n504 & n636;
  assign n638 = n386 & n637;
  assign n639 = n504 & n636;
  assign n640 = n507 & n635;
  assign n641 = n510 & ~n629;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n639 & n642;
  assign n644 = ~n638 & n643;
  assign n645 = ~n634 & n644;
  assign n646 = ~n616 & n645;
  assign \V149(0)  = n610 | ~n646;
  assign n648 = ~\V133(7)  & ~\V133(10) ;
  assign n649 = ~\V133(9)  & n648;
  assign n650 = ~\V133(10)  & ~\V133(2) ;
  assign n651 = \V133(7)  & n650;
  assign n652 = ~\V133(9)  & n651;
  assign n653 = ~\V133(1)  & ~\V133(10) ;
  assign n654 = \V133(7)  & n653;
  assign n655 = ~\V133(9)  & n654;
  assign n656 = ~\V133(10)  & ~n655;
  assign n657 = ~n652 & n656;
  assign n658 = ~n649 & n657;
  assign n659 = ~n228 & n658;
  assign n660 = \V84(0)  & \V133(10) ;
  assign n661 = ~n655 & n660;
  assign n662 = ~n652 & n661;
  assign n663 = ~n649 & n662;
  assign n664 = ~n228 & n663;
  assign n665 = \V116(0)  & ~n655;
  assign n666 = ~n652 & n665;
  assign n667 = ~n649 & n666;
  assign n668 = n228 & n667;
  assign n669 = \V49(0)  & ~n655;
  assign n670 = ~n652 & n669;
  assign n671 = n649 & n670;
  assign n672 = \V48(0)  & ~n655;
  assign n673 = n652 & n672;
  assign n674 = \V48(0)  & n655;
  assign n675 = ~n673 & ~n674;
  assign n676 = ~n671 & n675;
  assign n677 = ~n668 & n676;
  assign n678 = ~n664 & n677;
  assign \V134(0)  = n659 | ~n678;
  assign n680 = ~\V133(7)  & n650;
  assign n681 = ~\V133(9)  & n680;
  assign n682 = ~\V133(7)  & n653;
  assign n683 = ~\V133(9)  & n682;
  assign n684 = \V133(8)  & ~\V133(10) ;
  assign n685 = ~\V133(9)  & n684;
  assign n686 = \V133(7)  & ~\V133(8) ;
  assign n687 = ~\V133(9)  & n686;
  assign n688 = ~\V133(8)  & n374;
  assign n689 = ~\V133(9)  & n688;
  assign n690 = ~\V133(4)  & n689;
  assign n691 = \V52(0)  & ~\V133(10) ;
  assign n692 = ~n690 & n691;
  assign n693 = ~n687 & n692;
  assign n694 = ~n685 & n693;
  assign n695 = ~n683 & n694;
  assign n696 = n681 & n695;
  assign n697 = n683 & n694;
  assign n698 = n247 & ~n690;
  assign n699 = ~n687 & n698;
  assign n700 = ~n685 & n699;
  assign n701 = ~n683 & n700;
  assign n702 = ~n681 & n701;
  assign n703 = \V15(1)  & n422;
  assign n704 = n419 & n703;
  assign n705 = n406 & n704;
  assign n706 = ~n394 & n705;
  assign n707 = \V84(2)  & n422;
  assign n708 = n419 & n707;
  assign n709 = ~n406 & n708;
  assign n710 = \V47(2)  & ~n422;
  assign n711 = ~n425 & ~n710;
  assign n712 = ~n709 & n711;
  assign n713 = ~n706 & n712;
  assign n714 = \V133(10)  & ~n713;
  assign n715 = ~n690 & n714;
  assign n716 = ~n687 & n715;
  assign n717 = ~n690 & ~n713;
  assign n718 = n687 & n717;
  assign n719 = n690 & ~n713;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~n716 & n720;
  assign n722 = ~n702 & n721;
  assign n723 = ~n697 & n722;
  assign \V136(1)  = n696 | ~n723;
  assign n725 = n289 & ~n690;
  assign n726 = ~n687 & n725;
  assign n727 = ~n685 & n726;
  assign n728 = ~n683 & n727;
  assign n729 = ~n681 & n728;
  assign n730 = ~\V133(10)  & \V51(0) ;
  assign n731 = ~n690 & n730;
  assign n732 = ~n687 & n731;
  assign n733 = ~n685 & n732;
  assign n734 = ~n683 & n733;
  assign n735 = n681 & n734;
  assign n736 = n683 & n733;
  assign n737 = \V50(0)  & ~\V133(10) ;
  assign n738 = ~n690 & n737;
  assign n739 = ~n687 & n738;
  assign n740 = n685 & n739;
  assign n741 = \V15(0)  & n422;
  assign n742 = n419 & n741;
  assign n743 = n406 & n742;
  assign n744 = ~n394 & n743;
  assign n745 = \V84(1)  & n422;
  assign n746 = n419 & n745;
  assign n747 = ~n406 & n746;
  assign n748 = \V47(1)  & ~n422;
  assign n749 = ~n425 & ~n748;
  assign n750 = ~n747 & n749;
  assign n751 = ~n744 & n750;
  assign n752 = \V133(10)  & ~n751;
  assign n753 = ~n690 & n752;
  assign n754 = ~n687 & n753;
  assign n755 = ~n690 & ~n751;
  assign n756 = n687 & n755;
  assign n757 = n690 & ~n751;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n754 & n758;
  assign n760 = ~n740 & n759;
  assign n761 = ~n736 & n760;
  assign n762 = ~n735 & n761;
  assign \V136(0)  = n729 | ~n762;
  assign n764 = \V84(28)  & n511;
  assign n765 = ~\V133(9)  & n764;
  assign n766 = ~\V133(4)  & n765;
  assign n767 = ~n510 & n766;
  assign n768 = ~n507 & n767;
  assign n769 = ~n504 & n768;
  assign n770 = ~n386 & n769;
  assign n771 = ~n228 & n770;
  assign n772 = ~\V133(10)  & \V116(28) ;
  assign n773 = ~n510 & n772;
  assign n774 = ~n507 & n773;
  assign n775 = ~n504 & n774;
  assign n776 = ~n386 & n775;
  assign n777 = n228 & n776;
  assign n778 = \V47(13)  & n422;
  assign n779 = n419 & n778;
  assign n780 = n406 & n779;
  assign n781 = ~n394 & n780;
  assign n782 = \V47(17)  & n422;
  assign n783 = n419 & n782;
  assign n784 = ~n406 & n783;
  assign n785 = \V47(20)  & n422;
  assign n786 = ~n419 & n785;
  assign n787 = \V47(28)  & ~n422;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~n784 & n788;
  assign n790 = ~n781 & n789;
  assign n791 = ~n425 & n790;
  assign n792 = \V133(10)  & ~n791;
  assign n793 = ~n510 & n792;
  assign n794 = ~n507 & n793;
  assign n795 = ~n504 & n794;
  assign n796 = ~n386 & n795;
  assign n797 = ~n510 & ~n791;
  assign n798 = ~n507 & n797;
  assign n799 = ~n504 & n798;
  assign n800 = n386 & n799;
  assign n801 = n504 & n798;
  assign n802 = n507 & n797;
  assign n803 = n510 & ~n791;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n801 & n804;
  assign n806 = ~n800 & n805;
  assign n807 = ~n796 & n806;
  assign n808 = ~n777 & n807;
  assign \V165(11)  = n771 | ~n808;
  assign n810 = ~\V133(1)  & \V133(7) ;
  assign n811 = ~\V133(9)  & n810;
  assign n812 = ~\V133(6)  & n421;
  assign n813 = ~\V133(9)  & n812;
  assign n814 = ~\V133(4)  & n813;
  assign n815 = ~\V133(1)  & ~\V133(0) ;
  assign n816 = \V133(5)  & n815;
  assign n817 = ~\V133(9)  & n816;
  assign n818 = ~\V133(1)  & \V133(0) ;
  assign n819 = \V133(5)  & n818;
  assign n820 = ~\V133(9)  & n819;
  assign n821 = ~\V118(0)  & n820;
  assign n822 = ~\V133(5)  & ~\V133(1) ;
  assign n823 = ~\V133(6)  & n822;
  assign n824 = ~\V133(9)  & n823;
  assign n825 = ~\V133(4)  & n824;
  assign n826 = n229 & ~n825;
  assign n827 = ~n821 & n826;
  assign n828 = ~n817 & n827;
  assign n829 = ~n814 & n828;
  assign n830 = ~n811 & n829;
  assign n831 = n419 & n785;
  assign n832 = n406 & n831;
  assign n833 = ~n394 & n832;
  assign n834 = \V47(24)  & n422;
  assign n835 = n419 & n834;
  assign n836 = ~n406 & n835;
  assign n837 = \V47(27)  & n422;
  assign n838 = ~n419 & n837;
  assign n839 = \V84(3)  & ~n422;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n836 & n840;
  assign n842 = ~n833 & n841;
  assign n843 = ~n425 & n842;
  assign n844 = \V133(10)  & ~n843;
  assign n845 = ~n825 & n844;
  assign n846 = ~n821 & n845;
  assign n847 = ~n817 & n846;
  assign n848 = ~n814 & n847;
  assign n849 = ~n811 & n848;
  assign n850 = ~n825 & ~n843;
  assign n851 = ~n821 & n850;
  assign n852 = ~n817 & n851;
  assign n853 = ~n814 & n852;
  assign n854 = n811 & n853;
  assign n855 = n814 & n852;
  assign n856 = n817 & n851;
  assign n857 = n821 & n850;
  assign n858 = n825 & ~n843;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n856 & n859;
  assign n861 = ~n855 & n860;
  assign n862 = ~n854 & n861;
  assign n863 = ~n849 & n862;
  assign \V197(3)  = n830 | ~n863;
  assign n865 = \V84(27)  & n511;
  assign n866 = ~\V133(9)  & n865;
  assign n867 = ~\V133(4)  & n866;
  assign n868 = ~n510 & n867;
  assign n869 = ~n507 & n868;
  assign n870 = ~n504 & n869;
  assign n871 = ~n386 & n870;
  assign n872 = ~n228 & n871;
  assign n873 = ~\V133(10)  & \V116(27) ;
  assign n874 = ~n510 & n873;
  assign n875 = ~n507 & n874;
  assign n876 = ~n504 & n875;
  assign n877 = ~n386 & n876;
  assign n878 = n228 & n877;
  assign n879 = \V47(12)  & n422;
  assign n880 = n419 & n879;
  assign n881 = n406 & n880;
  assign n882 = ~n394 & n881;
  assign n883 = \V47(16)  & n422;
  assign n884 = n419 & n883;
  assign n885 = ~n406 & n884;
  assign n886 = \V47(19)  & n422;
  assign n887 = ~n419 & n886;
  assign n888 = \V47(27)  & ~n422;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n885 & n889;
  assign n891 = ~n882 & n890;
  assign n892 = ~n425 & n891;
  assign n893 = \V133(10)  & ~n892;
  assign n894 = ~n510 & n893;
  assign n895 = ~n507 & n894;
  assign n896 = ~n504 & n895;
  assign n897 = ~n386 & n896;
  assign n898 = ~n510 & ~n892;
  assign n899 = ~n507 & n898;
  assign n900 = ~n504 & n899;
  assign n901 = n386 & n900;
  assign n902 = n504 & n899;
  assign n903 = n507 & n898;
  assign n904 = n510 & ~n892;
  assign n905 = ~n903 & ~n904;
  assign n906 = ~n902 & n905;
  assign n907 = ~n901 & n906;
  assign n908 = ~n897 & n907;
  assign n909 = ~n878 & n908;
  assign \V165(10)  = n872 | ~n909;
  assign n911 = n247 & ~n825;
  assign n912 = ~n821 & n911;
  assign n913 = ~n817 & n912;
  assign n914 = ~n814 & n913;
  assign n915 = ~n811 & n914;
  assign n916 = n419 & n886;
  assign n917 = n406 & n916;
  assign n918 = ~n394 & n917;
  assign n919 = \V47(23)  & n422;
  assign n920 = n419 & n919;
  assign n921 = ~n406 & n920;
  assign n922 = \V47(26)  & n422;
  assign n923 = ~n419 & n922;
  assign n924 = \V84(2)  & ~n422;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n921 & n925;
  assign n927 = ~n918 & n926;
  assign n928 = ~n425 & n927;
  assign n929 = \V133(10)  & ~n928;
  assign n930 = ~n825 & n929;
  assign n931 = ~n821 & n930;
  assign n932 = ~n817 & n931;
  assign n933 = ~n814 & n932;
  assign n934 = ~n811 & n933;
  assign n935 = ~n825 & ~n928;
  assign n936 = ~n821 & n935;
  assign n937 = ~n817 & n936;
  assign n938 = ~n814 & n937;
  assign n939 = n811 & n938;
  assign n940 = n814 & n937;
  assign n941 = n817 & n936;
  assign n942 = n821 & n935;
  assign n943 = n825 & ~n928;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n941 & n944;
  assign n946 = ~n940 & n945;
  assign n947 = ~n939 & n946;
  assign n948 = ~n934 & n947;
  assign \V197(2)  = n915 | ~n948;
  assign n950 = \V84(30)  & n511;
  assign n951 = ~\V133(9)  & n950;
  assign n952 = ~\V133(4)  & n951;
  assign n953 = ~n510 & n952;
  assign n954 = ~n507 & n953;
  assign n955 = ~n504 & n954;
  assign n956 = ~n386 & n955;
  assign n957 = ~n228 & n956;
  assign n958 = \V116(30)  & ~\V133(10) ;
  assign n959 = ~n510 & n958;
  assign n960 = ~n507 & n959;
  assign n961 = ~n504 & n960;
  assign n962 = ~n386 & n961;
  assign n963 = n228 & n962;
  assign n964 = \V47(15)  & n422;
  assign n965 = n419 & n964;
  assign n966 = n406 & n965;
  assign n967 = ~n394 & n966;
  assign n968 = ~n406 & n916;
  assign n969 = \V47(22)  & n422;
  assign n970 = ~n419 & n969;
  assign n971 = \V47(30)  & ~n422;
  assign n972 = ~n970 & ~n971;
  assign n973 = ~n968 & n972;
  assign n974 = ~n967 & n973;
  assign n975 = ~n425 & n974;
  assign n976 = \V133(10)  & ~n975;
  assign n977 = ~n510 & n976;
  assign n978 = ~n507 & n977;
  assign n979 = ~n504 & n978;
  assign n980 = ~n386 & n979;
  assign n981 = ~n510 & ~n975;
  assign n982 = ~n507 & n981;
  assign n983 = ~n504 & n982;
  assign n984 = n386 & n983;
  assign n985 = n504 & n982;
  assign n986 = n507 & n981;
  assign n987 = n510 & ~n975;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n985 & n988;
  assign n990 = ~n984 & n989;
  assign n991 = ~n980 & n990;
  assign n992 = ~n963 & n991;
  assign \V165(13)  = n957 | ~n992;
  assign n994 = n261 & ~n825;
  assign n995 = ~n821 & n994;
  assign n996 = ~n817 & n995;
  assign n997 = ~n814 & n996;
  assign n998 = ~n811 & n997;
  assign n999 = n419 & n969;
  assign n1000 = n406 & n999;
  assign n1001 = ~n394 & n1000;
  assign n1002 = n419 & n922;
  assign n1003 = ~n406 & n1002;
  assign n1004 = \V47(29)  & n422;
  assign n1005 = ~n419 & n1004;
  assign n1006 = \V84(5)  & ~n422;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1003 & n1007;
  assign n1009 = ~n1001 & n1008;
  assign n1010 = ~n425 & n1009;
  assign n1011 = \V133(10)  & ~n1010;
  assign n1012 = ~n825 & n1011;
  assign n1013 = ~n821 & n1012;
  assign n1014 = ~n817 & n1013;
  assign n1015 = ~n814 & n1014;
  assign n1016 = ~n811 & n1015;
  assign n1017 = ~n825 & ~n1010;
  assign n1018 = ~n821 & n1017;
  assign n1019 = ~n817 & n1018;
  assign n1020 = ~n814 & n1019;
  assign n1021 = n811 & n1020;
  assign n1022 = n814 & n1019;
  assign n1023 = n817 & n1018;
  assign n1024 = n821 & n1017;
  assign n1025 = n825 & ~n1010;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n1023 & n1026;
  assign n1028 = ~n1022 & n1027;
  assign n1029 = ~n1021 & n1028;
  assign n1030 = ~n1016 & n1029;
  assign \V197(5)  = n998 | ~n1030;
  assign n1032 = \V84(29)  & n511;
  assign n1033 = ~\V133(9)  & n1032;
  assign n1034 = ~\V133(4)  & n1033;
  assign n1035 = ~n510 & n1034;
  assign n1036 = ~n507 & n1035;
  assign n1037 = ~n504 & n1036;
  assign n1038 = ~n386 & n1037;
  assign n1039 = ~n228 & n1038;
  assign n1040 = ~\V133(10)  & \V116(29) ;
  assign n1041 = ~n510 & n1040;
  assign n1042 = ~n507 & n1041;
  assign n1043 = ~n504 & n1042;
  assign n1044 = ~n386 & n1043;
  assign n1045 = n228 & n1044;
  assign n1046 = \V47(14)  & n422;
  assign n1047 = n419 & n1046;
  assign n1048 = n406 & n1047;
  assign n1049 = ~n394 & n1048;
  assign n1050 = \V47(18)  & n422;
  assign n1051 = n419 & n1050;
  assign n1052 = ~n406 & n1051;
  assign n1053 = \V47(21)  & n422;
  assign n1054 = ~n419 & n1053;
  assign n1055 = \V47(29)  & ~n422;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1052 & n1056;
  assign n1058 = ~n1049 & n1057;
  assign n1059 = ~n425 & n1058;
  assign n1060 = \V133(10)  & ~n1059;
  assign n1061 = ~n510 & n1060;
  assign n1062 = ~n507 & n1061;
  assign n1063 = ~n504 & n1062;
  assign n1064 = ~n386 & n1063;
  assign n1065 = ~n510 & ~n1059;
  assign n1066 = ~n507 & n1065;
  assign n1067 = ~n504 & n1066;
  assign n1068 = n386 & n1067;
  assign n1069 = n504 & n1066;
  assign n1070 = n507 & n1065;
  assign n1071 = n510 & ~n1059;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = ~n1069 & n1072;
  assign n1074 = ~n1068 & n1073;
  assign n1075 = ~n1064 & n1074;
  assign n1076 = ~n1045 & n1075;
  assign \V165(12)  = n1039 | ~n1076;
  assign n1078 = n275 & ~n825;
  assign n1079 = ~n821 & n1078;
  assign n1080 = ~n817 & n1079;
  assign n1081 = ~n814 & n1080;
  assign n1082 = ~n811 & n1081;
  assign n1083 = n419 & n1053;
  assign n1084 = n406 & n1083;
  assign n1085 = ~n394 & n1084;
  assign n1086 = \V47(25)  & n422;
  assign n1087 = n419 & n1086;
  assign n1088 = ~n406 & n1087;
  assign n1089 = \V47(28)  & n422;
  assign n1090 = ~n419 & n1089;
  assign n1091 = \V84(4)  & ~n422;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~n1088 & n1092;
  assign n1094 = ~n1085 & n1093;
  assign n1095 = ~n425 & n1094;
  assign n1096 = \V133(10)  & ~n1095;
  assign n1097 = ~n825 & n1096;
  assign n1098 = ~n821 & n1097;
  assign n1099 = ~n817 & n1098;
  assign n1100 = ~n814 & n1099;
  assign n1101 = ~n811 & n1100;
  assign n1102 = ~n825 & ~n1095;
  assign n1103 = ~n821 & n1102;
  assign n1104 = ~n817 & n1103;
  assign n1105 = ~n814 & n1104;
  assign n1106 = n811 & n1105;
  assign n1107 = n814 & n1104;
  assign n1108 = n817 & n1103;
  assign n1109 = n821 & n1102;
  assign n1110 = n825 & ~n1095;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1108 & n1111;
  assign n1113 = ~n1107 & n1112;
  assign n1114 = ~n1106 & n1113;
  assign n1115 = ~n1101 & n1114;
  assign \V197(4)  = n1082 | ~n1115;
  assign n1117 = \V116(27)  & n228;
  assign n1118 = ~n825 & n1117;
  assign n1119 = ~n821 & n1118;
  assign n1120 = ~n817 & n1119;
  assign n1121 = ~n814 & n1120;
  assign n1122 = ~n811 & n1121;
  assign n1123 = \V84(12)  & n422;
  assign n1124 = n419 & n1123;
  assign n1125 = n406 & n1124;
  assign n1126 = ~n394 & n1125;
  assign n1127 = \V84(16)  & n422;
  assign n1128 = n419 & n1127;
  assign n1129 = ~n406 & n1128;
  assign n1130 = \V84(19)  & n422;
  assign n1131 = ~n419 & n1130;
  assign n1132 = \V84(27)  & ~n422;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1129 & n1133;
  assign n1135 = ~n1126 & n1134;
  assign n1136 = ~n425 & n1135;
  assign n1137 = \V133(10)  & ~n1136;
  assign n1138 = ~n825 & n1137;
  assign n1139 = ~n821 & n1138;
  assign n1140 = ~n817 & n1139;
  assign n1141 = ~n814 & n1140;
  assign n1142 = ~n811 & n1141;
  assign n1143 = ~n825 & ~n1136;
  assign n1144 = ~n821 & n1143;
  assign n1145 = ~n817 & n1144;
  assign n1146 = ~n814 & n1145;
  assign n1147 = n811 & n1146;
  assign n1148 = n814 & n1145;
  assign n1149 = n817 & n1144;
  assign n1150 = n821 & n1143;
  assign n1151 = n825 & ~n1136;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n1149 & n1152;
  assign n1154 = ~n1148 & n1153;
  assign n1155 = ~n1147 & n1154;
  assign n1156 = ~n1142 & n1155;
  assign \V197(27)  = n1122 | ~n1156;
  assign n1158 = \V116(26)  & n228;
  assign n1159 = ~n825 & n1158;
  assign n1160 = ~n821 & n1159;
  assign n1161 = ~n817 & n1160;
  assign n1162 = ~n814 & n1161;
  assign n1163 = ~n811 & n1162;
  assign n1164 = n406 & n459;
  assign n1165 = ~n394 & n1164;
  assign n1166 = \V84(15)  & n422;
  assign n1167 = n419 & n1166;
  assign n1168 = ~n406 & n1167;
  assign n1169 = \V84(18)  & n422;
  assign n1170 = ~n419 & n1169;
  assign n1171 = \V84(26)  & ~n422;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1168 & n1172;
  assign n1174 = ~n1165 & n1173;
  assign n1175 = ~n425 & n1174;
  assign n1176 = \V133(10)  & ~n1175;
  assign n1177 = ~n825 & n1176;
  assign n1178 = ~n821 & n1177;
  assign n1179 = ~n817 & n1178;
  assign n1180 = ~n814 & n1179;
  assign n1181 = ~n811 & n1180;
  assign n1182 = ~n825 & ~n1175;
  assign n1183 = ~n821 & n1182;
  assign n1184 = ~n817 & n1183;
  assign n1185 = ~n814 & n1184;
  assign n1186 = n811 & n1185;
  assign n1187 = n814 & n1184;
  assign n1188 = n817 & n1183;
  assign n1189 = n821 & n1182;
  assign n1190 = n825 & ~n1175;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~n1188 & n1191;
  assign n1193 = ~n1187 & n1192;
  assign n1194 = ~n1186 & n1193;
  assign n1195 = ~n1181 & n1194;
  assign \V197(26)  = n1163 | ~n1195;
  assign n1197 = \V84(31)  & n511;
  assign n1198 = ~\V133(9)  & n1197;
  assign n1199 = ~\V133(4)  & n1198;
  assign n1200 = ~n510 & n1199;
  assign n1201 = ~n507 & n1200;
  assign n1202 = ~n504 & n1201;
  assign n1203 = ~n386 & n1202;
  assign n1204 = ~n228 & n1203;
  assign n1205 = \V116(31)  & ~\V133(10) ;
  assign n1206 = ~n510 & n1205;
  assign n1207 = ~n507 & n1206;
  assign n1208 = ~n504 & n1207;
  assign n1209 = ~n386 & n1208;
  assign n1210 = n228 & n1209;
  assign n1211 = n406 & n884;
  assign n1212 = ~n394 & n1211;
  assign n1213 = ~n406 & n831;
  assign n1214 = ~n419 & n919;
  assign n1215 = \V47(31)  & ~n422;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1213 & n1216;
  assign n1218 = ~n1212 & n1217;
  assign n1219 = ~n425 & n1218;
  assign n1220 = \V133(10)  & ~n1219;
  assign n1221 = ~n510 & n1220;
  assign n1222 = ~n507 & n1221;
  assign n1223 = ~n504 & n1222;
  assign n1224 = ~n386 & n1223;
  assign n1225 = ~n510 & ~n1219;
  assign n1226 = ~n507 & n1225;
  assign n1227 = ~n504 & n1226;
  assign n1228 = n386 & n1227;
  assign n1229 = n504 & n1226;
  assign n1230 = n507 & n1225;
  assign n1231 = n510 & ~n1219;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = ~n1228 & n1233;
  assign n1235 = ~n1224 & n1234;
  assign n1236 = ~n1210 & n1235;
  assign \V165(14)  = n1204 | ~n1236;
  assign n1238 = \V116(29)  & n228;
  assign n1239 = ~n825 & n1238;
  assign n1240 = ~n821 & n1239;
  assign n1241 = ~n817 & n1240;
  assign n1242 = ~n814 & n1241;
  assign n1243 = ~n811 & n1242;
  assign n1244 = \V84(14)  & n422;
  assign n1245 = n419 & n1244;
  assign n1246 = n406 & n1245;
  assign n1247 = ~n394 & n1246;
  assign n1248 = n419 & n1169;
  assign n1249 = ~n406 & n1248;
  assign n1250 = \V84(21)  & n422;
  assign n1251 = ~n419 & n1250;
  assign n1252 = \V84(29)  & ~n422;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1249 & n1253;
  assign n1255 = ~n1247 & n1254;
  assign n1256 = ~n425 & n1255;
  assign n1257 = \V133(10)  & ~n1256;
  assign n1258 = ~n825 & n1257;
  assign n1259 = ~n821 & n1258;
  assign n1260 = ~n817 & n1259;
  assign n1261 = ~n814 & n1260;
  assign n1262 = ~n811 & n1261;
  assign n1263 = ~n825 & ~n1256;
  assign n1264 = ~n821 & n1263;
  assign n1265 = ~n817 & n1264;
  assign n1266 = ~n814 & n1265;
  assign n1267 = n811 & n1266;
  assign n1268 = n814 & n1265;
  assign n1269 = n817 & n1264;
  assign n1270 = n821 & n1263;
  assign n1271 = n825 & ~n1256;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1269 & n1272;
  assign n1274 = ~n1268 & n1273;
  assign n1275 = ~n1267 & n1274;
  assign n1276 = ~n1262 & n1275;
  assign \V197(29)  = n1243 | ~n1276;
  assign n1278 = n289 & ~n825;
  assign n1279 = ~n821 & n1278;
  assign n1280 = ~n817 & n1279;
  assign n1281 = ~n814 & n1280;
  assign n1282 = ~n811 & n1281;
  assign n1283 = n406 & n1051;
  assign n1284 = ~n394 & n1283;
  assign n1285 = ~n406 & n999;
  assign n1286 = ~n419 & n1086;
  assign n1287 = \V84(1)  & ~n422;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = ~n1285 & n1288;
  assign n1290 = ~n1284 & n1289;
  assign n1291 = ~n425 & n1290;
  assign n1292 = \V133(10)  & ~n1291;
  assign n1293 = ~n825 & n1292;
  assign n1294 = ~n821 & n1293;
  assign n1295 = ~n817 & n1294;
  assign n1296 = ~n814 & n1295;
  assign n1297 = ~n811 & n1296;
  assign n1298 = ~n825 & ~n1291;
  assign n1299 = ~n821 & n1298;
  assign n1300 = ~n817 & n1299;
  assign n1301 = ~n814 & n1300;
  assign n1302 = n811 & n1301;
  assign n1303 = n814 & n1300;
  assign n1304 = n817 & n1299;
  assign n1305 = n821 & n1298;
  assign n1306 = n825 & ~n1291;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1304 & n1307;
  assign n1309 = ~n1303 & n1308;
  assign n1310 = ~n1302 & n1309;
  assign n1311 = ~n1297 & n1310;
  assign \V197(1)  = n1282 | ~n1311;
  assign n1313 = \V116(28)  & n228;
  assign n1314 = ~n825 & n1313;
  assign n1315 = ~n821 & n1314;
  assign n1316 = ~n817 & n1315;
  assign n1317 = ~n814 & n1316;
  assign n1318 = ~n811 & n1317;
  assign n1319 = \V84(13)  & n422;
  assign n1320 = n419 & n1319;
  assign n1321 = n406 & n1320;
  assign n1322 = ~n394 & n1321;
  assign n1323 = \V84(17)  & n422;
  assign n1324 = n419 & n1323;
  assign n1325 = ~n406 & n1324;
  assign n1326 = \V84(20)  & n422;
  assign n1327 = ~n419 & n1326;
  assign n1328 = \V84(28)  & ~n422;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = ~n1325 & n1329;
  assign n1331 = ~n1322 & n1330;
  assign n1332 = ~n425 & n1331;
  assign n1333 = \V133(10)  & ~n1332;
  assign n1334 = ~n825 & n1333;
  assign n1335 = ~n821 & n1334;
  assign n1336 = ~n817 & n1335;
  assign n1337 = ~n814 & n1336;
  assign n1338 = ~n811 & n1337;
  assign n1339 = ~n825 & ~n1332;
  assign n1340 = ~n821 & n1339;
  assign n1341 = ~n817 & n1340;
  assign n1342 = ~n814 & n1341;
  assign n1343 = n811 & n1342;
  assign n1344 = n814 & n1341;
  assign n1345 = n817 & n1340;
  assign n1346 = n821 & n1339;
  assign n1347 = n825 & ~n1332;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1345 & n1348;
  assign n1350 = ~n1344 & n1349;
  assign n1351 = ~n1343 & n1350;
  assign n1352 = ~n1338 & n1351;
  assign \V197(28)  = n1318 | ~n1352;
  assign n1354 = n304 & ~n825;
  assign n1355 = ~n821 & n1354;
  assign n1356 = ~n817 & n1355;
  assign n1357 = ~n814 & n1356;
  assign n1358 = ~n811 & n1357;
  assign n1359 = n406 & n783;
  assign n1360 = ~n394 & n1359;
  assign n1361 = ~n406 & n1083;
  assign n1362 = ~n419 & n834;
  assign n1363 = \V84(0)  & ~n422;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1361 & n1364;
  assign n1366 = ~n1360 & n1365;
  assign n1367 = ~n425 & n1366;
  assign n1368 = \V133(10)  & ~n1367;
  assign n1369 = ~n825 & n1368;
  assign n1370 = ~n821 & n1369;
  assign n1371 = ~n817 & n1370;
  assign n1372 = ~n814 & n1371;
  assign n1373 = ~n811 & n1372;
  assign n1374 = ~n825 & ~n1367;
  assign n1375 = ~n821 & n1374;
  assign n1376 = ~n817 & n1375;
  assign n1377 = ~n814 & n1376;
  assign n1378 = n811 & n1377;
  assign n1379 = n814 & n1376;
  assign n1380 = n817 & n1375;
  assign n1381 = n821 & n1374;
  assign n1382 = n825 & ~n1367;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n1380 & n1383;
  assign n1385 = ~n1379 & n1384;
  assign n1386 = ~n1378 & n1385;
  assign n1387 = ~n1373 & n1386;
  assign \V197(0)  = n1358 | ~n1387;
  assign n1389 = n318 & ~n825;
  assign n1390 = ~n821 & n1389;
  assign n1391 = ~n817 & n1390;
  assign n1392 = ~n814 & n1391;
  assign n1393 = ~n811 & n1392;
  assign n1394 = n406 & n835;
  assign n1395 = ~n394 & n1394;
  assign n1396 = n419 & n1089;
  assign n1397 = ~n406 & n1396;
  assign n1398 = \V47(31)  & n422;
  assign n1399 = ~n419 & n1398;
  assign n1400 = \V84(7)  & ~n422;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1397 & n1401;
  assign n1403 = ~n1395 & n1402;
  assign n1404 = ~n425 & n1403;
  assign n1405 = \V133(10)  & ~n1404;
  assign n1406 = ~n825 & n1405;
  assign n1407 = ~n821 & n1406;
  assign n1408 = ~n817 & n1407;
  assign n1409 = ~n814 & n1408;
  assign n1410 = ~n811 & n1409;
  assign n1411 = ~n825 & ~n1404;
  assign n1412 = ~n821 & n1411;
  assign n1413 = ~n817 & n1412;
  assign n1414 = ~n814 & n1413;
  assign n1415 = n811 & n1414;
  assign n1416 = n814 & n1413;
  assign n1417 = n817 & n1412;
  assign n1418 = n821 & n1411;
  assign n1419 = n825 & ~n1404;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~n1417 & n1420;
  assign n1422 = ~n1416 & n1421;
  assign n1423 = ~n1415 & n1422;
  assign n1424 = ~n1410 & n1423;
  assign \V197(7)  = n1393 | ~n1424;
  assign n1426 = n332 & ~n825;
  assign n1427 = ~n821 & n1426;
  assign n1428 = ~n817 & n1427;
  assign n1429 = ~n814 & n1428;
  assign n1430 = ~n811 & n1429;
  assign n1431 = n406 & n920;
  assign n1432 = ~n394 & n1431;
  assign n1433 = n419 & n837;
  assign n1434 = ~n406 & n1433;
  assign n1435 = \V47(30)  & n422;
  assign n1436 = ~n419 & n1435;
  assign n1437 = \V84(6)  & ~n422;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = ~n1434 & n1438;
  assign n1440 = ~n1432 & n1439;
  assign n1441 = ~n425 & n1440;
  assign n1442 = \V133(10)  & ~n1441;
  assign n1443 = ~n825 & n1442;
  assign n1444 = ~n821 & n1443;
  assign n1445 = ~n817 & n1444;
  assign n1446 = ~n814 & n1445;
  assign n1447 = ~n811 & n1446;
  assign n1448 = ~n825 & ~n1441;
  assign n1449 = ~n821 & n1448;
  assign n1450 = ~n817 & n1449;
  assign n1451 = ~n814 & n1450;
  assign n1452 = n811 & n1451;
  assign n1453 = n814 & n1450;
  assign n1454 = n817 & n1449;
  assign n1455 = n821 & n1448;
  assign n1456 = n825 & ~n1441;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1454 & n1457;
  assign n1459 = ~n1453 & n1458;
  assign n1460 = ~n1452 & n1459;
  assign n1461 = ~n1447 & n1460;
  assign \V197(6)  = n1430 | ~n1461;
  assign n1463 = \V116(21)  & n228;
  assign n1464 = ~n825 & n1463;
  assign n1465 = ~n821 & n1464;
  assign n1466 = ~n817 & n1465;
  assign n1467 = ~n814 & n1466;
  assign n1468 = ~n811 & n1467;
  assign n1469 = \V84(6)  & n422;
  assign n1470 = n419 & n1469;
  assign n1471 = n406 & n1470;
  assign n1472 = ~n394 & n1471;
  assign n1473 = ~n419 & n1319;
  assign n1474 = \V84(21)  & ~n422;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n486 & n1475;
  assign n1477 = ~n1472 & n1476;
  assign n1478 = ~n425 & n1477;
  assign n1479 = \V133(10)  & ~n1478;
  assign n1480 = ~n825 & n1479;
  assign n1481 = ~n821 & n1480;
  assign n1482 = ~n817 & n1481;
  assign n1483 = ~n814 & n1482;
  assign n1484 = ~n811 & n1483;
  assign n1485 = ~n825 & ~n1478;
  assign n1486 = ~n821 & n1485;
  assign n1487 = ~n817 & n1486;
  assign n1488 = ~n814 & n1487;
  assign n1489 = n811 & n1488;
  assign n1490 = n814 & n1487;
  assign n1491 = n817 & n1486;
  assign n1492 = n821 & n1485;
  assign n1493 = n825 & ~n1478;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = ~n1491 & n1494;
  assign n1496 = ~n1490 & n1495;
  assign n1497 = ~n1489 & n1496;
  assign n1498 = ~n1484 & n1497;
  assign \V197(21)  = n1468 | ~n1498;
  assign n1500 = n346 & ~n825;
  assign n1501 = ~n821 & n1500;
  assign n1502 = ~n817 & n1501;
  assign n1503 = ~n814 & n1502;
  assign n1504 = ~n811 & n1503;
  assign n1505 = n406 & n1002;
  assign n1506 = ~n394 & n1505;
  assign n1507 = n419 & n1435;
  assign n1508 = ~n406 & n1507;
  assign n1509 = ~n419 & n745;
  assign n1510 = \V84(9)  & ~n422;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1508 & n1511;
  assign n1513 = ~n1506 & n1512;
  assign n1514 = ~n425 & n1513;
  assign n1515 = \V133(10)  & ~n1514;
  assign n1516 = ~n825 & n1515;
  assign n1517 = ~n821 & n1516;
  assign n1518 = ~n817 & n1517;
  assign n1519 = ~n814 & n1518;
  assign n1520 = ~n811 & n1519;
  assign n1521 = ~n825 & ~n1514;
  assign n1522 = ~n821 & n1521;
  assign n1523 = ~n817 & n1522;
  assign n1524 = ~n814 & n1523;
  assign n1525 = n811 & n1524;
  assign n1526 = n814 & n1523;
  assign n1527 = n817 & n1522;
  assign n1528 = n821 & n1521;
  assign n1529 = n825 & ~n1514;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1527 & n1530;
  assign n1532 = ~n1526 & n1531;
  assign n1533 = ~n1525 & n1532;
  assign n1534 = ~n1520 & n1533;
  assign \V197(9)  = n1504 | ~n1534;
  assign n1536 = \V116(20)  & n228;
  assign n1537 = ~n825 & n1536;
  assign n1538 = ~n821 & n1537;
  assign n1539 = ~n817 & n1538;
  assign n1540 = ~n814 & n1539;
  assign n1541 = ~n811 & n1540;
  assign n1542 = \V84(5)  & n422;
  assign n1543 = n419 & n1542;
  assign n1544 = n406 & n1543;
  assign n1545 = ~n394 & n1544;
  assign n1546 = ~n419 & n1123;
  assign n1547 = \V84(20)  & ~n422;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~n432 & n1548;
  assign n1550 = ~n1545 & n1549;
  assign n1551 = ~n425 & n1550;
  assign n1552 = \V133(10)  & ~n1551;
  assign n1553 = ~n825 & n1552;
  assign n1554 = ~n821 & n1553;
  assign n1555 = ~n817 & n1554;
  assign n1556 = ~n814 & n1555;
  assign n1557 = ~n811 & n1556;
  assign n1558 = ~n825 & ~n1551;
  assign n1559 = ~n821 & n1558;
  assign n1560 = ~n817 & n1559;
  assign n1561 = ~n814 & n1560;
  assign n1562 = n811 & n1561;
  assign n1563 = n814 & n1560;
  assign n1564 = n817 & n1559;
  assign n1565 = n821 & n1558;
  assign n1566 = n825 & ~n1551;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1564 & n1567;
  assign n1569 = ~n1563 & n1568;
  assign n1570 = ~n1562 & n1569;
  assign n1571 = ~n1557 & n1570;
  assign \V197(20)  = n1541 | ~n1571;
  assign n1573 = n360 & ~n825;
  assign n1574 = ~n821 & n1573;
  assign n1575 = ~n817 & n1574;
  assign n1576 = ~n814 & n1575;
  assign n1577 = ~n811 & n1576;
  assign n1578 = n406 & n1087;
  assign n1579 = ~n394 & n1578;
  assign n1580 = n419 & n1004;
  assign n1581 = ~n406 & n1580;
  assign n1582 = \V84(0)  & n422;
  assign n1583 = ~n419 & n1582;
  assign n1584 = \V84(8)  & ~n422;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = ~n1581 & n1585;
  assign n1587 = ~n1579 & n1586;
  assign n1588 = ~n425 & n1587;
  assign n1589 = \V133(10)  & ~n1588;
  assign n1590 = ~n825 & n1589;
  assign n1591 = ~n821 & n1590;
  assign n1592 = ~n817 & n1591;
  assign n1593 = ~n814 & n1592;
  assign n1594 = ~n811 & n1593;
  assign n1595 = ~n825 & ~n1588;
  assign n1596 = ~n821 & n1595;
  assign n1597 = ~n817 & n1596;
  assign n1598 = ~n814 & n1597;
  assign n1599 = n811 & n1598;
  assign n1600 = n814 & n1597;
  assign n1601 = n817 & n1596;
  assign n1602 = n821 & n1595;
  assign n1603 = n825 & ~n1588;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = ~n1601 & n1604;
  assign n1606 = ~n1600 & n1605;
  assign n1607 = ~n1599 & n1606;
  assign n1608 = ~n1594 & n1607;
  assign \V197(8)  = n1577 | ~n1608;
  assign n1610 = \V116(23)  & n228;
  assign n1611 = ~n825 & n1610;
  assign n1612 = ~n821 & n1611;
  assign n1613 = ~n817 & n1612;
  assign n1614 = ~n814 & n1613;
  assign n1615 = ~n811 & n1614;
  assign n1616 = \V84(8)  & n422;
  assign n1617 = n419 & n1616;
  assign n1618 = n406 & n1617;
  assign n1619 = ~n394 & n1618;
  assign n1620 = ~n406 & n1124;
  assign n1621 = ~n419 & n1166;
  assign n1622 = \V84(23)  & ~n422;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n1620 & n1623;
  assign n1625 = ~n1619 & n1624;
  assign n1626 = ~n425 & n1625;
  assign n1627 = \V133(10)  & ~n1626;
  assign n1628 = ~n825 & n1627;
  assign n1629 = ~n821 & n1628;
  assign n1630 = ~n817 & n1629;
  assign n1631 = ~n814 & n1630;
  assign n1632 = ~n811 & n1631;
  assign n1633 = ~n825 & ~n1626;
  assign n1634 = ~n821 & n1633;
  assign n1635 = ~n817 & n1634;
  assign n1636 = ~n814 & n1635;
  assign n1637 = n811 & n1636;
  assign n1638 = n814 & n1635;
  assign n1639 = n817 & n1634;
  assign n1640 = n821 & n1633;
  assign n1641 = n825 & ~n1626;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = ~n1639 & n1642;
  assign n1644 = ~n1638 & n1643;
  assign n1645 = ~n1637 & n1644;
  assign n1646 = ~n1632 & n1645;
  assign \V197(23)  = n1615 | ~n1646;
  assign n1648 = \V116(22)  & n228;
  assign n1649 = ~n825 & n1648;
  assign n1650 = ~n821 & n1649;
  assign n1651 = ~n817 & n1650;
  assign n1652 = ~n814 & n1651;
  assign n1653 = ~n811 & n1652;
  assign n1654 = \V84(7)  & n422;
  assign n1655 = n419 & n1654;
  assign n1656 = n406 & n1655;
  assign n1657 = ~n394 & n1656;
  assign n1658 = ~n419 & n1244;
  assign n1659 = \V84(22)  & ~n422;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n460 & n1660;
  assign n1662 = ~n1657 & n1661;
  assign n1663 = ~n425 & n1662;
  assign n1664 = \V133(10)  & ~n1663;
  assign n1665 = ~n825 & n1664;
  assign n1666 = ~n821 & n1665;
  assign n1667 = ~n817 & n1666;
  assign n1668 = ~n814 & n1667;
  assign n1669 = ~n811 & n1668;
  assign n1670 = ~n825 & ~n1663;
  assign n1671 = ~n821 & n1670;
  assign n1672 = ~n817 & n1671;
  assign n1673 = ~n814 & n1672;
  assign n1674 = n811 & n1673;
  assign n1675 = n814 & n1672;
  assign n1676 = n817 & n1671;
  assign n1677 = n821 & n1670;
  assign n1678 = n825 & ~n1663;
  assign n1679 = ~n1677 & ~n1678;
  assign n1680 = ~n1676 & n1679;
  assign n1681 = ~n1675 & n1680;
  assign n1682 = ~n1674 & n1681;
  assign n1683 = ~n1669 & n1682;
  assign \V197(22)  = n1653 | ~n1683;
  assign n1685 = \V116(25)  & n228;
  assign n1686 = ~n825 & n1685;
  assign n1687 = ~n821 & n1686;
  assign n1688 = ~n817 & n1687;
  assign n1689 = ~n814 & n1688;
  assign n1690 = ~n811 & n1689;
  assign n1691 = n406 & n485;
  assign n1692 = ~n394 & n1691;
  assign n1693 = ~n406 & n1245;
  assign n1694 = ~n419 & n1323;
  assign n1695 = \V84(25)  & ~n422;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = ~n1693 & n1696;
  assign n1698 = ~n1692 & n1697;
  assign n1699 = ~n425 & n1698;
  assign n1700 = \V133(10)  & ~n1699;
  assign n1701 = ~n825 & n1700;
  assign n1702 = ~n821 & n1701;
  assign n1703 = ~n817 & n1702;
  assign n1704 = ~n814 & n1703;
  assign n1705 = ~n811 & n1704;
  assign n1706 = ~n825 & ~n1699;
  assign n1707 = ~n821 & n1706;
  assign n1708 = ~n817 & n1707;
  assign n1709 = ~n814 & n1708;
  assign n1710 = n811 & n1709;
  assign n1711 = n814 & n1708;
  assign n1712 = n817 & n1707;
  assign n1713 = n821 & n1706;
  assign n1714 = n825 & ~n1699;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1712 & n1715;
  assign n1717 = ~n1711 & n1716;
  assign n1718 = ~n1710 & n1717;
  assign n1719 = ~n1705 & n1718;
  assign \V197(25)  = n1690 | ~n1719;
  assign n1721 = \V116(24)  & n228;
  assign n1722 = ~n825 & n1721;
  assign n1723 = ~n821 & n1722;
  assign n1724 = ~n817 & n1723;
  assign n1725 = ~n814 & n1724;
  assign n1726 = ~n811 & n1725;
  assign n1727 = n406 & n431;
  assign n1728 = ~n394 & n1727;
  assign n1729 = ~n406 & n1320;
  assign n1730 = ~n419 & n1127;
  assign n1731 = \V84(24)  & ~n422;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1729 & n1732;
  assign n1734 = ~n1728 & n1733;
  assign n1735 = ~n425 & n1734;
  assign n1736 = \V133(10)  & ~n1735;
  assign n1737 = ~n825 & n1736;
  assign n1738 = ~n821 & n1737;
  assign n1739 = ~n817 & n1738;
  assign n1740 = ~n814 & n1739;
  assign n1741 = ~n811 & n1740;
  assign n1742 = ~n825 & ~n1735;
  assign n1743 = ~n821 & n1742;
  assign n1744 = ~n817 & n1743;
  assign n1745 = ~n814 & n1744;
  assign n1746 = n811 & n1745;
  assign n1747 = n814 & n1744;
  assign n1748 = n817 & n1743;
  assign n1749 = n821 & n1742;
  assign n1750 = n825 & ~n1735;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = ~n1748 & n1751;
  assign n1753 = ~n1747 & n1752;
  assign n1754 = ~n1746 & n1753;
  assign n1755 = ~n1741 & n1754;
  assign \V197(24)  = n1726 | ~n1755;
  assign n1757 = ~\V133(8)  & n377;
  assign n1758 = ~\V133(9)  & n1757;
  assign n1759 = ~\V133(10)  & ~n1758;
  assign n1760 = ~n228 & n1759;
  assign n1761 = ~n375 & n1760;
  assign n1762 = n685 & n1761;
  assign n1763 = \V133(10)  & \V119(0) ;
  assign n1764 = ~n1758 & n1763;
  assign n1765 = ~n228 & n1764;
  assign n1766 = ~n375 & n1765;
  assign n1767 = ~n685 & n1761;
  assign n1768 = n683 & n1767;
  assign n1769 = ~n683 & n1767;
  assign n1770 = \V121(16)  & n1758;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = ~n1768 & n1771;
  assign n1773 = ~n1766 & n1772;
  assign \V213(0)  = n1762 | ~n1773;
  assign n1775 = \V116(17)  & n228;
  assign n1776 = ~n825 & n1775;
  assign n1777 = ~n821 & n1776;
  assign n1778 = ~n817 & n1777;
  assign n1779 = ~n814 & n1778;
  assign n1780 = ~n811 & n1779;
  assign n1781 = n406 & n708;
  assign n1782 = ~n394 & n1781;
  assign n1783 = ~n406 & n1470;
  assign n1784 = ~n419 & n430;
  assign n1785 = \V84(17)  & ~n422;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1783 & n1786;
  assign n1788 = ~n1782 & n1787;
  assign n1789 = ~n425 & n1788;
  assign n1790 = \V133(10)  & ~n1789;
  assign n1791 = ~n825 & n1790;
  assign n1792 = ~n821 & n1791;
  assign n1793 = ~n817 & n1792;
  assign n1794 = ~n814 & n1793;
  assign n1795 = ~n811 & n1794;
  assign n1796 = ~n825 & ~n1789;
  assign n1797 = ~n821 & n1796;
  assign n1798 = ~n817 & n1797;
  assign n1799 = ~n814 & n1798;
  assign n1800 = n811 & n1799;
  assign n1801 = n814 & n1798;
  assign n1802 = n817 & n1797;
  assign n1803 = n821 & n1796;
  assign n1804 = n825 & ~n1789;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = ~n1802 & n1805;
  assign n1807 = ~n1801 & n1806;
  assign n1808 = ~n1800 & n1807;
  assign n1809 = ~n1795 & n1808;
  assign \V197(17)  = n1780 | ~n1809;
  assign n1811 = \V116(16)  & n228;
  assign n1812 = ~n825 & n1811;
  assign n1813 = ~n821 & n1812;
  assign n1814 = ~n817 & n1813;
  assign n1815 = ~n814 & n1814;
  assign n1816 = ~n811 & n1815;
  assign n1817 = n406 & n746;
  assign n1818 = ~n394 & n1817;
  assign n1819 = ~n406 & n1543;
  assign n1820 = ~n419 & n1616;
  assign n1821 = \V84(16)  & ~n422;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1819 & n1822;
  assign n1824 = ~n1818 & n1823;
  assign n1825 = ~n425 & n1824;
  assign n1826 = \V133(10)  & ~n1825;
  assign n1827 = ~n825 & n1826;
  assign n1828 = ~n821 & n1827;
  assign n1829 = ~n817 & n1828;
  assign n1830 = ~n814 & n1829;
  assign n1831 = ~n811 & n1830;
  assign n1832 = ~n825 & ~n1825;
  assign n1833 = ~n821 & n1832;
  assign n1834 = ~n817 & n1833;
  assign n1835 = ~n814 & n1834;
  assign n1836 = n811 & n1835;
  assign n1837 = n814 & n1834;
  assign n1838 = n817 & n1833;
  assign n1839 = n821 & n1832;
  assign n1840 = n825 & ~n1825;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~n1838 & n1841;
  assign n1843 = ~n1837 & n1842;
  assign n1844 = ~n1836 & n1843;
  assign n1845 = ~n1831 & n1844;
  assign \V197(16)  = n1816 | ~n1845;
  assign n1847 = \V116(19)  & n228;
  assign n1848 = ~n825 & n1847;
  assign n1849 = ~n821 & n1848;
  assign n1850 = ~n817 & n1849;
  assign n1851 = ~n814 & n1850;
  assign n1852 = ~n811 & n1851;
  assign n1853 = \V84(4)  & n422;
  assign n1854 = n419 & n1853;
  assign n1855 = n406 & n1854;
  assign n1856 = ~n394 & n1855;
  assign n1857 = ~n406 & n1617;
  assign n1858 = ~n419 & n458;
  assign n1859 = \V84(19)  & ~n422;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & n1860;
  assign n1862 = ~n1856 & n1861;
  assign n1863 = ~n425 & n1862;
  assign n1864 = \V133(10)  & ~n1863;
  assign n1865 = ~n825 & n1864;
  assign n1866 = ~n821 & n1865;
  assign n1867 = ~n817 & n1866;
  assign n1868 = ~n814 & n1867;
  assign n1869 = ~n811 & n1868;
  assign n1870 = ~n825 & ~n1863;
  assign n1871 = ~n821 & n1870;
  assign n1872 = ~n817 & n1871;
  assign n1873 = ~n814 & n1872;
  assign n1874 = n811 & n1873;
  assign n1875 = n814 & n1872;
  assign n1876 = n817 & n1871;
  assign n1877 = n821 & n1870;
  assign n1878 = n825 & ~n1863;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = ~n1876 & n1879;
  assign n1881 = ~n1875 & n1880;
  assign n1882 = ~n1874 & n1881;
  assign n1883 = ~n1869 & n1882;
  assign \V197(19)  = n1852 | ~n1883;
  assign n1885 = \V116(18)  & n228;
  assign n1886 = ~n825 & n1885;
  assign n1887 = ~n821 & n1886;
  assign n1888 = ~n817 & n1887;
  assign n1889 = ~n814 & n1888;
  assign n1890 = ~n811 & n1889;
  assign n1891 = \V84(3)  & n422;
  assign n1892 = n419 & n1891;
  assign n1893 = n406 & n1892;
  assign n1894 = ~n394 & n1893;
  assign n1895 = ~n406 & n1655;
  assign n1896 = ~n419 & n484;
  assign n1897 = \V84(18)  & ~n422;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1895 & n1898;
  assign n1900 = ~n1894 & n1899;
  assign n1901 = ~n425 & n1900;
  assign n1902 = \V133(10)  & ~n1901;
  assign n1903 = ~n825 & n1902;
  assign n1904 = ~n821 & n1903;
  assign n1905 = ~n817 & n1904;
  assign n1906 = ~n814 & n1905;
  assign n1907 = ~n811 & n1906;
  assign n1908 = ~n825 & ~n1901;
  assign n1909 = ~n821 & n1908;
  assign n1910 = ~n817 & n1909;
  assign n1911 = ~n814 & n1910;
  assign n1912 = n811 & n1911;
  assign n1913 = n814 & n1910;
  assign n1914 = n817 & n1909;
  assign n1915 = n821 & n1908;
  assign n1916 = n825 & ~n1901;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n1914 & n1917;
  assign n1919 = ~n1913 & n1918;
  assign n1920 = ~n1912 & n1919;
  assign n1921 = ~n1907 & n1920;
  assign \V197(18)  = n1890 | ~n1921;
  assign n1923 = n451 & ~n825;
  assign n1924 = ~n821 & n1923;
  assign n1925 = ~n817 & n1924;
  assign n1926 = ~n814 & n1925;
  assign n1927 = ~n811 & n1926;
  assign n1928 = n406 & n1396;
  assign n1929 = ~n394 & n1928;
  assign n1930 = n419 & n1582;
  assign n1931 = ~n406 & n1930;
  assign n1932 = ~n419 & n1891;
  assign n1933 = \V84(11)  & ~n422;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = ~n1931 & n1934;
  assign n1936 = ~n1929 & n1935;
  assign n1937 = ~n425 & n1936;
  assign n1938 = \V133(10)  & ~n1937;
  assign n1939 = ~n825 & n1938;
  assign n1940 = ~n821 & n1939;
  assign n1941 = ~n817 & n1940;
  assign n1942 = ~n814 & n1941;
  assign n1943 = ~n811 & n1942;
  assign n1944 = ~n825 & ~n1937;
  assign n1945 = ~n821 & n1944;
  assign n1946 = ~n817 & n1945;
  assign n1947 = ~n814 & n1946;
  assign n1948 = n811 & n1947;
  assign n1949 = n814 & n1946;
  assign n1950 = n817 & n1945;
  assign n1951 = n821 & n1944;
  assign n1952 = n825 & ~n1937;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = ~n1950 & n1953;
  assign n1955 = ~n1949 & n1954;
  assign n1956 = ~n1948 & n1955;
  assign n1957 = ~n1943 & n1956;
  assign \V197(11)  = n1927 | ~n1957;
  assign n1959 = n477 & ~n825;
  assign n1960 = ~n821 & n1959;
  assign n1961 = ~n817 & n1960;
  assign n1962 = ~n814 & n1961;
  assign n1963 = ~n811 & n1962;
  assign n1964 = n406 & n1433;
  assign n1965 = ~n394 & n1964;
  assign n1966 = n419 & n1398;
  assign n1967 = ~n406 & n1966;
  assign n1968 = ~n419 & n707;
  assign n1969 = \V84(10)  & ~n422;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n1967 & n1970;
  assign n1972 = ~n1965 & n1971;
  assign n1973 = ~n425 & n1972;
  assign n1974 = \V133(10)  & ~n1973;
  assign n1975 = ~n825 & n1974;
  assign n1976 = ~n821 & n1975;
  assign n1977 = ~n817 & n1976;
  assign n1978 = ~n814 & n1977;
  assign n1979 = ~n811 & n1978;
  assign n1980 = ~n825 & ~n1973;
  assign n1981 = ~n821 & n1980;
  assign n1982 = ~n817 & n1981;
  assign n1983 = ~n814 & n1982;
  assign n1984 = n811 & n1983;
  assign n1985 = n814 & n1982;
  assign n1986 = n817 & n1981;
  assign n1987 = n821 & n1980;
  assign n1988 = n825 & ~n1973;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1986 & n1989;
  assign n1991 = ~n1985 & n1990;
  assign n1992 = ~n1984 & n1991;
  assign n1993 = ~n1979 & n1992;
  assign \V197(10)  = n1963 | ~n1993;
  assign n1995 = \V116(13)  & n228;
  assign n1996 = ~n825 & n1995;
  assign n1997 = ~n821 & n1996;
  assign n1998 = ~n817 & n1997;
  assign n1999 = ~n814 & n1998;
  assign n2000 = ~n811 & n1999;
  assign n2001 = n406 & n1507;
  assign n2002 = ~n394 & n2001;
  assign n2003 = ~n419 & n1542;
  assign n2004 = \V84(13)  & ~n422;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n709 & n2005;
  assign n2007 = ~n2002 & n2006;
  assign n2008 = ~n425 & n2007;
  assign n2009 = \V133(10)  & ~n2008;
  assign n2010 = ~n825 & n2009;
  assign n2011 = ~n821 & n2010;
  assign n2012 = ~n817 & n2011;
  assign n2013 = ~n814 & n2012;
  assign n2014 = ~n811 & n2013;
  assign n2015 = ~n825 & ~n2008;
  assign n2016 = ~n821 & n2015;
  assign n2017 = ~n817 & n2016;
  assign n2018 = ~n814 & n2017;
  assign n2019 = n811 & n2018;
  assign n2020 = n814 & n2017;
  assign n2021 = n817 & n2016;
  assign n2022 = n821 & n2015;
  assign n2023 = n825 & ~n2008;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~n2021 & n2024;
  assign n2026 = ~n2020 & n2025;
  assign n2027 = ~n2019 & n2026;
  assign n2028 = ~n2014 & n2027;
  assign \V197(13)  = n2000 | ~n2028;
  assign n2030 = \V116(12)  & n228;
  assign n2031 = ~n825 & n2030;
  assign n2032 = ~n821 & n2031;
  assign n2033 = ~n817 & n2032;
  assign n2034 = ~n814 & n2033;
  assign n2035 = ~n811 & n2034;
  assign n2036 = n406 & n1580;
  assign n2037 = ~n394 & n2036;
  assign n2038 = ~n419 & n1853;
  assign n2039 = \V84(12)  & ~n422;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~n747 & n2040;
  assign n2042 = ~n2037 & n2041;
  assign n2043 = ~n425 & n2042;
  assign n2044 = \V133(10)  & ~n2043;
  assign n2045 = ~n825 & n2044;
  assign n2046 = ~n821 & n2045;
  assign n2047 = ~n817 & n2046;
  assign n2048 = ~n814 & n2047;
  assign n2049 = ~n811 & n2048;
  assign n2050 = ~n825 & ~n2043;
  assign n2051 = ~n821 & n2050;
  assign n2052 = ~n817 & n2051;
  assign n2053 = ~n814 & n2052;
  assign n2054 = n811 & n2053;
  assign n2055 = n814 & n2052;
  assign n2056 = n817 & n2051;
  assign n2057 = n821 & n2050;
  assign n2058 = n825 & ~n2043;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~n2056 & n2059;
  assign n2061 = ~n2055 & n2060;
  assign n2062 = ~n2054 & n2061;
  assign n2063 = ~n2049 & n2062;
  assign \V197(12)  = n2035 | ~n2063;
  assign n2065 = \V116(15)  & n228;
  assign n2066 = ~n825 & n2065;
  assign n2067 = ~n821 & n2066;
  assign n2068 = ~n817 & n2067;
  assign n2069 = ~n814 & n2068;
  assign n2070 = ~n811 & n2069;
  assign n2071 = n406 & n1930;
  assign n2072 = ~n394 & n2071;
  assign n2073 = ~n406 & n1854;
  assign n2074 = ~n419 & n1654;
  assign n2075 = \V84(15)  & ~n422;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = ~n2073 & n2076;
  assign n2078 = ~n2072 & n2077;
  assign n2079 = ~n425 & n2078;
  assign n2080 = \V133(10)  & ~n2079;
  assign n2081 = ~n825 & n2080;
  assign n2082 = ~n821 & n2081;
  assign n2083 = ~n817 & n2082;
  assign n2084 = ~n814 & n2083;
  assign n2085 = ~n811 & n2084;
  assign n2086 = ~n825 & ~n2079;
  assign n2087 = ~n821 & n2086;
  assign n2088 = ~n817 & n2087;
  assign n2089 = ~n814 & n2088;
  assign n2090 = n811 & n2089;
  assign n2091 = n814 & n2088;
  assign n2092 = n817 & n2087;
  assign n2093 = n821 & n2086;
  assign n2094 = n825 & ~n2079;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n2092 & n2095;
  assign n2097 = ~n2091 & n2096;
  assign n2098 = ~n2090 & n2097;
  assign n2099 = ~n2085 & n2098;
  assign \V197(15)  = n2070 | ~n2099;
  assign n2101 = \V116(14)  & n228;
  assign n2102 = ~n825 & n2101;
  assign n2103 = ~n821 & n2102;
  assign n2104 = ~n817 & n2103;
  assign n2105 = ~n814 & n2104;
  assign n2106 = ~n811 & n2105;
  assign n2107 = n406 & n1966;
  assign n2108 = ~n394 & n2107;
  assign n2109 = ~n406 & n1892;
  assign n2110 = ~n419 & n1469;
  assign n2111 = \V84(14)  & ~n422;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~n2109 & n2112;
  assign n2114 = ~n2108 & n2113;
  assign n2115 = ~n425 & n2114;
  assign n2116 = \V133(10)  & ~n2115;
  assign n2117 = ~n825 & n2116;
  assign n2118 = ~n821 & n2117;
  assign n2119 = ~n817 & n2118;
  assign n2120 = ~n814 & n2119;
  assign n2121 = ~n811 & n2120;
  assign n2122 = ~n825 & ~n2115;
  assign n2123 = ~n821 & n2122;
  assign n2124 = ~n817 & n2123;
  assign n2125 = ~n814 & n2124;
  assign n2126 = n811 & n2125;
  assign n2127 = n814 & n2124;
  assign n2128 = n817 & n2123;
  assign n2129 = n821 & n2122;
  assign n2130 = n825 & ~n2115;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = ~n2128 & n2131;
  assign n2133 = ~n2127 & n2132;
  assign n2134 = ~n2126 & n2133;
  assign n2135 = ~n2121 & n2134;
  assign \V197(14)  = n2106 | ~n2135;
  assign n2137 = n332 & ~n450;
  assign n2138 = ~n386 & n2137;
  assign n2139 = \V15(5)  & n422;
  assign n2140 = n419 & n2139;
  assign n2141 = n406 & n2140;
  assign n2142 = ~n394 & n2141;
  assign n2143 = \V47(6)  & ~n422;
  assign n2144 = ~n425 & ~n2143;
  assign n2145 = ~n1783 & n2144;
  assign n2146 = ~n2142 & n2145;
  assign n2147 = \V133(10)  & ~n2146;
  assign n2148 = ~n450 & n2147;
  assign n2149 = ~n386 & n2148;
  assign n2150 = ~n450 & ~n2146;
  assign n2151 = n386 & n2150;
  assign n2152 = n450 & ~n2146;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2149 & n2153;
  assign \V142(3)  = n2138 | ~n2154;
  assign n2156 = n261 & ~n450;
  assign n2157 = ~n386 & n2156;
  assign n2158 = \V15(4)  & n422;
  assign n2159 = n419 & n2158;
  assign n2160 = n406 & n2159;
  assign n2161 = ~n394 & n2160;
  assign n2162 = \V47(5)  & ~n422;
  assign n2163 = ~n425 & ~n2162;
  assign n2164 = ~n1819 & n2163;
  assign n2165 = ~n2161 & n2164;
  assign n2166 = \V133(10)  & ~n2165;
  assign n2167 = ~n450 & n2166;
  assign n2168 = ~n386 & n2167;
  assign n2169 = ~n450 & ~n2165;
  assign n2170 = n386 & n2169;
  assign n2171 = n450 & ~n2165;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n2168 & n2172;
  assign \V142(2)  = n2157 | ~n2173;
  assign n2175 = n360 & ~n450;
  assign n2176 = ~n386 & n2175;
  assign n2177 = \V15(7)  & n422;
  assign n2178 = n419 & n2177;
  assign n2179 = n406 & n2178;
  assign n2180 = ~n394 & n2179;
  assign n2181 = \V47(0)  & n422;
  assign n2182 = ~n419 & n2181;
  assign n2183 = \V47(8)  & ~n422;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~n1857 & n2184;
  assign n2186 = ~n2180 & n2185;
  assign n2187 = ~n425 & n2186;
  assign n2188 = \V133(10)  & ~n2187;
  assign n2189 = ~n450 & n2188;
  assign n2190 = ~n386 & n2189;
  assign n2191 = ~n450 & ~n2187;
  assign n2192 = n386 & n2191;
  assign n2193 = n450 & ~n2187;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = ~n2190 & n2194;
  assign \V142(5)  = n2176 | ~n2195;
  assign n2197 = n318 & ~n450;
  assign n2198 = ~n386 & n2197;
  assign n2199 = \V15(6)  & n422;
  assign n2200 = n419 & n2199;
  assign n2201 = n406 & n2200;
  assign n2202 = ~n394 & n2201;
  assign n2203 = \V47(7)  & ~n422;
  assign n2204 = ~n425 & ~n2203;
  assign n2205 = ~n1895 & n2204;
  assign n2206 = ~n2202 & n2205;
  assign n2207 = \V133(10)  & ~n2206;
  assign n2208 = ~n450 & n2207;
  assign n2209 = ~n386 & n2208;
  assign n2210 = ~n450 & ~n2206;
  assign n2211 = n386 & n2210;
  assign n2212 = n450 & ~n2206;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = ~n2209 & n2213;
  assign \V142(4)  = n2198 | ~n2214;
  assign n2216 = \V116(31)  & n228;
  assign n2217 = ~n825 & n2216;
  assign n2218 = ~n821 & n2217;
  assign n2219 = ~n817 & n2218;
  assign n2220 = ~n814 & n2219;
  assign n2221 = ~n811 & n2220;
  assign n2222 = n406 & n1128;
  assign n2223 = ~n394 & n2222;
  assign n2224 = n419 & n1326;
  assign n2225 = ~n406 & n2224;
  assign n2226 = \V84(23)  & n422;
  assign n2227 = ~n419 & n2226;
  assign n2228 = \V84(31)  & ~n422;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2225 & n2229;
  assign n2231 = ~n2223 & n2230;
  assign n2232 = ~n425 & n2231;
  assign n2233 = \V133(10)  & ~n2232;
  assign n2234 = ~n825 & n2233;
  assign n2235 = ~n821 & n2234;
  assign n2236 = ~n817 & n2235;
  assign n2237 = ~n814 & n2236;
  assign n2238 = ~n811 & n2237;
  assign n2239 = ~n825 & ~n2232;
  assign n2240 = ~n821 & n2239;
  assign n2241 = ~n817 & n2240;
  assign n2242 = ~n814 & n2241;
  assign n2243 = n811 & n2242;
  assign n2244 = n814 & n2241;
  assign n2245 = n817 & n2240;
  assign n2246 = n821 & n2239;
  assign n2247 = n825 & ~n2232;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = ~n2245 & n2248;
  assign n2250 = ~n2244 & n2249;
  assign n2251 = ~n2243 & n2250;
  assign n2252 = ~n2238 & n2251;
  assign \V197(31)  = n2221 | ~n2252;
  assign n2254 = n275 & ~n450;
  assign n2255 = ~n386 & n2254;
  assign n2256 = \V15(3)  & n422;
  assign n2257 = n419 & n2256;
  assign n2258 = n406 & n2257;
  assign n2259 = ~n394 & n2258;
  assign n2260 = \V47(4)  & ~n422;
  assign n2261 = ~n425 & ~n2260;
  assign n2262 = ~n2073 & n2261;
  assign n2263 = ~n2259 & n2262;
  assign n2264 = \V133(10)  & ~n2263;
  assign n2265 = ~n450 & n2264;
  assign n2266 = ~n386 & n2265;
  assign n2267 = ~n450 & ~n2263;
  assign n2268 = n386 & n2267;
  assign n2269 = n450 & ~n2263;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = ~n2266 & n2270;
  assign \V142(1)  = n2255 | ~n2271;
  assign n2273 = \V116(30)  & n228;
  assign n2274 = ~n825 & n2273;
  assign n2275 = ~n821 & n2274;
  assign n2276 = ~n817 & n2275;
  assign n2277 = ~n814 & n2276;
  assign n2278 = ~n811 & n2277;
  assign n2279 = n406 & n1167;
  assign n2280 = ~n394 & n2279;
  assign n2281 = n419 & n1130;
  assign n2282 = ~n406 & n2281;
  assign n2283 = \V84(22)  & n422;
  assign n2284 = ~n419 & n2283;
  assign n2285 = \V84(30)  & ~n422;
  assign n2286 = ~n2284 & ~n2285;
  assign n2287 = ~n2282 & n2286;
  assign n2288 = ~n2280 & n2287;
  assign n2289 = ~n425 & n2288;
  assign n2290 = \V133(10)  & ~n2289;
  assign n2291 = ~n825 & n2290;
  assign n2292 = ~n821 & n2291;
  assign n2293 = ~n817 & n2292;
  assign n2294 = ~n814 & n2293;
  assign n2295 = ~n811 & n2294;
  assign n2296 = ~n825 & ~n2289;
  assign n2297 = ~n821 & n2296;
  assign n2298 = ~n817 & n2297;
  assign n2299 = ~n814 & n2298;
  assign n2300 = n811 & n2299;
  assign n2301 = n814 & n2298;
  assign n2302 = n817 & n2297;
  assign n2303 = n821 & n2296;
  assign n2304 = n825 & ~n2289;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n2302 & n2305;
  assign n2307 = ~n2301 & n2306;
  assign n2308 = ~n2300 & n2307;
  assign n2309 = ~n2295 & n2308;
  assign \V197(30)  = n2278 | ~n2309;
  assign n2311 = n229 & ~n450;
  assign n2312 = ~n386 & n2311;
  assign n2313 = \V15(2)  & n422;
  assign n2314 = n419 & n2313;
  assign n2315 = n406 & n2314;
  assign n2316 = ~n394 & n2315;
  assign n2317 = \V47(3)  & ~n422;
  assign n2318 = ~n425 & ~n2317;
  assign n2319 = ~n2109 & n2318;
  assign n2320 = ~n2316 & n2319;
  assign n2321 = \V133(10)  & ~n2320;
  assign n2322 = ~n450 & n2321;
  assign n2323 = ~n386 & n2322;
  assign n2324 = ~n450 & ~n2320;
  assign n2325 = n386 & n2324;
  assign n2326 = n450 & ~n2320;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = ~n2323 & n2327;
  assign \V142(0)  = n2312 | ~n2328;
  assign n2330 = \V84(20)  & n511;
  assign n2331 = ~\V133(9)  & n2330;
  assign n2332 = ~\V133(4)  & n2331;
  assign n2333 = ~n510 & n2332;
  assign n2334 = ~n507 & n2333;
  assign n2335 = ~n504 & n2334;
  assign n2336 = ~n386 & n2335;
  assign n2337 = ~n228 & n2336;
  assign n2338 = ~\V133(10)  & \V116(20) ;
  assign n2339 = ~n510 & n2338;
  assign n2340 = ~n507 & n2339;
  assign n2341 = ~n504 & n2340;
  assign n2342 = ~n386 & n2341;
  assign n2343 = n228 & n2342;
  assign n2344 = n419 & n623;
  assign n2345 = n406 & n2344;
  assign n2346 = ~n394 & n2345;
  assign n2347 = \V47(9)  & n422;
  assign n2348 = n419 & n2347;
  assign n2349 = ~n406 & n2348;
  assign n2350 = ~n419 & n879;
  assign n2351 = \V47(20)  & ~n422;
  assign n2352 = ~n2350 & ~n2351;
  assign n2353 = ~n2349 & n2352;
  assign n2354 = ~n2346 & n2353;
  assign n2355 = ~n425 & n2354;
  assign n2356 = \V133(10)  & ~n2355;
  assign n2357 = ~n510 & n2356;
  assign n2358 = ~n507 & n2357;
  assign n2359 = ~n504 & n2358;
  assign n2360 = ~n386 & n2359;
  assign n2361 = ~n510 & ~n2355;
  assign n2362 = ~n507 & n2361;
  assign n2363 = ~n504 & n2362;
  assign n2364 = n386 & n2363;
  assign n2365 = n504 & n2362;
  assign n2366 = n507 & n2361;
  assign n2367 = n510 & ~n2355;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n2365 & n2368;
  assign n2370 = ~n2364 & n2369;
  assign n2371 = ~n2360 & n2370;
  assign n2372 = ~n2343 & n2371;
  assign \V165(3)  = n2337 | ~n2372;
  assign n2374 = ~n227 & n451;
  assign n2375 = ~n223 & n2374;
  assign n2376 = ~n221 & n2375;
  assign n2377 = \V84(28)  & \V133(10) ;
  assign n2378 = ~n227 & n2377;
  assign n2379 = ~n223 & n2378;
  assign n2380 = \V84(28)  & ~n227;
  assign n2381 = n223 & n2380;
  assign n2382 = \V84(28)  & n227;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2379 & n2383;
  assign n2385 = ~n235 & n2384;
  assign \V212(11)  = n2376 | ~n2385;
  assign n2387 = \V84(19)  & n511;
  assign n2388 = ~\V133(9)  & n2387;
  assign n2389 = ~\V133(4)  & n2388;
  assign n2390 = ~n510 & n2389;
  assign n2391 = ~n507 & n2390;
  assign n2392 = ~n504 & n2391;
  assign n2393 = ~n386 & n2392;
  assign n2394 = ~n228 & n2393;
  assign n2395 = ~\V133(10)  & \V116(19) ;
  assign n2396 = ~n510 & n2395;
  assign n2397 = ~n507 & n2396;
  assign n2398 = ~n504 & n2397;
  assign n2399 = ~n386 & n2398;
  assign n2400 = n228 & n2399;
  assign n2401 = n406 & n531;
  assign n2402 = ~n394 & n2401;
  assign n2403 = \V47(8)  & n422;
  assign n2404 = n419 & n2403;
  assign n2405 = ~n406 & n2404;
  assign n2406 = \V47(11)  & n422;
  assign n2407 = ~n419 & n2406;
  assign n2408 = \V47(19)  & ~n422;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~n2405 & n2409;
  assign n2411 = ~n2402 & n2410;
  assign n2412 = ~n425 & n2411;
  assign n2413 = \V133(10)  & ~n2412;
  assign n2414 = ~n510 & n2413;
  assign n2415 = ~n507 & n2414;
  assign n2416 = ~n504 & n2415;
  assign n2417 = ~n386 & n2416;
  assign n2418 = ~n510 & ~n2412;
  assign n2419 = ~n507 & n2418;
  assign n2420 = ~n504 & n2419;
  assign n2421 = n386 & n2420;
  assign n2422 = n504 & n2419;
  assign n2423 = n507 & n2418;
  assign n2424 = n510 & ~n2412;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~n2422 & n2425;
  assign n2427 = ~n2421 & n2426;
  assign n2428 = ~n2417 & n2427;
  assign n2429 = ~n2400 & n2428;
  assign \V165(2)  = n2394 | ~n2429;
  assign n2431 = ~n227 & n477;
  assign n2432 = ~n223 & n2431;
  assign n2433 = ~n221 & n2432;
  assign n2434 = \V84(27)  & \V133(10) ;
  assign n2435 = ~n227 & n2434;
  assign n2436 = ~n223 & n2435;
  assign n2437 = \V84(27)  & ~n227;
  assign n2438 = n223 & n2437;
  assign n2439 = \V84(27)  & n227;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = ~n2436 & n2440;
  assign n2442 = ~n235 & n2441;
  assign \V212(10)  = n2433 | ~n2442;
  assign n2444 = \V84(22)  & n511;
  assign n2445 = ~\V133(9)  & n2444;
  assign n2446 = ~\V133(4)  & n2445;
  assign n2447 = ~n510 & n2446;
  assign n2448 = ~n507 & n2447;
  assign n2449 = ~n504 & n2448;
  assign n2450 = ~n386 & n2449;
  assign n2451 = ~n228 & n2450;
  assign n2452 = ~\V133(10)  & \V116(22) ;
  assign n2453 = ~n510 & n2452;
  assign n2454 = ~n507 & n2453;
  assign n2455 = ~n504 & n2454;
  assign n2456 = ~n386 & n2455;
  assign n2457 = n228 & n2456;
  assign n2458 = n419 & n533;
  assign n2459 = n406 & n2458;
  assign n2460 = ~n394 & n2459;
  assign n2461 = n419 & n2406;
  assign n2462 = ~n406 & n2461;
  assign n2463 = ~n419 & n1046;
  assign n2464 = \V47(22)  & ~n422;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~n2462 & n2465;
  assign n2467 = ~n2460 & n2466;
  assign n2468 = ~n425 & n2467;
  assign n2469 = \V133(10)  & ~n2468;
  assign n2470 = ~n510 & n2469;
  assign n2471 = ~n507 & n2470;
  assign n2472 = ~n504 & n2471;
  assign n2473 = ~n386 & n2472;
  assign n2474 = ~n510 & ~n2468;
  assign n2475 = ~n507 & n2474;
  assign n2476 = ~n504 & n2475;
  assign n2477 = n386 & n2476;
  assign n2478 = n504 & n2475;
  assign n2479 = n507 & n2474;
  assign n2480 = n510 & ~n2468;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = ~n2478 & n2481;
  assign n2483 = ~n2477 & n2482;
  assign n2484 = ~n2473 & n2483;
  assign n2485 = ~n2457 & n2484;
  assign \V165(5)  = n2451 | ~n2485;
  assign n2487 = ~n227 & n1995;
  assign n2488 = ~n223 & n2487;
  assign n2489 = ~n221 & n2488;
  assign n2490 = \V84(30)  & \V133(10) ;
  assign n2491 = ~n227 & n2490;
  assign n2492 = ~n223 & n2491;
  assign n2493 = \V84(30)  & ~n227;
  assign n2494 = n223 & n2493;
  assign n2495 = \V84(30)  & n227;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = ~n2492 & n2496;
  assign n2498 = ~n235 & n2497;
  assign \V212(13)  = n2489 | ~n2498;
  assign n2500 = \V84(21)  & n511;
  assign n2501 = ~\V133(9)  & n2500;
  assign n2502 = ~\V133(4)  & n2501;
  assign n2503 = ~n510 & n2502;
  assign n2504 = ~n507 & n2503;
  assign n2505 = ~n504 & n2504;
  assign n2506 = ~n386 & n2505;
  assign n2507 = ~n228 & n2506;
  assign n2508 = ~\V133(10)  & \V116(21) ;
  assign n2509 = ~n510 & n2508;
  assign n2510 = ~n507 & n2509;
  assign n2511 = ~n504 & n2510;
  assign n2512 = ~n386 & n2511;
  assign n2513 = n228 & n2512;
  assign n2514 = n419 & n578;
  assign n2515 = n406 & n2514;
  assign n2516 = ~n394 & n2515;
  assign n2517 = \V47(10)  & n422;
  assign n2518 = n419 & n2517;
  assign n2519 = ~n406 & n2518;
  assign n2520 = ~n419 & n778;
  assign n2521 = \V47(21)  & ~n422;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = ~n2519 & n2522;
  assign n2524 = ~n2516 & n2523;
  assign n2525 = ~n425 & n2524;
  assign n2526 = \V133(10)  & ~n2525;
  assign n2527 = ~n510 & n2526;
  assign n2528 = ~n507 & n2527;
  assign n2529 = ~n504 & n2528;
  assign n2530 = ~n386 & n2529;
  assign n2531 = ~n510 & ~n2525;
  assign n2532 = ~n507 & n2531;
  assign n2533 = ~n504 & n2532;
  assign n2534 = n386 & n2533;
  assign n2535 = n504 & n2532;
  assign n2536 = n507 & n2531;
  assign n2537 = n510 & ~n2525;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = ~n2535 & n2538;
  assign n2540 = ~n2534 & n2539;
  assign n2541 = ~n2530 & n2540;
  assign n2542 = ~n2513 & n2541;
  assign \V165(4)  = n2507 | ~n2542;
  assign n2544 = ~n227 & n2030;
  assign n2545 = ~n223 & n2544;
  assign n2546 = ~n221 & n2545;
  assign n2547 = \V84(29)  & \V133(10) ;
  assign n2548 = ~n227 & n2547;
  assign n2549 = ~n223 & n2548;
  assign n2550 = \V84(29)  & ~n227;
  assign n2551 = n223 & n2550;
  assign n2552 = \V84(29)  & n227;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~n2549 & n2553;
  assign n2555 = ~n235 & n2554;
  assign \V212(12)  = n2546 | ~n2555;
  assign n2557 = ~\V133(1)  & ~\V133(9) ;
  assign n2558 = ~\V133(4)  & n2557;
  assign n2559 = \V84(12)  & n511;
  assign n2560 = ~\V133(9)  & n2559;
  assign n2561 = ~\V133(4)  & n2560;
  assign n2562 = ~n2558 & n2561;
  assign n2563 = ~n507 & n2562;
  assign n2564 = ~n504 & n2563;
  assign n2565 = ~n386 & n2564;
  assign n2566 = ~n228 & n2565;
  assign n2567 = \V116(12)  & ~\V133(10) ;
  assign n2568 = ~n2558 & n2567;
  assign n2569 = ~n507 & n2568;
  assign n2570 = ~n504 & n2569;
  assign n2571 = ~n386 & n2570;
  assign n2572 = n228 & n2571;
  assign n2573 = \V15(11)  & n422;
  assign n2574 = n419 & n2573;
  assign n2575 = n406 & n2574;
  assign n2576 = ~n394 & n2575;
  assign n2577 = n419 & n433;
  assign n2578 = ~n406 & n2577;
  assign n2579 = ~n419 & n530;
  assign n2580 = \V47(12)  & ~n422;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2578 & n2581;
  assign n2583 = ~n2576 & n2582;
  assign n2584 = ~n425 & n2583;
  assign n2585 = \V133(10)  & ~n2584;
  assign n2586 = ~n2558 & n2585;
  assign n2587 = ~n507 & n2586;
  assign n2588 = ~n504 & n2587;
  assign n2589 = ~n386 & n2588;
  assign n2590 = ~n2558 & ~n2584;
  assign n2591 = ~n507 & n2590;
  assign n2592 = ~n504 & n2591;
  assign n2593 = n386 & n2592;
  assign n2594 = n504 & n2591;
  assign n2595 = n507 & n2590;
  assign n2596 = n2558 & ~n2584;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~n2594 & n2597;
  assign n2599 = ~n2593 & n2598;
  assign n2600 = ~n2589 & n2599;
  assign n2601 = ~n2572 & n2600;
  assign \V146(0)  = n2566 | ~n2601;
  assign n2603 = ~n227 & n2101;
  assign n2604 = ~n223 & n2603;
  assign n2605 = ~n221 & n2604;
  assign n2606 = \V84(31)  & \V133(10) ;
  assign n2607 = ~n227 & n2606;
  assign n2608 = ~n223 & n2607;
  assign n2609 = \V84(31)  & ~n227;
  assign n2610 = n223 & n2609;
  assign n2611 = \V84(31)  & n227;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2608 & n2612;
  assign n2614 = ~n235 & n2613;
  assign \V212(14)  = n2605 | ~n2614;
  assign n2616 = \V84(18)  & n511;
  assign n2617 = ~\V133(9)  & n2616;
  assign n2618 = ~\V133(4)  & n2617;
  assign n2619 = ~n510 & n2618;
  assign n2620 = ~n507 & n2619;
  assign n2621 = ~n504 & n2620;
  assign n2622 = ~n386 & n2621;
  assign n2623 = ~n228 & n2622;
  assign n2624 = ~\V133(10)  & \V116(18) ;
  assign n2625 = ~n510 & n2624;
  assign n2626 = ~n507 & n2625;
  assign n2627 = ~n504 & n2626;
  assign n2628 = ~n386 & n2627;
  assign n2629 = n228 & n2628;
  assign n2630 = n406 & n576;
  assign n2631 = ~n394 & n2630;
  assign n2632 = ~n406 & n2458;
  assign n2633 = ~n419 & n2517;
  assign n2634 = \V47(18)  & ~n422;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = ~n2632 & n2635;
  assign n2637 = ~n2631 & n2636;
  assign n2638 = ~n425 & n2637;
  assign n2639 = \V133(10)  & ~n2638;
  assign n2640 = ~n510 & n2639;
  assign n2641 = ~n507 & n2640;
  assign n2642 = ~n504 & n2641;
  assign n2643 = ~n386 & n2642;
  assign n2644 = ~n510 & ~n2638;
  assign n2645 = ~n507 & n2644;
  assign n2646 = ~n504 & n2645;
  assign n2647 = n386 & n2646;
  assign n2648 = n504 & n2645;
  assign n2649 = n507 & n2644;
  assign n2650 = n510 & ~n2638;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = ~n2648 & n2651;
  assign n2653 = ~n2647 & n2652;
  assign n2654 = ~n2643 & n2653;
  assign n2655 = ~n2629 & n2654;
  assign \V165(1)  = n2623 | ~n2655;
  assign n2657 = \V84(17)  & n511;
  assign n2658 = ~\V133(9)  & n2657;
  assign n2659 = ~\V133(4)  & n2658;
  assign n2660 = ~n510 & n2659;
  assign n2661 = ~n507 & n2660;
  assign n2662 = ~n504 & n2661;
  assign n2663 = ~n386 & n2662;
  assign n2664 = ~n228 & n2663;
  assign n2665 = ~\V133(10)  & \V116(17) ;
  assign n2666 = ~n510 & n2665;
  assign n2667 = ~n507 & n2666;
  assign n2668 = ~n504 & n2667;
  assign n2669 = ~n386 & n2668;
  assign n2670 = n228 & n2669;
  assign n2671 = n406 & n621;
  assign n2672 = ~n394 & n2671;
  assign n2673 = ~n406 & n2514;
  assign n2674 = ~n419 & n2347;
  assign n2675 = \V47(17)  & ~n422;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2673 & n2676;
  assign n2678 = ~n2672 & n2677;
  assign n2679 = ~n425 & n2678;
  assign n2680 = \V133(10)  & ~n2679;
  assign n2681 = ~n510 & n2680;
  assign n2682 = ~n507 & n2681;
  assign n2683 = ~n504 & n2682;
  assign n2684 = ~n386 & n2683;
  assign n2685 = ~n510 & ~n2679;
  assign n2686 = ~n507 & n2685;
  assign n2687 = ~n504 & n2686;
  assign n2688 = n386 & n2687;
  assign n2689 = n504 & n2686;
  assign n2690 = n507 & n2685;
  assign n2691 = n510 & ~n2679;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~n2689 & n2692;
  assign n2694 = ~n2688 & n2693;
  assign n2695 = ~n2684 & n2694;
  assign n2696 = ~n2670 & n2695;
  assign \V165(0)  = n2664 | ~n2696;
  assign n2698 = \V84(24)  & n511;
  assign n2699 = ~\V133(9)  & n2698;
  assign n2700 = ~\V133(4)  & n2699;
  assign n2701 = ~n510 & n2700;
  assign n2702 = ~n507 & n2701;
  assign n2703 = ~n504 & n2702;
  assign n2704 = ~n386 & n2703;
  assign n2705 = ~n228 & n2704;
  assign n2706 = ~\V133(10)  & \V116(24) ;
  assign n2707 = ~n510 & n2706;
  assign n2708 = ~n507 & n2707;
  assign n2709 = ~n504 & n2708;
  assign n2710 = ~n386 & n2709;
  assign n2711 = n228 & n2710;
  assign n2712 = n406 & n2348;
  assign n2713 = ~n394 & n2712;
  assign n2714 = ~n406 & n779;
  assign n2715 = ~n419 & n883;
  assign n2716 = \V47(24)  & ~n422;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = ~n2714 & n2717;
  assign n2719 = ~n2713 & n2718;
  assign n2720 = ~n425 & n2719;
  assign n2721 = \V133(10)  & ~n2720;
  assign n2722 = ~n510 & n2721;
  assign n2723 = ~n507 & n2722;
  assign n2724 = ~n504 & n2723;
  assign n2725 = ~n386 & n2724;
  assign n2726 = ~n510 & ~n2720;
  assign n2727 = ~n507 & n2726;
  assign n2728 = ~n504 & n2727;
  assign n2729 = n386 & n2728;
  assign n2730 = n504 & n2727;
  assign n2731 = n507 & n2726;
  assign n2732 = n510 & ~n2720;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = ~n2730 & n2733;
  assign n2735 = ~n2729 & n2734;
  assign n2736 = ~n2725 & n2735;
  assign n2737 = ~n2711 & n2736;
  assign \V165(7)  = n2705 | ~n2737;
  assign n2739 = \V84(23)  & n511;
  assign n2740 = ~\V133(9)  & n2739;
  assign n2741 = ~\V133(4)  & n2740;
  assign n2742 = ~n510 & n2741;
  assign n2743 = ~n507 & n2742;
  assign n2744 = ~n504 & n2743;
  assign n2745 = ~n386 & n2744;
  assign n2746 = ~n228 & n2745;
  assign n2747 = ~\V133(10)  & \V116(23) ;
  assign n2748 = ~n510 & n2747;
  assign n2749 = ~n507 & n2748;
  assign n2750 = ~n504 & n2749;
  assign n2751 = ~n386 & n2750;
  assign n2752 = n228 & n2751;
  assign n2753 = n406 & n2404;
  assign n2754 = ~n394 & n2753;
  assign n2755 = ~n406 & n880;
  assign n2756 = ~n419 & n964;
  assign n2757 = \V47(23)  & ~n422;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = ~n2755 & n2758;
  assign n2760 = ~n2754 & n2759;
  assign n2761 = ~n425 & n2760;
  assign n2762 = \V133(10)  & ~n2761;
  assign n2763 = ~n510 & n2762;
  assign n2764 = ~n507 & n2763;
  assign n2765 = ~n504 & n2764;
  assign n2766 = ~n386 & n2765;
  assign n2767 = ~n510 & ~n2761;
  assign n2768 = ~n507 & n2767;
  assign n2769 = ~n504 & n2768;
  assign n2770 = n386 & n2769;
  assign n2771 = n504 & n2768;
  assign n2772 = n507 & n2767;
  assign n2773 = n510 & ~n2761;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = ~n2771 & n2774;
  assign n2776 = ~n2770 & n2775;
  assign n2777 = ~n2766 & n2776;
  assign n2778 = ~n2752 & n2777;
  assign \V165(6)  = n2746 | ~n2778;
  assign n2780 = \V84(26)  & n511;
  assign n2781 = ~\V133(9)  & n2780;
  assign n2782 = ~\V133(4)  & n2781;
  assign n2783 = ~n510 & n2782;
  assign n2784 = ~n507 & n2783;
  assign n2785 = ~n504 & n2784;
  assign n2786 = ~n386 & n2785;
  assign n2787 = ~n228 & n2786;
  assign n2788 = ~\V133(10)  & \V116(26) ;
  assign n2789 = ~n510 & n2788;
  assign n2790 = ~n507 & n2789;
  assign n2791 = ~n504 & n2790;
  assign n2792 = ~n386 & n2791;
  assign n2793 = n228 & n2792;
  assign n2794 = n406 & n2461;
  assign n2795 = ~n394 & n2794;
  assign n2796 = ~n406 & n965;
  assign n2797 = ~n419 & n1050;
  assign n2798 = \V47(26)  & ~n422;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = ~n2796 & n2799;
  assign n2801 = ~n2795 & n2800;
  assign n2802 = ~n425 & n2801;
  assign n2803 = \V133(10)  & ~n2802;
  assign n2804 = ~n510 & n2803;
  assign n2805 = ~n507 & n2804;
  assign n2806 = ~n504 & n2805;
  assign n2807 = ~n386 & n2806;
  assign n2808 = ~n510 & ~n2802;
  assign n2809 = ~n507 & n2808;
  assign n2810 = ~n504 & n2809;
  assign n2811 = n386 & n2810;
  assign n2812 = n504 & n2809;
  assign n2813 = n507 & n2808;
  assign n2814 = n510 & ~n2802;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~n2812 & n2815;
  assign n2817 = ~n2811 & n2816;
  assign n2818 = ~n2807 & n2817;
  assign n2819 = ~n2793 & n2818;
  assign \V165(9)  = n2787 | ~n2819;
  assign n2821 = \V84(25)  & n511;
  assign n2822 = ~\V133(9)  & n2821;
  assign n2823 = ~\V133(4)  & n2822;
  assign n2824 = ~n510 & n2823;
  assign n2825 = ~n507 & n2824;
  assign n2826 = ~n504 & n2825;
  assign n2827 = ~n386 & n2826;
  assign n2828 = ~n228 & n2827;
  assign n2829 = ~\V133(10)  & \V116(25) ;
  assign n2830 = ~n510 & n2829;
  assign n2831 = ~n507 & n2830;
  assign n2832 = ~n504 & n2831;
  assign n2833 = ~n386 & n2832;
  assign n2834 = n228 & n2833;
  assign n2835 = n406 & n2518;
  assign n2836 = ~n394 & n2835;
  assign n2837 = ~n406 & n1047;
  assign n2838 = ~n419 & n782;
  assign n2839 = \V47(25)  & ~n422;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = ~n2837 & n2840;
  assign n2842 = ~n2836 & n2841;
  assign n2843 = ~n425 & n2842;
  assign n2844 = \V133(10)  & ~n2843;
  assign n2845 = ~n510 & n2844;
  assign n2846 = ~n507 & n2845;
  assign n2847 = ~n504 & n2846;
  assign n2848 = ~n386 & n2847;
  assign n2849 = ~n510 & ~n2843;
  assign n2850 = ~n507 & n2849;
  assign n2851 = ~n504 & n2850;
  assign n2852 = n386 & n2851;
  assign n2853 = n504 & n2850;
  assign n2854 = n507 & n2849;
  assign n2855 = n510 & ~n2843;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = ~n2853 & n2856;
  assign n2858 = ~n2852 & n2857;
  assign n2859 = ~n2848 & n2858;
  assign n2860 = ~n2834 & n2859;
  assign \V165(8)  = n2828 | ~n2860;
  assign n2862 = ~\V133(9)  & n215;
  assign n2863 = ~\V133(4)  & n2862;
  assign n2864 = \V84(16)  & n511;
  assign n2865 = ~\V133(9)  & n2864;
  assign n2866 = ~\V133(4)  & n2865;
  assign n2867 = ~n2863 & n2866;
  assign n2868 = ~n510 & n2867;
  assign n2869 = ~n507 & n2868;
  assign n2870 = ~n504 & n2869;
  assign n2871 = ~n386 & n2870;
  assign n2872 = ~n228 & n2871;
  assign n2873 = ~\V133(10)  & \V116(16) ;
  assign n2874 = ~n2863 & n2873;
  assign n2875 = ~n510 & n2874;
  assign n2876 = ~n507 & n2875;
  assign n2877 = ~n504 & n2876;
  assign n2878 = ~n386 & n2877;
  assign n2879 = n228 & n2878;
  assign n2880 = n406 & n2577;
  assign n2881 = ~n394 & n2880;
  assign n2882 = ~n406 & n2344;
  assign n2883 = ~n419 & n2403;
  assign n2884 = \V47(16)  & ~n422;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2882 & n2885;
  assign n2887 = ~n2881 & n2886;
  assign n2888 = ~n425 & n2887;
  assign n2889 = \V133(10)  & ~n2888;
  assign n2890 = ~n2863 & n2889;
  assign n2891 = ~n510 & n2890;
  assign n2892 = ~n507 & n2891;
  assign n2893 = ~n504 & n2892;
  assign n2894 = ~n386 & n2893;
  assign n2895 = ~n2863 & ~n2888;
  assign n2896 = ~n510 & n2895;
  assign n2897 = ~n507 & n2896;
  assign n2898 = ~n504 & n2897;
  assign n2899 = n386 & n2898;
  assign n2900 = n504 & n2897;
  assign n2901 = n507 & n2896;
  assign n2902 = n510 & n2895;
  assign n2903 = n2863 & ~n2888;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = ~n2901 & n2904;
  assign n2906 = ~n2900 & n2905;
  assign n2907 = ~n2899 & n2906;
  assign n2908 = ~n2894 & n2907;
  assign n2909 = ~n2879 & n2908;
  assign \V150(0)  = n2872 | ~n2909;
endmodule


