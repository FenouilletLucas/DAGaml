// Benchmark "TOP" written by ABC on Sun Apr 24 20:33:51 2016

module TOP ( clock, 
    Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227, Pg3226,
    Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218, Pg3217,
    Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249, Pg563,
    Pg51, PCLK,
    Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435, Pg25420,
    Pg24734, Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275, Pg8274,
    Pg8273, Pg8272, Pg8271, Pg8270, Pg8269, Pg8268, Pg8267, Pg8266, Pg8265,
    Pg8264, Pg8263, Pg8262, Pg8261, Pg8260, Pg8259, Pg8258, Pg8251, Pg8249,
    Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, Pg8082, Pg8030, Pg8023, Pg8021,
    Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, Pg7487, Pg7425, Pg7390,
    Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, Pg7084, Pg7052,
    Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750, Pg6712,
    Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368, Pg6313,
    Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657, Pg5648,
    Pg5637, Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472, Pg5437,
    Pg5388, Pg4590, Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088, Pg3993  );
  input  clock;
  input  Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227,
    Pg3226, Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218,
    Pg3217, Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249,
    Pg563, Pg51, PCLK;
  output Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435,
    Pg25420, Pg24734, Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275,
    Pg8274, Pg8273, Pg8272, Pg8271, Pg8270, Pg8269, Pg8268, Pg8267, Pg8266,
    Pg8265, Pg8264, Pg8263, Pg8262, Pg8261, Pg8260, Pg8259, Pg8258, Pg8251,
    Pg8249, Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, Pg8082, Pg8030, Pg8023,
    Pg8021, Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, Pg7487, Pg7425,
    Pg7390, Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, Pg7084,
    Pg7052, Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750,
    Pg6712, Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368,
    Pg6313, Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657,
    Pg5648, Pg5637, Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472,
    Pg5437, Pg5388, Pg4590, Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088,
    Pg3993;
  reg Pg8021, Ng2817, Ng2933, Ng13457, Ng2883, Ng2888, Ng2896, Ng2892,
    Ng2903, Ng2900, Ng2908, Ng2912, Ng2917, Ng2924, Ng2920, Ng2984, Ng2985,
    Ng2929, Ng2879, Ng2934, Ng2935, Ng2938, Ng2941, Ng2944, Ng2947, Ng2953,
    Ng2956, Ng2959, Ng2962, Ng2963, Ng2966, Ng2969, Ng2972, Ng2975, Ng2978,
    Ng2981, Ng2874, Ng1506, Ng1501, Ng1496, Ng1491, Ng1486, Ng1481, Ng1476,
    Ng1471, Ng13439, Pg8251, Ng813, Pg4090, Ng809, Pg4323, Ng805, Pg4590,
    Ng801, Pg6225, Ng797, Pg6442, Ng793, Pg6895, Ng789, Pg7334, Ng785,
    Pg7519, Ng13423, Pg8249, Ng125, Pg4088, Ng121, Pg4321, Ng117, Pg8023,
    Ng113, Pg8175, Ng109, Pg3993, Ng105, Pg4200, Ng101, Pg4450, Ng97,
    Pg8096, Ng13407, Ng2200, Ng2195, Ng2190, Ng2185, Ng2180, Ng2175,
    Ng2170, Ng2165, Ng13455, Ng3210, Ng3211, Ng3084, Ng3085, Ng3086,
    Ng3087, Ng3091, Ng3092, Ng3093, Ng3094, Ng3095, Ng3096, Ng3097, Ng3098,
    Ng3099, Ng3100, Ng3101, Ng3102, Ng3103, Ng3104, Ng3105, Ng3106, Ng3107,
    Ng3108, Ng3155, Ng3158, Ng3161, Ng3164, Ng3167, Ng3170, Ng3173, Ng3176,
    Ng3179, Ng3182, Ng3185, Ng3088, Ng3191, Ng3128, Ng3126, Ng3125, Ng3123,
    Ng3120, Ng3110, Ng3139, Ng3135, Ng3147, Ng185, Ng130, Ng131, Ng129,
    Ng133, Ng134, Ng132, Ng142, Ng143, Ng141, Ng145, Ng146, Ng144, Ng148,
    Ng149, Ng147, Ng151, Ng152, Ng150, Ng154, Ng155, Ng153, Ng157, Ng158,
    Ng156, Ng160, Ng161, Ng159, Ng163, Ng164, Ng162, Ng169, Ng170, Ng168,
    Ng172, Ng173, Ng171, Ng175, Ng176, Ng174, Ng178, Ng179, Ng177, Ng186,
    Ng189, Ng192, Ng231, Ng234, Ng237, Ng195, Ng198, Ng201, Ng240, Ng243,
    Ng246, Ng204, Ng207, Ng210, Ng249, Ng252, Ng255, Ng213, Ng216, Ng219,
    Ng258, Ng261, Ng264, Ng222, Ng225, Ng228, Ng267, Ng270, Ng273, Ng92,
    Ng88, Ng83, Ng79, Ng74, Ng70, Ng65, Ng61, Ng56, Ng52, Ng11497, Ng11498,
    Ng11499, Ng11500, Ng11501, Ng11502, Ng11503, Ng11504, Ng11505, Ng11506,
    Ng11507, Ng11508, Ng408, Ng411, Ng414, Ng417, Ng420, Ng423, Ng427,
    Ng428, Ng426, Ng429, Ng432, Ng435, Ng438, Ng441, Ng444, Ng448, Ng449,
    Ng447, Ng312, Ng313, Ng314, Ng315, Ng316, Ng317, Ng318, Ng319, Ng320,
    Ng322, Ng323, Ng321, Ng403, Ng404, Ng402, Ng450, Ng451, Ng452, Ng453,
    Ng454, Ng279, Ng280, Ng281, Ng282, Ng283, Ng284, Ng285, Ng286, Ng287,
    Ng288, Ng289, Ng290, Ng291, Ng299, Ng305, Ng298, Ng342, Ng349, Ng350,
    Ng351, Ng352, Ng353, Ng357, Ng364, Ng365, Ng366, Ng367, Ng368, Ng372,
    Ng379, Ng380, Ng381, Ng382, Ng383, Ng387, Ng394, Ng395, Ng396, Ng397,
    Ng324, Ng554, Ng557, Ng510, Ng513, Ng523, Ng524, Ng564, Ng569, Ng570,
    Ng571, Ng572, Ng573, Ng574, Ng565, Ng566, Ng567, Ng568, Ng489, Ng486,
    Ng487, Ng488, Ng11512, Ng11515, Ng11516, Ng477, Ng478, Ng479, Ng480,
    Ng484, Ng464, Ng11517, Ng11513, Ng11514, Ng528, Ng535, Ng542, Ng543,
    Ng544, Ng548, Ng549, Ng8284, Ng558, Ng559, Ng576, Ng577, Ng575, Ng579,
    Ng580, Ng578, Ng582, Ng583, Ng581, Ng585, Ng586, Ng584, Ng587, Ng590,
    Ng593, Ng596, Ng599, Ng602, Ng614, Ng617, Ng620, Ng605, Ng608, Ng611,
    Ng490, Ng493, Ng496, Ng506, Ng507, Pg16297, Ng525, Ng529, Ng530, Ng531,
    Ng532, Ng533, Ng534, Ng536, Ng537, Ng538, Ng541, Ng630, Ng659, Ng640,
    Ng633, Ng653, Ng646, Ng660, Ng672, Ng666, Ng679, Ng686, Ng692, Ng699,
    Ng700, Ng698, Ng702, Ng703, Ng701, Ng705, Ng706, Ng704, Ng708, Ng709,
    Ng707, Ng711, Ng712, Ng710, Ng714, Ng715, Ng713, Ng717, Ng718, Ng716,
    Ng720, Ng721, Ng719, Ng723, Ng724, Ng722, Ng726, Ng727, Ng725, Ng729,
    Ng730, Ng728, Ng732, Ng733, Ng731, Ng735, Ng736, Ng734, Ng738, Ng739,
    Ng737, \[1612] , \[1594] , Ng853, Ng818, Ng819, Ng817, Ng821, Ng822,
    Ng820, Ng830, Ng831, Ng829, Ng833, Ng834, Ng832, Ng836, Ng837, Ng835,
    Ng839, Ng840, Ng838, Ng842, Ng843, Ng841, Ng845, Ng846, Ng844, Ng848,
    Ng849, Ng847, Ng851, Ng852, Ng850, Ng857, Ng858, Ng856, Ng860, Ng861,
    Ng859, Ng863, Ng864, Ng862, Ng866, Ng867, Ng865, Ng873, Ng876, Ng879,
    Ng918, Ng921, Ng924, Ng882, Ng885, Ng888, Ng927, Ng930, Ng933, Ng891,
    Ng894, Ng897, Ng936, Ng939, Ng942, Ng900, Ng903, Ng906, Ng945, Ng948,
    Ng951, Ng909, Ng912, Ng915, Ng954, Ng957, Ng960, Ng780, Ng776, Ng771,
    Ng767, Ng762, Ng758, Ng753, Ng749, Ng744, Ng740, Ng11524, Ng11525,
    Ng11526, Ng11527, Ng11528, Ng11529, Ng11530, Ng11531, Ng11532, Ng11533,
    Ng11534, Ng11535, Ng1095, Ng1098, Ng1101, Ng1104, Ng1107, Ng1110,
    Ng1114, Ng1115, Ng1113, Ng1116, Ng1119, Ng1122, Ng1125, Ng1128, Ng1131,
    Ng1135, Ng1136, Ng1134, Ng999, Ng1000, Ng1001, Ng1002, Ng1003, Ng1004,
    Ng1005, Ng1006, Ng1007, Ng1009, Ng1010, Ng1008, Ng1090, Ng1091, Ng1089,
    Ng1137, Ng1138, Ng1139, Ng1140, Ng1141, Ng966, Ng967, Ng968, Ng969,
    Ng970, Ng971, Ng972, Ng973, Ng974, Ng975, Ng976, Ng977, Ng978, Ng986,
    Ng992, Ng985, Ng1029, Ng1036, Ng1037, Ng1038, Ng1039, Ng1040, Ng1044,
    Ng1051, Ng1052, Ng1053, Ng1054, Ng1055, Ng1059, Ng1066, Ng1067, Ng1068,
    Ng1069, Ng1070, Ng1074, Ng1081, Ng1082, Ng1083, Ng1084, Ng1011, Ng1240,
    Ng1243, Ng1196, Ng1199, Ng1209, Ng1210, Ng1250, Ng1255, Ng1256, Ng1257,
    Ng1258, Ng1259, Ng1260, Ng1251, Ng1252, Ng1253, Ng1254, Ng1176, Ng1173,
    Ng1174, Ng1175, Ng11539, Ng11542, Ng11543, Ng1164, Ng1165, Ng1166,
    Ng1167, Ng1171, Ng1151, Ng11544, Ng11540, Ng11541, Ng1214, Ng1221,
    Ng1228, Ng1229, Ng1230, Ng1234, Ng1235, Ng8293, Ng1244, Ng1245, Ng1262,
    Ng1263, Ng1261, Ng1265, Ng1266, Ng1264, Ng1268, Ng1269, Ng1267, Ng1271,
    Ng1272, Ng1270, Ng1273, Ng1276, Ng1279, Ng1282, Ng1285, Ng1288, Ng1300,
    Ng1303, Ng1306, Ng1291, Ng1294, Ng1297, Ng1177, Ng1180, Ng1183, Ng1192,
    Ng1193, Pg16355, Ng1211, Ng1215, Ng1216, Ng1217, Ng1218, Ng1219,
    Ng1220, Ng1222, Ng1223, Ng1224, Ng1227, \[1605] , \[1603] , Ng1315,
    Ng1316, Ng1345, Ng1326, Ng1319, Ng1339, Ng1332, Ng1346, Ng1358, Ng1352,
    Ng1365, Ng1372, Ng1378, Ng1385, Ng1386, Ng1384, Ng1388, Ng1389, Ng1387,
    Ng1391, Ng1392, Ng1390, Ng1394, Ng1395, Ng1393, Ng1397, Ng1398, Ng1396,
    Ng1400, Ng1401, Ng1399, Ng1403, Ng1404, Ng1402, Ng1406, Ng1407, Ng1405,
    Ng1409, Ng1410, Ng1408, Ng1412, Ng1413, Ng1411, Ng1415, Ng1416, Ng1414,
    Ng1418, Ng1419, Ng1417, Ng1421, Ng1422, Ng1420, Ng1424, Ng1425, Ng1423,
    Ng1512, Ng1513, Ng1511, Ng1515, Ng1516, Ng1514, Ng1524, Ng1525, Ng1523,
    Ng1527, Ng1528, Ng1526, Ng1530, Ng1531, Ng1529, Ng1533, Ng1534, Ng1532,
    Ng1536, Ng1537, Ng1535, Ng1539, Ng1540, Ng1538, Ng1542, Ng1543, Ng1541,
    Ng1545, Ng1546, Ng1544, Ng1551, Ng1552, Ng1550, Ng1554, Ng1555, Ng1553,
    Ng1557, Ng1558, Ng1556, Ng1560, Ng1561, Ng1559, Ng1567, Ng1570, Ng1573,
    Ng1612, Ng1615, Ng1618, Ng1576, Ng1579, Ng1582, Ng1621, Ng1624, Ng1627,
    Ng1585, Ng1588, Ng1591, Ng1630, Ng1633, Ng1636, Ng1594, Ng1597, Ng1600,
    Ng1639, Ng1642, Ng1645, Ng1603, Ng1606, Ng1609, Ng1648, Ng1651, Ng1654,
    Ng1466, Ng1462, Ng1457, Ng1453, Ng1448, Ng1444, Ng1439, Ng1435, Ng1430,
    Ng1426, Ng11551, Ng11552, Ng11553, Ng11554, Ng11555, Ng11556, Ng11557,
    Ng11558, Ng11559, Ng11560, Ng11561, Ng11562, Ng1789, Ng1792, Ng1795,
    Ng1798, Ng1801, Ng1804, Ng1808, Ng1809, Ng1807, Ng1810, Ng1813, Ng1816,
    Ng1819, Ng1822, Ng1825, Ng1829, Ng1830, Ng1828, Ng1693, Ng1694, Ng1695,
    Ng1696, Ng1697, Ng1698, Ng1699, Ng1700, Ng1701, Ng1703, Ng1704, Ng1702,
    Ng1784, Ng1785, Ng1783, Ng1831, Ng1832, Ng1833, Ng1834, Ng1835, Ng1660,
    Ng1661, Ng1662, Ng1663, Ng1664, Ng1665, Ng1666, Ng1667, Ng1668, Ng1669,
    Ng1670, Ng1671, Ng1672, Ng1680, Ng1686, Ng1679, Ng1723, Ng1730, Ng1731,
    Ng1732, Ng1733, Ng1734, Ng1738, Ng1745, Ng1746, Ng1747, Ng1748, Ng1749,
    Ng1753, Ng1760, Ng1761, Ng1762, Ng1763, Ng1764, Ng1768, Ng1775, Ng1776,
    Ng1777, Ng1778, Ng1705, Ng1934, Ng1937, Ng1890, Ng1893, Ng1903, Ng1904,
    Ng1944, Ng1949, Ng1950, Ng1951, Ng1952, Ng1953, Ng1954, Ng1945, Ng1946,
    Ng1947, Ng1948, Ng1870, Ng1867, Ng1868, Ng1869, Ng11566, Ng11569,
    Ng11570, Ng1858, Ng1859, Ng1860, Ng1861, Ng1865, Ng1845, Ng11571,
    Ng11567, Ng11568, Ng1908, Ng1915, Ng1922, Ng1923, Ng1924, Ng1928,
    Ng1929, Ng8302, Ng1938, Ng1939, Ng1956, Ng1957, Ng1955, Ng1959, Ng1960,
    Ng1958, Ng1962, Ng1963, Ng1961, Ng1965, Ng1966, Ng1964, Ng1967, Ng1970,
    Ng1973, Ng1976, Ng1979, Ng1982, Ng1994, Ng1997, Ng2000, Ng1985, Ng1988,
    Ng1991, Ng1871, Ng1874, Ng1877, Ng1886, Ng1887, Pg16399, Ng1905,
    Ng1909, Ng1910, Ng1911, Ng1912, Ng1913, Ng1914, Ng1916, Ng1917, Ng1918,
    Ng1921, Ng2010, Ng2039, Ng2020, Ng2013, Ng2033, Ng2026, Ng2040, Ng2052,
    Ng2046, Ng2059, Ng2066, Ng2072, Ng2079, Ng2080, Ng2078, Ng2082, Ng2083,
    Ng2081, Ng2085, Ng2086, Ng2084, Ng2088, Ng2089, Ng2087, Ng2091, Ng2092,
    Ng2090, Ng2094, Ng2095, Ng2093, Ng2097, Ng2098, Ng2096, Ng2100, Ng2101,
    Ng2099, Ng2103, Ng2104, Ng2102, Ng2106, Ng2107, Ng2105, Ng2109, Ng2110,
    Ng2108, Ng2112, Ng2113, Ng2111, Ng2115, Ng2116, Ng2114, Ng2118, Ng2119,
    Ng2117, Ng2206, Ng2207, Ng2205, Ng2209, Ng2210, Ng2208, Ng2218, Ng2219,
    Ng2217, Ng2221, Ng2222, Ng2220, Ng2224, Ng2225, Ng2223, Ng2227, Ng2228,
    Ng2226, Ng2230, Ng2231, Ng2229, Ng2233, Ng2234, Ng2232, Ng2236, Ng2237,
    Ng2235, Ng2239, Ng2240, Ng2238, Ng2245, Ng2246, Ng2244, Ng2248, Ng2249,
    Ng2247, Ng2251, Ng2252, Ng2250, Ng2254, Ng2255, Ng2253, Ng2261, Ng2264,
    Ng2267, Ng2306, Ng2309, Ng2312, Ng2270, Ng2273, Ng2276, Ng2315, Ng2318,
    Ng2321, Ng2279, Ng2282, Ng2285, Ng2324, Ng2327, Ng2330, Ng2288, Ng2291,
    Ng2294, Ng2333, Ng2336, Ng2339, Ng2297, Ng2300, Ng2303, Ng2342, Ng2345,
    Ng2348, Ng2160, Ng2156, Ng2151, Ng2147, Ng2142, Ng2138, Ng2133, Ng2129,
    Ng2124, Ng2120, Ng2256, \[1609] , Ng2257, Ng11578, Ng11579, Ng11580,
    Ng11581, Ng11582, Ng11583, Ng11584, Ng11585, Ng11586, Ng11587, Ng11588,
    Ng11589, Ng2483, Ng2486, Ng2489, Ng2492, Ng2495, Ng2498, Ng2502,
    Ng2503, Ng2501, Ng2504, Ng2507, Ng2510, Ng2513, Ng2516, Ng2519, Ng2523,
    Ng2524, Ng2522, Ng2387, Ng2388, Ng2389, Ng2390, Ng2391, Ng2392, Ng2393,
    Ng2394, Ng2395, Ng2397, Ng2398, Ng2396, Ng2478, Ng2479, Ng2477, Ng2525,
    Ng2526, Ng2527, Ng2528, Ng2529, Ng2354, Ng2355, Ng2356, Ng2357, Ng2358,
    Ng2359, Ng2360, Ng2361, Ng2362, Ng2363, Ng2364, Ng2365, Ng2366, Ng2374,
    Ng2380, Ng2373, Ng2417, Ng2424, Ng2425, Ng2426, Ng2427, Ng2428, Ng2432,
    Ng2439, Ng2440, Ng2441, Ng2442, Ng2443, Ng2447, Ng2454, Ng2455, Ng2456,
    Ng2457, Ng2458, Ng2462, Ng2469, Ng2470, Ng2471, Ng2472, Ng2399, Ng2628,
    Ng2631, Ng2584, Ng2587, Ng2597, Ng2598, Ng2638, Ng2643, Ng2644, Ng2645,
    Ng2646, Ng2647, Ng2648, Ng2639, Ng2640, Ng2641, Ng2642, Ng2564, Ng2561,
    Ng2562, Ng2563, Ng11593, Ng11596, Ng11597, Ng2552, Ng2553, Ng2554,
    Ng2555, Ng2559, Ng2539, Ng11598, Ng11594, Ng11595, Ng2602, Ng2609,
    Ng2616, Ng2617, Ng2618, Ng2622, Ng2623, Ng8311, Ng2632, Ng2633, Ng2650,
    Ng2651, Ng2649, Ng2653, Ng2654, Ng2652, Ng2656, Ng2657, Ng2655, Ng2659,
    Ng2660, Ng2658, Ng2661, Ng2664, Ng2667, Ng2670, Ng2673, Ng2676, Ng2688,
    Ng2691, Ng2694, Ng2679, Ng2682, Ng2685, Ng2565, Ng2568, Ng2571, Ng2580,
    Ng2581, Pg16437, Ng2599, Ng2603, Ng2604, Ng2605, Ng2606, Ng2607,
    Ng2608, Ng2610, Ng2611, Ng2612, Ng2615, Ng2704, Ng2733, Ng2714, Ng2707,
    Ng2727, Ng2720, Ng2734, Ng2746, Ng2740, Ng2753, Ng2760, Ng2766, Ng2773,
    Ng2774, Ng2772, Ng2776, Ng2777, Ng2775, Ng2779, Ng2780, Ng2778, Ng2782,
    Ng2783, Ng2781, Ng2785, Ng2786, Ng2784, Ng2788, Ng2789, Ng2787, Ng2791,
    Ng2792, Ng2790, Ng2794, Ng2795, Ng2793, Ng2797, Ng2798, Ng2796, Ng2800,
    Ng2801, Ng2799, Ng2803, Ng2804, Ng2802, Ng2806, Ng2807, Ng2805, Ng2809,
    Ng2810, Ng2808, Ng2812, Ng2813, Ng2811, Ng3054, Ng3079, Ng13475,
    Ng3043, Ng3044, Ng3045, Ng3046, Ng3047, Ng3048, Ng3049, Ng3050, Ng3051,
    Ng3052, Ng3053, Ng3055, Ng3056, Ng3057, Ng3058, Ng3059, Ng3060, Ng3061,
    Ng3062, Ng3063, Ng3064, Ng3065, Ng3066, Ng3067, Ng3068, Ng3069, Ng3070,
    Ng3071, Ng3072, Ng3073, Ng3074, Ng3075, Ng3076, Ng3077, Ng3078, Ng2997,
    Ng2993, Ng2998, Ng3006, Ng3002, Ng3013, Ng3010, Ng3024, Ng3018, Ng3028,
    Ng3036, Ng3032, Pg5388, Ng2986, Ng2987, Pg8275, Pg8274, Pg8273, Pg8272,
    Pg8268, Pg8269, Pg8270, Pg8271, Ng3083, Pg8267, Ng2992, Pg8266, Pg8265,
    Pg8264, Pg8262, Pg8263, Pg8260, Pg8261, Pg8259, Ng2990, Ng2991, Pg8258;
  wire n4522_1, n4523, n4524, n4525, n4526, n4527_1, n4528, n4529, n4530,
    n4531, n4532_1, n4533, n4534, n4535, n4536, n4537_1, n4538, n4539,
    n4540, n4541, n4542_1, n4543, n4545, n4547_1, n4548, n4549, n4550,
    n4551_1, n4552, n4553, n4554, n4555, n4556_1, n4557, n4558, n4559,
    n4560_1, n4561, n4562, n4563, n4564, n4565_1, n4566, n4567, n4568,
    n4569_1, n4570, n4571, n4572, n4573, n4574_1, n4575, n4576, n4577,
    n4578_1, n4579, n4580, n4581, n4582, n4583_1, n4584, n4585, n4586,
    n4587_1, n4588, n4589, n4590, n4591, n4592_1, n4594, n4595, n4596_1,
    n4597, n4598, n4599, n4600, n4601_1, n4602, n4603, n4604, n4605_1,
    n4606, n4607, n4608, n4609, n4610_1, n4611, n4612, n4613, n4614_1,
    n4615, n4616, n4617, n4618_1, n4619, n4620, n4621, n4622_1, n4623,
    n4625, n4626, n4627_1, n4628, n4629, n4630, n4631, n4632_1, n4633,
    n4634, n4635, n4636, n4637_1, n4638, n4639, n4640, n4641_1, n4642,
    n4643, n4644, n4645_1, n4646, n4647, n4648, n4649_1, n4650, n4651,
    n4652, n4653_1, n4655, n4656, n4657_1, n4658, n4659, n4660, n4662,
    n4664, n4666, n4671, n4672, n4673_1, n4675, n4676, n4677_1, n4678,
    n4679, n4680, n4681_1, n4682, n4683, n4684, n4685_1, n4687, n4688,
    n4689_1, n4691, n4692, n4693_1, n4695, n4696, n4697_1, n4699, n4700,
    n4701_1, n4703, n4704, n4705_1, n4707, n4708, n4709_1, n4710, n4711,
    n4712, n4713_1, n4715, n4716, n4717_1, n4719, n4720, n4721_1, n4723,
    n4724, n4725_1, n4727, n4728, n4729_1, n4730, n4731, n4732, n4733_1,
    n4734, n4735, n4736, n4737, n4738_1, n4739, n4740, n4741, n4742,
    n4743_1, n4744, n4745, n4746, n4747, n4748_1, n4749, n4751, n4752,
    n4753_1, n4754, n4755, n4756, n4757_1, n4758, n4759, n4760, n4761_1,
    n4762, n4763, n4764, n4765, n4766_1, n4767, n4768, n4769, n4770_1,
    n4771, n4772, n4773, n4775_1, n4777, n4778, n4780, n4781, n4783,
    n4784_1, n4786, n4787, n4789, n4790, n4792, n4793_1, n4795, n4796,
    n4798, n4799, n4801, n4802_1, n4803, n4804, n4805, n4806_1, n4808,
    n4809, n4811_1, n4812, n4814, n4815_1, n4817, n4818, n4820_1, n4821,
    n4823, n4824, n4826, n4827, n4829, n4830_1, n4832, n4833, n4834,
    n4835_1, n4836, n4838, n4839_1, n4841, n4842, n4844, n4845, n4847_1,
    n4848, n4850, n4851, n4853, n4854, n4856, n4857_1, n4859, n4860,
    n4862_1, n4863, n4865, n4866, n4868, n4869, n4871, n4872, n4874, n4875,
    n4877_1, n4878, n4880, n4881_1, n4883, n4884, n4886, n4887, n4889_1,
    n4890, n4892, n4893, n4895, n4896, n4898, n4899, n4901, n4902_1, n4904,
    n4905, n4907, n4908, n4910, n4911_1, n4913, n4914, n4916_1, n4917,
    n4919, n4920_1, n4922, n4923, n4925_1, n4926, n4928, n4929_1, n4930,
    n4932, n4933, n4934_1, n4936, n4938, n4939_1, n4941, n4942, n4943,
    n4944_1, n4946, n4947, n4949_1, n4950, n4952, n4953, n4955, n4956,
    n4957, n4958, n4960, n4961, n4963, n4964_1, n4966, n4967, n4969_1,
    n4970, n4971, n4972, n4973, n4975, n4977, n4978, n4980, n4981, n4983,
    n4984_1, n4986, n4987, n4989_1, n4990, n4992, n4993, n4995, n4996,
    n4998, n4999_1, n5001, n5002, n5004_1, n5005, n5007, n5008, n5010,
    n5011, n5013, n5014_1, n5016, n5017, n5019_1, n5020, n5021, n5023,
    n5024_1, n5025, n5027, n5028, n5029_1, n5031, n5032, n5034_1, n5035,
    n5037, n5038, n5040, n5041, n5043, n5044_1, n5046, n5047, n5049_1,
    n5050, n5052, n5053, n5055, n5056, n5058, n5059_1, n5061, n5062,
    n5064_1, n5065, n5067, n5068_1, n5070, n5071, n5073_1, n5074, n5076,
    n5077, n5079, n5080, n5082, n5083, n5085, n5086_1, n5088, n5089,
    n5091_1, n5092, n5094, n5095, n5096_1, n5097, n5098, n5099, n5100,
    n5102, n5103, n5105, n5106_1, n5108, n5109, n5110, n5111_1, n5112,
    n5113, n5114, n5116_1, n5117, n5119, n5120, n5122, n5123, n5124, n5125,
    n5126_1, n5127, n5128, n5129, n5131_1, n5132, n5133, n5134, n5135,
    n5136_1, n5138, n5139, n5140, n5142, n5143, n5144, n5146_1, n5147,
    n5149, n5150, n5152, n5153, n5155, n5156_1, n5158, n5159, n5161_1,
    n5162, n5164, n5165, n5166_1, n5167, n5168, n5169, n5170, n5171_1,
    n5173, n5174, n5176_1, n5177, n5179, n5180, n5181_1, n5182, n5183,
    n5184, n5185, n5186_1, n5187, n5188, n5189, n5190, n5191_1, n5192,
    n5193, n5194, n5195, n5196_1, n5197, n5198, n5199, n5200, n5201_1,
    n5202, n5203, n5204, n5205, n5206_1, n5207, n5208, n5209, n5210,
    n5211_1, n5212, n5213, n5214, n5215, n5216_1, n5217, n5218, n5219,
    n5220, n5221_1, n5222, n5223, n5224, n5225, n5226_1, n5227, n5228,
    n5229, n5230, n5231_1, n5232, n5233, n5234, n5235, n5236_1, n5237,
    n5238, n5239, n5240, n5241_1, n5242, n5243, n5244, n5245, n5246_1,
    n5247, n5248, n5249, n5250, n5251_1, n5252, n5253, n5254, n5255,
    n5256_1, n5257, n5258, n5259, n5260, n5261_1, n5262, n5263, n5264,
    n5265, n5266_1, n5267, n5268, n5269, n5270, n5271_1, n5272, n5273,
    n5274, n5275, n5276_1, n5277, n5278, n5279, n5280, n5281_1, n5282,
    n5283, n5284, n5285, n5286_1, n5287, n5288, n5289, n5290, n5291_1,
    n5292, n5293, n5294, n5295, n5296_1, n5297, n5298, n5299, n5300,
    n5301_1, n5302, n5303, n5304, n5305, n5306_1, n5307, n5308, n5309,
    n5310, n5311_1, n5312, n5313, n5314, n5315, n5316_1, n5317, n5318,
    n5319, n5320, n5321_1, n5322, n5323, n5324, n5325, n5326_1, n5327,
    n5328, n5329, n5330, n5331_1, n5332, n5333, n5334, n5335, n5336_1,
    n5337, n5338, n5339, n5340, n5341_1, n5342, n5343, n5344, n5345,
    n5346_1, n5347, n5348, n5349, n5350, n5351_1, n5352, n5353, n5354,
    n5355, n5356_1, n5357, n5358, n5359, n5360, n5361_1, n5362, n5363,
    n5364, n5365, n5366_1, n5367, n5368, n5369, n5370, n5371_1, n5372,
    n5373, n5374, n5375, n5376_1, n5377, n5378, n5379, n5380, n5381_1,
    n5382, n5383, n5384, n5385, n5386_1, n5387, n5388, n5389, n5390,
    n5391_1, n5392, n5393, n5394, n5395, n5396_1, n5397, n5398, n5399,
    n5400, n5401_1, n5402, n5403, n5404, n5405, n5406_1, n5407, n5408,
    n5409, n5410, n5411_1, n5412, n5413, n5414, n5415, n5416_1, n5417,
    n5418, n5419, n5420, n5421_1, n5422, n5423, n5424, n5425, n5426_1,
    n5427, n5428, n5429, n5430, n5431_1, n5432, n5433, n5434, n5435,
    n5436_1, n5437, n5438, n5439, n5440, n5441_1, n5442, n5443, n5444,
    n5445, n5446_1, n5447, n5448, n5449, n5450, n5451_1, n5452, n5453,
    n5455, n5456_1, n5458, n5459, n5461_1, n5462, n5463, n5464, n5465,
    n5466_1, n5467, n5468, n5469, n5470, n5471_1, n5472, n5473, n5475,
    n5476_1, n5478, n5479, n5481_1, n5482, n5483, n5484, n5485, n5486_1,
    n5487, n5488, n5489, n5490, n5491_1, n5492, n5493, n5495, n5496_1,
    n5498, n5499, n5501_1, n5502, n5503, n5504, n5505, n5506_1, n5507,
    n5508, n5509, n5510, n5511_1, n5512, n5514, n5515, n5517, n5518, n5520,
    n5521_1, n5522, n5523, n5524, n5525, n5526_1, n5527, n5528, n5529,
    n5530, n5531_1, n5533, n5534, n5536_1, n5537, n5539, n5540, n5541_1,
    n5542, n5543, n5544, n5545, n5546_1, n5547, n5548, n5549, n5550, n5552,
    n5553, n5555, n5556_1, n5558, n5559, n5560, n5561_1, n5562, n5563,
    n5564, n5565, n5566_1, n5567, n5568, n5569, n5571_1, n5572, n5574,
    n5575, n5577, n5578, n5579, n5580, n5581_1, n5582, n5583, n5584, n5585,
    n5586_1, n5587, n5588, n5590, n5591_1, n5593, n5594, n5596_1, n5597,
    n5598, n5599, n5600, n5601_1, n5602, n5603, n5604, n5605, n5606_1,
    n5607, n5608, n5610, n5611_1, n5613, n5614, n5616_1, n5617, n5618,
    n5619, n5620, n5621_1, n5622, n5623, n5624, n5625, n5626_1, n5627,
    n5629, n5630, n5632, n5633, n5635, n5636_1, n5637, n5638, n5640,
    n5641_1, n5642, n5643, n5645, n5646_1, n5647, n5649, n5650, n5651_1,
    n5653, n5654, n5655, n5657, n5658, n5659, n5661_1, n5662, n5663, n5665,
    n5666_1, n5667, n5669, n5670, n5671_1, n5673, n5674, n5675, n5677,
    n5678, n5679, n5680, n5681_1, n5682, n5683, n5684, n5685, n5686_1,
    n5687, n5688, n5689, n5690, n5691_1, n5692, n5693, n5694, n5695,
    n5696_1, n5697, n5698, n5699, n5700, n5701_1, n5702, n5703, n5704,
    n5705, n5706_1, n5707, n5708, n5709, n5710, n5711_1, n5713, n5714,
    n5715, n5717, n5718, n5719, n5721_1, n5722, n5723, n5724, n5725,
    n5726_1, n5727, n5729, n5730, n5732, n5733, n5735, n5736_1, n5737,
    n5738, n5739, n5740, n5742, n5743, n5745, n5746_1, n5748, n5749, n5750,
    n5752, n5753, n5755, n5756_1, n5758, n5759, n5760, n5761_1, n5762,
    n5763, n5765, n5766_1, n5767, n5768, n5769, n5770, n5771_1, n5772,
    n5773, n5774, n5775, n5776_1, n5777, n5778, n5779, n5780, n5781_1,
    n5782, n5783, n5784, n5785, n5786_1, n5788, n5789, n5791_1, n5792,
    n5794, n5795, n5796_1, n5797, n5798, n5799, n5800, n5801_1, n5803,
    n5804, n5806_1, n5807, n5809, n5810, n5811_1, n5812, n5814, n5815,
    n5816_1, n5818, n5819, n5820_1, n5822, n5823, n5824_1, n5825, n5826,
    n5827, n5828, n5829_1, n5830, n5831, n5832, n5833, n5834_1, n5835,
    n5836, n5837, n5839_1, n5840, n5842, n5843, n5845, n5846, n5847, n5848,
    n5849_1, n5850, n5851, n5852, n5853, n5854_1, n5855, n5856, n5857,
    n5858, n5859_1, n5860, n5861, n5862, n5863, n5864_1, n5865, n5866,
    n5868, n5869_1, n5871, n5872, n5874_1, n5875, n5876, n5877, n5878,
    n5879_1, n5880, n5881, n5883, n5884_1, n5885, n5887, n5888, n5889_1,
    n5891, n5892, n5893, n5894_1, n5895, n5896, n5897, n5899_1, n5900,
    n5902, n5903, n5905, n5906, n5907, n5908, n5909_1, n5910, n5911, n5912,
    n5913, n5914_1, n5915, n5916, n5917, n5918, n5919_1, n5920, n5921,
    n5922, n5923, n5924_1, n5925, n5926, n5927, n5928, n5930, n5931, n5933,
    n5934_1, n5936, n5937, n5938, n5939_1, n5940, n5941, n5942, n5943,
    n5944_1, n5945, n5946, n5948, n5949_1, n5951, n5952, n5954_1, n5955,
    n5956, n5957, n5958, n5960, n5961, n5962, n5964_1, n5965, n5966, n5968,
    n5969_1, n5970, n5972, n5973, n5975, n5976, n5978, n5979_1, n5980,
    n5982, n5983, n5984_1, n5985, n5986, n5987, n5988, n5989_1, n5990,
    n5991, n5992, n5993, n5994_1, n5995, n5996, n5997, n5998, n5999_1,
    n6000, n6001, n6002, n6003, n6004_1, n6005, n6006, n6007, n6008,
    n6009_1, n6010, n6011, n6012, n6013, n6014_1, n6015, n6016, n6017,
    n6018, n6019_1, n6020, n6021, n6023, n6024_1, n6025, n6026, n6027,
    n6028, n6029_1, n6030, n6031, n6032, n6033, n6034_1, n6036, n6037,
    n6039_1, n6040, n6042, n6043, n6044_1, n6045, n6047, n6048, n6050,
    n6051, n6053, n6054_1, n6056, n6057, n6059, n6060, n6062, n6063_1,
    n6065, n6066, n6068, n6069, n6071, n6072_1, n6074, n6075, n6077, n6078,
    n6080, n6081_1, n6083, n6084, n6086, n6087, n6089, n6090_1, n6092,
    n6093, n6094_1, n6095, n6097, n6098, n6099_1, n6100, n6102, n6103_1,
    n6104, n6105, n6107, n6108_1, n6109, n6110, n6112_1, n6113, n6114,
    n6115, n6116, n6117_1, n6118, n6119, n6120, n6121_1, n6122, n6123,
    n6124, n6125_1, n6126, n6127, n6128, n6129_1, n6130, n6131, n6132,
    n6133, n6135, n6136, n6137, n6138, n6139_1, n6140, n6141, n6142, n6143,
    n6144_1, n6145, n6146, n6147, n6148_1, n6149, n6150, n6151, n6152_1,
    n6153, n6154, n6155, n6156_1, n6157, n6158, n6159, n6160_1, n6161,
    n6162, n6163, n6164_1, n6166, n6167, n6168_1, n6170, n6171, n6172_1,
    n6174, n6175, n6176_1, n6177, n6178, n6179, n6180_1, n6182, n6183,
    n6185, n6186, n6188_1, n6189, n6190, n6191, n6192_1, n6193, n6195,
    n6196_1, n6198, n6199, n6201, n6202, n6203, n6204_1, n6206, n6207,
    n6209, n6210, n6212_1, n6213, n6214, n6215, n6216_1, n6217, n6218,
    n6219, n6220_1, n6221, n6222, n6224_1, n6225, n6227, n6228_1, n6230,
    n6231, n6232_1, n6233, n6234, n6235, n6236_1, n6237, n6238, n6239,
    n6240_1, n6242, n6243, n6245_1, n6246, n6248, n6249, n6250_1, n6251,
    n6252, n6253, n6254, n6255_1, n6256, n6257, n6258, n6259, n6260_1,
    n6261, n6262, n6263, n6264_1, n6265, n6266, n6267, n6268_1, n6269,
    n6270, n6271, n6272, n6273_1, n6274, n6275, n6276, n6277_1, n6278,
    n6279, n6280, n6281, n6282_1, n6283, n6284, n6285, n6286_1, n6287,
    n6288, n6289, n6290, n6291_1, n6292, n6293, n6294, n6295_1, n6296,
    n6297, n6298, n6299, n6300_1, n6301, n6302, n6303, n6304_1, n6305,
    n6306, n6307, n6308, n6309_1, n6310, n6311, n6312, n6313_1, n6314,
    n6315, n6316, n6317, n6318_1, n6319, n6320, n6321, n6322_1, n6323,
    n6324, n6325, n6326, n6327_1, n6328, n6329, n6330, n6331, n6333, n6334,
    n6336, n6337_1, n6339, n6340, n6341, n6342_1, n6343, n6344, n6345,
    n6347, n6348, n6350_1, n6351, n6353, n6354_1, n6355, n6357, n6358,
    n6360, n6361, n6363, n6364_1, n6365, n6366, n6368, n6369_1, n6371,
    n6372, n6374_1, n6375, n6377, n6378, n6379_1, n6380, n6381, n6383,
    n6384_1, n6385, n6387, n6388_1, n6389, n6391, n6392_1, n6393, n6395,
    n6396_1, n6397, n6399, n6400_1, n6401, n6403, n6404_1, n6405, n6407,
    n6408, n6409_1, n6411, n6412, n6413_1, n6415, n6416, n6417, n6419,
    n6420, n6421, n6422, n6423_1, n6425, n6426, n6427_1, n6429, n6430,
    n6431, n6433, n6434, n6436_1, n6437, n6439, n6440, n6442, n6443, n6445,
    n6446_1, n6448, n6449, n6451_1, n6452, n6454, n6455, n6457, n6458,
    n6460, n6461_1, n6463, n6464, n6466_1, n6467, n6469, n6470, n6472,
    n6473, n6475, n6476_1, n6478, n6479, n6481_1, n6482, n6484, n6485,
    n6487, n6488, n6490, n6491_1, n6493, n6494, n6496_1, n6497, n6499,
    n6500, n6502, n6503, n6505, n6506_1, n6508, n6509, n6511_1, n6512,
    n6514, n6515, n6516_1, n6518, n6519, n6521_1, n6522, n6523, n6525,
    n6526_1, n6528, n6529, n6531_1, n6532, n6534, n6535, n6536_1, n6537,
    n6538, n6539, n6540, n6541_1, n6542, n6543, n6544, n6545, n6546_1,
    n6547, n6548, n6549, n6550, n6551_1, n6552, n6553, n6554, n6555,
    n6556_1, n6557, n6558, n6559, n6560, n6561_1, n6562, n6563, n6564,
    n6565, n6566_1, n6567, n6568, n6569, n6570, n6571_1, n6572, n6573,
    n6574, n6575_1, n6576, n6577, n6578, n6579, n6580_1, n6581, n6582,
    n6583, n6584, n6585_1, n6586, n6587, n6588_1, n6589, n6590, n6591,
    n6592, n6593_1, n6594, n6595, n6596, n6597, n6598_1, n6599, n6600,
    n6601, n6602, n6603_1, n6604, n6605, n6606, n6607, n6608_1, n6609,
    n6610, n6611, n6612, n6613_1, n6614, n6615, n6616, n6617, n6618_1,
    n6619, n6620, n6621, n6622, n6623_1, n6624, n6625, n6626, n6627,
    n6628_1, n6629, n6630, n6631, n6632, n6633_1, n6634, n6635, n6636,
    n6638_1, n6639, n6641, n6642, n6644, n6646, n6648_1, n6650, n6651,
    n6653_1, n6654, n6656, n6657, n6659, n6660, n6662, n6663_1, n6665,
    n6666, n6668_1, n6669, n6671, n6672, n6674, n6675, n6677, n6678_1,
    n6680, n6681, n6683_1, n6684, n6686, n6687, n6689, n6690, n6692,
    n6693_1, n6695, n6696, n6698_1, n6699, n6701, n6702, n6704, n6705,
    n6707, n6708_1, n6710, n6711, n6713_1, n6714, n6716, n6717, n6719,
    n6720, n6722, n6723_1, n6724, n6725, n6726, n6727, n6728_1, n6730,
    n6731, n6733_1, n6734, n6736, n6737, n6738_1, n6739, n6740, n6741,
    n6742, n6744, n6745, n6747, n6748_1, n6750, n6751, n6752, n6753_1,
    n6754, n6756, n6757, n6759, n6760, n6762, n6763_1, n6765, n6766,
    n6768_1, n6769, n6771, n6772, n6774, n6775, n6777, n6778_1, n6780,
    n6781, n6782, n6783_1, n6784, n6785, n6786, n6787, n6789, n6790, n6792,
    n6793_1, n6795, n6796, n6797, n6798_1, n6799, n6800, n6801, n6802,
    n6803_1, n6804, n6805, n6806, n6807, n6808_1, n6809, n6810, n6811,
    n6812, n6813_1, n6814, n6815, n6816, n6817, n6818_1, n6819, n6820,
    n6821, n6822, n6823_1, n6824, n6825, n6826, n6827, n6828_1, n6829,
    n6830, n6831, n6832, n6833_1, n6834, n6835, n6836, n6837, n6838_1,
    n6839, n6840, n6841, n6842, n6843_1, n6844, n6845, n6846, n6847,
    n6848_1, n6849, n6850, n6851, n6852, n6853_1, n6854, n6855, n6856,
    n6857, n6858_1, n6859, n6860, n6861, n6862, n6863_1, n6864, n6865,
    n6866, n6867, n6868_1, n6869, n6870, n6871, n6872, n6873_1, n6874,
    n6875, n6876, n6877, n6878_1, n6879, n6880, n6881, n6882, n6883_1,
    n6884, n6885, n6886, n6887, n6888_1, n6889, n6890, n6891, n6892,
    n6893_1, n6894, n6895, n6896, n6897, n6898_1, n6899, n6900, n6901,
    n6902, n6903_1, n6904, n6905, n6906, n6907, n6908_1, n6909, n6910,
    n6911, n6912, n6913_1, n6914, n6915, n6916, n6917, n6918_1, n6919,
    n6920, n6921, n6922, n6923_1, n6924, n6925, n6926, n6927_1, n6928,
    n6929, n6930, n6931, n6932_1, n6933, n6934, n6935, n6936, n6937_1,
    n6938, n6939, n6940, n6941, n6942_1, n6943, n6944, n6945, n6946,
    n6947_1, n6948, n6949, n6950, n6951, n6952_1, n6953, n6954, n6955,
    n6956, n6957_1, n6958, n6959, n6960, n6961, n6962_1, n6963, n6964,
    n6965, n6966, n6967_1, n6968, n6969, n6970, n6971, n6972_1, n6973,
    n6974, n6975, n6976, n6977_1, n6978, n6979, n6980, n6981, n6982_1,
    n6983, n6984, n6985, n6986, n6987_1, n6988, n6989, n6990, n6991,
    n6992_1, n6993, n6994, n6995, n6996, n6997_1, n6998, n6999, n7000,
    n7001, n7002_1, n7003, n7004, n7005, n7006, n7007_1, n7008, n7009,
    n7010, n7011, n7012_1, n7013, n7014, n7015, n7016, n7017_1, n7018,
    n7019, n7020, n7021, n7022_1, n7023, n7024, n7025, n7026, n7027_1,
    n7028, n7029, n7030, n7031, n7032_1, n7033, n7034, n7035, n7036,
    n7037_1, n7038, n7039, n7040, n7041, n7042_1, n7043, n7044, n7045,
    n7046, n7047_1, n7048, n7049, n7050, n7051, n7052_1, n7053, n7054,
    n7055, n7056, n7057_1, n7058, n7059, n7060, n7061, n7062_1, n7063,
    n7064, n7065, n7066, n7067_1, n7068, n7069, n7071, n7072_1, n7074,
    n7075, n7077_1, n7078, n7079, n7080, n7081, n7082_1, n7083, n7084,
    n7085, n7086, n7087_1, n7088, n7089, n7091, n7092_1, n7094, n7095,
    n7097_1, n7098, n7099, n7100, n7101, n7102_1, n7103, n7104, n7105,
    n7106, n7107_1, n7108, n7109, n7111, n7112_1, n7114, n7115, n7117_1,
    n7118, n7119, n7120, n7121, n7122_1, n7123, n7124, n7125, n7126,
    n7127_1, n7128, n7130, n7131, n7133, n7134, n7136, n7137_1, n7138,
    n7139, n7140, n7141, n7142_1, n7143, n7144, n7145, n7146, n7147_1,
    n7149, n7150, n7152_1, n7153, n7155, n7156, n7157_1, n7158, n7159,
    n7160, n7161_1, n7162, n7163, n7164_1, n7165, n7166, n7168_1, n7169,
    n7171, n7172, n7174, n7175, n7176, n7177_1, n7178, n7179, n7180,
    n7181_1, n7182, n7183, n7184, n7185_1, n7187, n7188, n7190, n7191,
    n7193_1, n7194, n7195, n7196, n7197_1, n7198, n7199, n7200, n7201_1,
    n7202, n7203, n7204, n7206, n7207, n7209, n7210_1, n7212, n7213,
    n7214_1, n7215, n7216, n7217, n7218, n7219_1, n7220, n7221, n7222,
    n7223_1, n7224, n7226, n7227_1, n7229, n7230, n7232, n7233, n7234,
    n7235_1, n7236, n7237, n7238, n7239_1, n7240, n7241, n7242, n7243_1,
    n7245, n7246, n7248, n7249, n7251_1, n7252, n7253, n7255, n7256_1,
    n7257, n7259, n7260, n7261_1, n7263, n7264, n7265, n7267, n7268, n7269,
    n7271, n7272, n7273, n7275, n7276, n7277, n7279, n7280, n7281, n7283,
    n7284, n7285, n7287, n7288, n7289, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
    n7327, n7328, n7329, n7331, n7332, n7333, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7343, n7344, n7346, n7347, n7349, n7350, n7351,
    n7352, n7353, n7354, n7356, n7357, n7359, n7360, n7362, n7363, n7364,
    n7366, n7367, n7369, n7370, n7372, n7373, n7374, n7375, n7376, n7377,
    n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7402, n7403, n7405, n7406, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7415, n7417, n7418, n7420, n7421, n7423, n7424,
    n7425, n7426, n7428, n7429, n7430, n7432, n7433, n7434, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7453, n7454, n7456, n7457, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7482, n7483, n7485, n7486, n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7497, n7498, n7499, n7501, n7502, n7503, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7513, n7514, n7516, n7517, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7545, n7546, n7548, n7549, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7563,
    n7564, n7566, n7567, n7569, n7570, n7571, n7572, n7573, n7575, n7576,
    n7577, n7579, n7580, n7581, n7583, n7584, n7585, n7587, n7588, n7590,
    n7591, n7593, n7594, n7595, n7596, n7597, n7599, n7600, n7601, n7602,
    n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
    n7633, n7634, n7635, n7636, n7637, n7638, n7640, n7642, n7643, n7645,
    n7646, n7648, n7649, n7650, n7651, n7653, n7654, n7656, n7657, n7659,
    n7660, n7662, n7663, n7665, n7666, n7668, n7669, n7671, n7672, n7674,
    n7675, n7677, n7678, n7680, n7681, n7683, n7684, n7686, n7687, n7689,
    n7690, n7692, n7693, n7695, n7696, n7698, n7699, n7700, n7701, n7703,
    n7704, n7705, n7706, n7708, n7709, n7710, n7711, n7713, n7714, n7715,
    n7716, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
    n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
    n7769, n7770, n7771, n7773, n7774, n7775, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7785, n7786, n7788, n7789, n7791, n7792, n7793,
    n7794, n7795, n7796, n7798, n7799, n7801, n7802, n7804, n7805, n7806,
    n7807, n7809, n7810, n7812, n7813, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7827, n7828, n7830, n7831,
    n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7845, n7846, n7848, n7849, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
    n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
    n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
    n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7936,
    n7937, n7939, n7940, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7950, n7951, n7953, n7954, n7956, n7957, n7958, n7960, n7961, n7963,
    n7964, n7966, n7967, n7968, n7969, n7971, n7972, n7974, n7975, n7977,
    n7979, n7980, n7981, n7982, n7983, n7985, n7986, n7987, n7989, n7990,
    n7991, n7993, n7994, n7995, n7997, n7998, n7999, n8001, n8002, n8003,
    n8005, n8006, n8007, n8009, n8010, n8011, n8013, n8014, n8015, n8017,
    n8018, n8019, n8021, n8022, n8023, n8024, n8025, n8027, n8028, n8029,
    n8031, n8032, n8033, n8035, n8036, n8038, n8039, n8041, n8042, n8044,
    n8045, n8047, n8048, n8050, n8051, n8053, n8054, n8056, n8057, n8059,
    n8060, n8062, n8063, n8065, n8066, n8068, n8069, n8071, n8072, n8074,
    n8075, n8077, n8078, n8080, n8081, n8083, n8084, n8086, n8087, n8089,
    n8090, n8092, n8093, n8095, n8096, n8098, n8099, n8101, n8102, n8104,
    n8105, n8107, n8108, n8110, n8111, n8113, n8114, n8116, n8117, n8118,
    n8120, n8121, n8123, n8124, n8125, n8127, n8128, n8130, n8131, n8133,
    n8134, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8240, n8241, n8243, n8244, n8246, n8248,
    n8250, n8252, n8253, n8255, n8256, n8258, n8259, n8261, n8262, n8264,
    n8265, n8267, n8268, n8270, n8271, n8273, n8274, n8276, n8277, n8279,
    n8280, n8282, n8283, n8285, n8286, n8288, n8289, n8291, n8292, n8294,
    n8295, n8297, n8298, n8300, n8301, n8303, n8304, n8306, n8307, n8309,
    n8310, n8312, n8313, n8315, n8316, n8318, n8319, n8321, n8322, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330, n8332, n8333, n8335, n8336,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8349,
    n8350, n8352, n8353, n8354, n8355, n8356, n8358, n8359, n8361, n8362,
    n8364, n8365, n8367, n8368, n8370, n8371, n8373, n8374, n8376, n8377,
    n8379, n8380, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8391, n8392, n8394, n8395, n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8669, n8670, n8672, n8673, n8675,
    n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
    n8686, n8687, n8689, n8690, n8692, n8693, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8709,
    n8710, n8712, n8713, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
    n8722, n8723, n8724, n8725, n8726, n8728, n8729, n8731, n8732, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8747, n8748, n8750, n8751, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8766, n8767, n8769,
    n8770, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8785, n8786, n8788, n8789, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8804,
    n8805, n8807, n8808, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822, n8824, n8825, n8827, n8828,
    n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8843, n8844, n8846, n8847, n8849, n8850, n8851, n8853,
    n8854, n8855, n8857, n8858, n8859, n8861, n8862, n8863, n8865, n8866,
    n8867, n8869, n8870, n8871, n8873, n8874, n8875, n8877, n8878, n8879,
    n8881, n8882, n8883, n8885, n8886, n8887, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8925, n8926, n8927, n8929, n8930, n8931, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8941, n8942, n8944, n8945, n8947, n8948,
    n8949, n8950, n8951, n8952, n8954, n8955, n8957, n8958, n8960, n8961,
    n8962, n8964, n8965, n8967, n8968, n8970, n8971, n8972, n8973, n8974,
    n8975, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n9000, n9001, n9003, n9004, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9015, n9016, n9018, n9019, n9021,
    n9022, n9023, n9024, n9026, n9027, n9028, n9030, n9031, n9032, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9051, n9052, n9054, n9055, n9057,
    n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9080, n9081, n9083, n9084, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9095, n9096, n9097, n9099, n9100, n9101, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109, n9111, n9112, n9114, n9115,
    n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9143, n9144, n9146, n9147, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9161, n9162, n9164, n9165, n9167, n9168, n9169, n9170, n9171, n9173,
    n9174, n9175, n9177, n9178, n9179, n9181, n9182, n9183, n9185, n9186,
    n9188, n9189, n9191, n9192, n9193, n9194, n9195, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9238, n9240, n9241,
    n9243, n9244, n9246, n9247, n9248, n9249, n9251, n9252, n9254, n9255,
    n9257, n9258, n9260, n9261, n9263, n9264, n9266, n9267, n9269, n9270,
    n9272, n9273, n9275, n9276, n9278, n9279, n9281, n9282, n9284, n9285,
    n9287, n9288, n9290, n9291, n9293, n9294, n9296, n9297, n9298, n9299,
    n9301, n9302, n9303, n9304, n9306, n9307, n9308, n9309, n9311, n9312,
    n9313, n9314, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9367, n9368, n9369, n9371, n9372, n9373, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9383, n9384, n9386, n9387, n9389, n9390,
    n9391, n9392, n9393, n9394, n9396, n9397, n9399, n9400, n9402, n9403,
    n9404, n9405, n9407, n9408, n9410, n9411, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9425, n9426, n9428,
    n9429, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9443, n9444, n9446, n9447, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
    n9534, n9535, n9537, n9538, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9548, n9549, n9551, n9552, n9554, n9555, n9556, n9558, n9559,
    n9561, n9562, n9564, n9565, n9566, n9567, n9568, n9570, n9571, n9573,
    n9574, n9576, n9578, n9579, n9580, n9581, n9582, n9584, n9585, n9586,
    n9588, n9589, n9590, n9592, n9593, n9594, n9596, n9597, n9598, n9600,
    n9601, n9602, n9604, n9605, n9606, n9608, n9609, n9610, n9612, n9613,
    n9614, n9616, n9617, n9618, n9620, n9621, n9622, n9623, n9624, n9626,
    n9627, n9628, n9630, n9631, n9632, n9634, n9635, n9637, n9638, n9640,
    n9641, n9643, n9644, n9646, n9647, n9649, n9650, n9652, n9653, n9655,
    n9656, n9658, n9659, n9661, n9662, n9664, n9665, n9667, n9668, n9670,
    n9671, n9673, n9674, n9676, n9677, n9679, n9680, n9682, n9683, n9685,
    n9686, n9688, n9689, n9691, n9692, n9694, n9695, n9697, n9698, n9700,
    n9701, n9703, n9704, n9706, n9707, n9709, n9710, n9712, n9713, n9715,
    n9716, n9717, n9719, n9720, n9722, n9723, n9724, n9726, n9727, n9729,
    n9730, n9732, n9733, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
    n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837, n9839, n9840, n9842, n9843,
    n9845, n9847, n9849, n9851, n9852, n9854, n9855, n9857, n9858, n9860,
    n9861, n9863, n9864, n9866, n9867, n9869, n9870, n9872, n9873, n9875,
    n9876, n9878, n9879, n9881, n9882, n9884, n9885, n9887, n9888, n9890,
    n9891, n9893, n9894, n9896, n9897, n9899, n9900, n9902, n9903, n9905,
    n9906, n9908, n9909, n9911, n9912, n9914, n9915, n9917, n9918, n9920,
    n9921, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9931, n9932,
    n9934, n9935, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9945,
    n9946, n9948, n9949, n9951, n9952, n9953, n9954, n9955, n9957, n9958,
    n9960, n9961, n9963, n9964, n9966, n9967, n9969, n9970, n9972, n9973,
    n9975, n9976, n9978, n9979, n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9990, n9991, n9993, n9994, n9996, n9997, n9998, n9999,
    n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
    n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
    n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
    n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
    n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
    n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
    n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10270,
    n10271, n10273, n10274, n10276, n10277, n10278, n10279, n10280, n10281,
    n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10290, n10291,
    n10293, n10294, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308, n10310, n10311, n10313,
    n10314, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10325, n10326, n10327, n10329, n10330, n10332, n10333, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10348, n10349, n10351, n10352, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
    n10367, n10368, n10370, n10371, n10373, n10374, n10375, n10376, n10377,
    n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10386, n10387,
    n10389, n10390, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10405, n10406, n10408, n10409,
    n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10425, n10426, n10428, n10429, n10431,
    n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10444, n10445, n10447, n10448, n10450, n10451, n10452,
    n10454, n10455, n10456, n10458, n10459, n10460, n10462, n10463, n10464,
    n10466, n10467, n10468, n10470, n10471, n10472, n10474, n10475, n10476,
    n10478, n10479, n10480, n10482, n10483, n10484, n10486, n10487, n10488,
    n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10526,
    n10527, n10528, n10530, n10531, n10532, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10542, n10543, n10545, n10546, n10548, n10549,
    n10550, n10551, n10552, n10553, n10555, n10556, n10558, n10559, n10561,
    n10562, n10563, n10565, n10566, n10568, n10569, n10571, n10572, n10573,
    n10574, n10575, n10576, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10601, n10602,
    n10604, n10605, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10616, n10617, n10619, n10620, n10622, n10623, n10624, n10625,
    n10627, n10628, n10629, n10631, n10632, n10633, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10652, n10653, n10655, n10656, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10681, n10682, n10684, n10685, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10696, n10697, n10698,
    n10700, n10701, n10702, n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10712, n10713, n10715, n10716, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10744, n10745, n10747, n10748, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
    n10762, n10763, n10765, n10766, n10768, n10769, n10770, n10771, n10772,
    n10774, n10775, n10776, n10778, n10779, n10780, n10782, n10783, n10784,
    n10786, n10787, n10789, n10790, n10792, n10793, n10794, n10795, n10796,
    n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10839, n10841, n10842, n10844, n10845,
    n10847, n10848, n10849, n10850, n10852, n10853, n10855, n10856, n10858,
    n10859, n10861, n10862, n10864, n10865, n10867, n10868, n10870, n10871,
    n10873, n10874, n10876, n10877, n10879, n10880, n10882, n10883, n10885,
    n10886, n10888, n10889, n10891, n10892, n10894, n10895, n10897, n10898,
    n10899, n10900, n10902, n10903, n10904, n10905, n10907, n10908, n10909,
    n10910, n10912, n10913, n10914, n10915, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10968, n10969, n10970, n10972, n10973, n10974, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10984, n10985, n10987, n10988, n10990,
    n10991, n10992, n10993, n10994, n10995, n10997, n10998, n11000, n11001,
    n11003, n11004, n11005, n11006, n11008, n11009, n11011, n11012, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11026, n11027, n11029, n11030, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11044, n11045,
    n11047, n11048, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
    n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11135, n11136, n11138, n11139,
    n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11149, n11150,
    n11152, n11153, n11155, n11156, n11157, n11159, n11160, n11162, n11163,
    n11165, n11166, n11167, n11168, n11169, n11171, n11172, n11174, n11175,
    n11177, n11179, n11180, n11181, n11182, n11183, n11185, n11186, n11187,
    n11189, n11190, n11191, n11193, n11194, n11195, n11197, n11198, n11199,
    n11201, n11202, n11203, n11205, n11206, n11207, n11209, n11210, n11211,
    n11213, n11214, n11215, n11217, n11218, n11219, n11221, n11222, n11223,
    n11224, n11225, n11227, n11228, n11229, n11231, n11232, n11233, n11235,
    n11236, n11238, n11239, n11241, n11242, n11244, n11245, n11247, n11248,
    n11250, n11251, n11253, n11254, n11256, n11257, n11259, n11260, n11262,
    n11263, n11265, n11266, n11268, n11269, n11271, n11272, n11274, n11275,
    n11277, n11278, n11280, n11281, n11283, n11284, n11286, n11287, n11289,
    n11290, n11292, n11293, n11295, n11296, n11298, n11299, n11301, n11302,
    n11304, n11305, n11307, n11308, n11310, n11311, n11313, n11314, n11316,
    n11317, n11318, n11320, n11321, n11323, n11324, n11325, n11327, n11328,
    n11330, n11331, n11333, n11334, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11440,
    n11441, n11443, n11444, n11446, n11448, n11450, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
    n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
    n11494, n11495, n11496, n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11540, n11541, n11542, n11543,
    n11544, n11545, n11546, n11547, n11548, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
    n11676, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
    n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
    n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
    n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11771, n11772,
    n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
    n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
    n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
    n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
    n11809, n11810, n11811, n11812, n11813, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834, n11836, n11837, n11838,
    n11839, n11840, n11841, n11842, n11843, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11866, n11867, n11868,
    n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
    n11878, n11879, n11880, n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
    n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11930, n11931, n11932, n11933, n11934,
    n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
    n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
    n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
    n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
    n11971, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
    n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12087,
    n12088, n12089, n12091, n12092, n12093, n12094, n12095, n12097, n12098,
    n12099, n12100, n12102, n12103, n12104, n12106, n12107, n12108, n12110,
    n12111, n12112, n12114, n12115, n12116, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12126, n12127, n12128, n12130, n12131, n12132,
    n12134, n12135, n12136, n12138, n12139, n12141, n12142, n12144, n12145,
    n12147, n12148, n12150, n12151, n12153, n12154, n12156, n12157, n12159,
    n12160, n12162, n12163, n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
    n12190, n12191, n12193, n12194, n12196, n12197, n12199, n12200, n12202,
    n12203, n12205, n12206, n12208, n12209, n12211, n12212, n12214, n12215,
    n12217, n12218, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12244, n12245,
    n271_1, n275_1, n280, n285_1, n290_1, n295_1, n300_1, n305_1, n310_1,
    n315, n320_1, n325_1, n330_1, n335_1, n340_1, n345_1, n350_1, n354_1,
    n359_1, n363_1, n367_1, n371_1, n375_1, n379_1, n383_1, n387_1, n391_1,
    n395_1, n399_1, n403_1, n407_1, n411_1, n415, n419_1, n423_1, n427,
    n431_1, n436, n441_1, n446_1, n451, n456, n461_1, n466_1, n471_1,
    n476_1, n481, n484, n489, n492_1, n497_1, n500, n505_1, n508_1, n513_1,
    n516_1, n521_1, n524_1, n529_1, n532_1, n537_1, n540_1, n545_1, n548_1,
    n553_1, n556_1, n561_1, n564_1, n569_1, n572_1, n577_1, n580_1, n585_1,
    n588, n593, n596_1, n601_1, n604_1, n609_1, n612_1, n617_1, n620_1,
    n625_1, n630, n635_1, n640_1, n645_1, n650, n655, n660, n665_1, n670,
    n675_1, n680, n685_1, n690, n695_1, n700_1, n705_1, n710_1, n715_1,
    n720, n725, n730_1, n735_1, n740_1, n745_1, n750_1, n755_1, n760_1,
    n765_1, n770_1, n775_1, n780_1, n785_1, n790_1, n795_1, n800_1, n805_1,
    n810_1, n815_1, n820, n825_1, n830_1, n835_1, n840_1, n845_1, n849_1,
    n854_1, n859_1, n864_1, n869_1, n873_1, n877_1, n881_1, n885_1, n889_1,
    n894_1, n899_1, n904_1, n909_1, n914_1, n919_1, n924_1, n929_1, n934,
    n939_1, n944_1, n949_1, n954_1, n959_1, n964_1, n969_1, n974_1, n979_1,
    n984_1, n989_1, n994_1, n999_1, n1004_1, n1009_1, n1014, n1019_1,
    n1024_1, n1029, n1034_1, n1039_1, n1044, n1049, n1054_1, n1059_1,
    n1064_1, n1069, n1074_1, n1079, n1084_1, n1089_1, n1094_1, n1099_1,
    n1104_1, n1109_1, n1114, n1119_1, n1124_1, n1129_1, n1134_1, n1139_1,
    n1144_1, n1149_1, n1154_1, n1159_1, n1164, n1169_1, n1174_1, n1179_1,
    n1184_1, n1189_1, n1194, n1199_1, n1204_1, n1209_1, n1214_1, n1219_1,
    n1224_1, n1229_1, n1234_1, n1239_1, n1244_1, n1249_1, n1254_1, n1259_1,
    n1264_1, n1269, n1274, n1279, n1284_1, n1289, n1294, n1299, n1304,
    n1309, n1314_1, n1319, n1324_1, n1329_1, n1334_1, n1339_1, n1344_1,
    n1349_1, n1354, n1359, n1364, n1369, n1374_1, n1379, n1384_1, n1389_1,
    n1394_1, n1399_1, n1404_1, n1409_1, n1414, n1419, n1424_1, n1429_1,
    n1434, n1439_1, n1444_1, n1449, n1454, n1459_1, n1464, n1469_1,
    n1474_1, n1479_1, n1484_1, n1489, n1494_1, n1499, n1504, n1509_1,
    n1514_1, n1519_1, n1524_1, n1529_1, n1534, n1538_1, n1543, n1547_1,
    n1552_1, n1556_1, n1561_1, n1565_1, n1570_1, n1574, n1579_1, n1583,
    n1588, n1592, n1597_1, n1601, n1605_1, n1609_1, n1614_1, n1619_1,
    n1624_1, n1628_1, n1632, n1636_1, n1640_1, n1644_1, n1648_1, n1652_1,
    n1656_1, n1660, n1664_1, n1668, n1672, n1676_1, n1680, n1684, n1688_1,
    n1692_1, n1696_1, n1700_1, n1704_1, n1708, n1712, n1716_1, n1720_1,
    n1725, n1730, n1735_1, n1740, n1744_1, n1748, n1753_1, n1757_1,
    n1762_1, n1766_1, n1771_1, n1775_1, n1780_1, n1784_1, n1789_1, n1793,
    n1798, n1802_1, n1807_1, n1812_1, n1817_1, n1822_1, n1826_1, n1830_1,
    n1834_1, n1839, n1844_1, n1849_1, n1854, n1859_1, n1864_1, n1868_1,
    n1872_1, n1876_1, n1880_1, n1884_1, n1889_1, n1893_1, n1898_1, n1903,
    n1907_1, n1912_1, n1916_1, n1921, n1926_1, n1931, n1936_1, n1941_1,
    n1946_1, n1951_1, n1956_1, n1961, n1966_1, n1971, n1976_1, n1981,
    n1986, n1991_1, n1996_1, n2001, n2006_1, n2011_1, n2016, n2021_1,
    n2026_1, n2031_1, n2036_1, n2041_1, n2046, n2051_1, n2055_1, n2060_1,
    n2065, n2068_1, n2073, n2078_1, n2083_1, n2088_1, n2093_1, n2098,
    n2103, n2108_1, n2113_1, n2118, n2123_1, n2128, n2133, n2138_1,
    n2143_1, n2148_1, n2153_1, n2158_1, n2163_1, n2168_1, n2173_1, n2178_1,
    n2183_1, n2188, n2193, n2198_1, n2203_1, n2208_1, n2213, n2218,
    n2223_1, n2228, n2233_1, n2238, n2243_1, n2248, n2253_1, n2258, n2263,
    n2268, n2273, n2278_1, n2283, n2288, n2293, n2298, n2303, n2308, n2313,
    n2318, n2323_1, n2328, n2333, n2338, n2343, n2348, n2353, n2358_1,
    n2363, n2368, n2373, n2378, n2383, n2388, n2392, n2396_1, n2400_1,
    n2405, n2410, n2415, n2420, n2425_1, n2430_1, n2435, n2440, n2445,
    n2450_1, n2455_1, n2460_1, n2465, n2470, n2475, n2480, n2485, n2490,
    n2495_1, n2500_1, n2505_1, n2510_1, n2515_1, n2520_1, n2525, n2530,
    n2535, n2540, n2545_1, n2550, n2555, n2560_1, n2565, n2570, n2575_1,
    n2580, n2585, n2590, n2595_1, n2600, n2605, n2610, n2615, n2620_1,
    n2625, n2630, n2635, n2640, n2645, n2650, n2655, n2660, n2665, n2670,
    n2675, n2680_1, n2685, n2690, n2695_1, n2700, n2705_1, n2710_1,
    n2715_1, n2720, n2725_1, n2730_1, n2735_1, n2740_1, n2745_1, n2750_1,
    n2755_1, n2760_1, n2765_1, n2770_1, n2775_1, n2780_1, n2785_1, n2790_1,
    n2795_1, n2800_1, n2805_1, n2810_1, n2815_1, n2820_1, n2825_1, n2830_1,
    n2835, n2840_1, n2845_1, n2850_1, n2855_1, n2860_1, n2865_1, n2870_1,
    n2875_1, n2880_1, n2885_1, n2890_1, n2895_1, n2900_1, n2905_1, n2910_1,
    n2915_1, n2920_1, n2925_1, n2930_1, n2935_1, n2940_1, n2945_1, n2950_1,
    n2955_1, n2960_1, n2965_1, n2970_1, n2975_1, n2980_1, n2985_1, n2990_1,
    n2995_1, n3000_1, n3005_1, n3010_1, n3015, n3020_1, n3025, n3030_1,
    n3035_1, n3040, n3044_1, n3049_1, n3053_1, n3058_1, n3062_1, n3067_1,
    n3071_1, n3076_1, n3080_1, n3085_1, n3089_1, n3094_1, n3098_1, n3103_1,
    n3107, n3111_1, n3115_1, n3120_1, n3125_1, n3130_1, n3134, n3138_1,
    n3142_1, n3146_1, n3150, n3154_1, n3158_1, n3162_1, n3166, n3170_1,
    n3174_1, n3178_1, n3182_1, n3186_1, n3190_1, n3194_1, n3198_1, n3202_1,
    n3206_1, n3210_1, n3214_1, n3218_1, n3222_1, n3226_1, n3231_1, n3236_1,
    n3241_1, n3246_1, n3250_1, n3254_1, n3259_1, n3263_1, n3268_1, n3272_1,
    n3277_1, n3281_1, n3286_1, n3290_1, n3295_1, n3299_1, n3304_1, n3308_1,
    n3313_1, n3318_1, n3323_1, n3328_1, n3332_1, n3336_1, n3340_1, n3345_1,
    n3350_1, n3355_1, n3360_1, n3365_1, n3370_1, n3374_1, n3378_1, n3382_1,
    n3386_1, n3390_1, n3395_1, n3399_1, n3404_1, n3409_1, n3413_1, n3418_1,
    n3422_1, n3427_1, n3432_1, n3437_1, n3442_1, n3447_1, n3452_1, n3457_1,
    n3462_1, n3467_1, n3472_1, n3477_1, n3482_1, n3487_1, n3492_1, n3497_1,
    n3502_1, n3507_1, n3512_1, n3517_1, n3522_1, n3527_1, n3532_1, n3537_1,
    n3542_1, n3547_1, n3552_1, n3557_1, n3561_1, n3566_1, n3571_1, n3574_1,
    n3579_1, n3584_1, n3589_1, n3594_1, n3599_1, n3604_1, n3609_1, n3614_1,
    n3619_1, n3624_1, n3629_1, n3633_1, n3637_1, n3642_1, n3647_1, n3652_1,
    n3657_1, n3662_1, n3667_1, n3672_1, n3677_1, n3682_1, n3687_1, n3692_1,
    n3697_1, n3702_1, n3707_1, n3712_1, n3717_1, n3722_1, n3727_1, n3732_1,
    n3737_1, n3742_1, n3747, n3752_1, n3757, n3762_1, n3767, n3772_1,
    n3777, n3782, n3787_1, n3792_1, n3797, n3802_1, n3807_1, n3812, n3817,
    n3822_1, n3827, n3832_1, n3837, n3842_1, n3847_1, n3852_1, n3857_1,
    n3862_1, n3867, n3872_1, n3877_1, n3882, n3887, n3892_1, n3897_1,
    n3902, n3907_1, n3912_1, n3917, n3922, n3927, n3932_1, n3937, n3942_1,
    n3947, n3952, n3957_1, n3962, n3967, n3972, n3977, n3982, n3987, n3992,
    n3997_1, n4002_1, n4007_1, n4012, n4017, n4022_1, n4027, n4032_1,
    n4037_1, n4042, n4047, n4052, n4057_1, n4062_1, n4067, n4072_1, n4077,
    n4082, n4087, n4092, n4097, n4102_1, n4107_1, n4112_1, n4117, n4122_1,
    n4127_1, n4132_1, n4137_1, n4142_1, n4147_1, n4152, n4157, n4162,
    n4167_1, n4172, n4177, n4182, n4187_1, n4192, n4197_1, n4202, n4207,
    n4212_1, n4217_1, n4222, n4227, n4232, n4237, n4242, n4247, n4252_1,
    n4257_1, n4262, n4267, n4272, n4277, n4282, n4287, n4292, n4297, n4302,
    n4307, n4312, n4317, n4322_1, n4327, n4332_1, n4337_1, n4342, n4347_1,
    n4352_1, n4357_1, n4362_1, n4367, n4372, n4377, n4382, n4387, n4392,
    n4397, n4402, n4407, n4412, n4417, n4422, n4427, n4432, n4437, n4442_1,
    n4447_1, n4452_1, n4457, n4462, n4467, n4472, n4477, n4482, n4487,
    n4492, n4497, n4502, n4507, n4512, n4517, n4522, n4527, n4532, n4537,
    n4542, n4547, n4551, n4556, n4560, n4565, n4569, n4574, n4578, n4583,
    n4587, n4592, n4596, n4601, n4605, n4610, n4614, n4618, n4622, n4627,
    n4632, n4637, n4641, n4645, n4649, n4653, n4657, n4661, n4665, n4669,
    n4673, n4677, n4681, n4685, n4689, n4693, n4697, n4701, n4705, n4709,
    n4713, n4717, n4721, n4725, n4729, n4733, n4738, n4743, n4748, n4753,
    n4757, n4761, n4766, n4770, n4775, n4779, n4784, n4788, n4793, n4797,
    n4802, n4806, n4811, n4815, n4820, n4825, n4830, n4835, n4839, n4843,
    n4847, n4852, n4857, n4862, n4867, n4872_1, n4877, n4881, n4885, n4889,
    n4893_1, n4897_1, n4902, n4906_1, n4911, n4916, n4920, n4925, n4929,
    n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979,
    n4984, n4989, n4994, n4999, n5004, n5009, n5014, n5019, n5024, n5029,
    n5034, n5039, n5044, n5049, n5054, n5059, n5064, n5068, n5073, n5078,
    n5081, n5086, n5091, n5096, n5101, n5106, n5111, n5116, n5121, n5126,
    n5131, n5136, n5141, n5146, n5151, n5156, n5161, n5166, n5171, n5176,
    n5181, n5186, n5191, n5196, n5201, n5206, n5211, n5216, n5221, n5226,
    n5231, n5236, n5241, n5246, n5251, n5256, n5261, n5266, n5271, n5276,
    n5281, n5286, n5291, n5296, n5301, n5306, n5311, n5316, n5321, n5326,
    n5331, n5336, n5341, n5346, n5351, n5356, n5361, n5366, n5371, n5376,
    n5381, n5386, n5391, n5396, n5401, n5406, n5411, n5416, n5421, n5426,
    n5431, n5436, n5441, n5446, n5451, n5456, n5461, n5466, n5471, n5476,
    n5481, n5486, n5491, n5496, n5501, n5506, n5511, n5516, n5521, n5526,
    n5531, n5536, n5541, n5546, n5551, n5556, n5561, n5566, n5571, n5576,
    n5581, n5586, n5591, n5596, n5601, n5606, n5611, n5616, n5621, n5626,
    n5631, n5636, n5641, n5646, n5651, n5656, n5661, n5666, n5671, n5676,
    n5681, n5686, n5691, n5696, n5701, n5706, n5711, n5716, n5721, n5726,
    n5731, n5736, n5741, n5746, n5751, n5756, n5761, n5766, n5771, n5776,
    n5781, n5786, n5791, n5796, n5801, n5806, n5811, n5816, n5820, n5824,
    n5829, n5834, n5839, n5844, n5849, n5854, n5859, n5864, n5869, n5874,
    n5879, n5884, n5889, n5894, n5899, n5904, n5909, n5914, n5919, n5924,
    n5929, n5934, n5939, n5944, n5949, n5954, n5959, n5964, n5969, n5974,
    n5979, n5984, n5989, n5994, n5999, n6004, n6009, n6014, n6019, n6024,
    n6029, n6034, n6039, n6044, n6049, n6054, n6058, n6063, n6067, n6072,
    n6076, n6081, n6085, n6090, n6094, n6099, n6103, n6108, n6112, n6117,
    n6121, n6125, n6129, n6134, n6139, n6144, n6148, n6152, n6156, n6160,
    n6164, n6168, n6172, n6176, n6180, n6184, n6188, n6192, n6196, n6200,
    n6204, n6208, n6212, n6216, n6220, n6224, n6228, n6232, n6236, n6240,
    n6245, n6250, n6255, n6260, n6264, n6268, n6273, n6277, n6282, n6286,
    n6291, n6295, n6300, n6304, n6309, n6313, n6318, n6322, n6327, n6332,
    n6337, n6342, n6346, n6350, n6354, n6359, n6364, n6369, n6374, n6379,
    n6384, n6388, n6392, n6396, n6400, n6404, n6409, n6413, n6418, n6423,
    n6427, n6432, n6436, n6441, n6446, n6451, n6456, n6461, n6466, n6471,
    n6476, n6481, n6486, n6491, n6496, n6501, n6506, n6511, n6516, n6521,
    n6526, n6531, n6536, n6541, n6546, n6551, n6556, n6561, n6566, n6571,
    n6575, n6580, n6585, n6588, n6593, n6598, n6603, n6608, n6613, n6618,
    n6623, n6628, n6633, n6638, n6643, n6648, n6653, n6658, n6663, n6668,
    n6673, n6678, n6683, n6688, n6693, n6698, n6703, n6708, n6713, n6718,
    n6723, n6728, n6733, n6738, n6743, n6748, n6753, n6758, n6763, n6768,
    n6773, n6778, n6783, n6788, n6793, n6798, n6803, n6808, n6813, n6818,
    n6823, n6828, n6833, n6838, n6843, n6848, n6853, n6858, n6863, n6868,
    n6873, n6878, n6883, n6888, n6893, n6898, n6903, n6908, n6913, n6918,
    n6923, n6927, n6932, n6937, n6942, n6947, n6952, n6957, n6962, n6967,
    n6972, n6977, n6982, n6987, n6992, n6997, n7002, n7007, n7012, n7017,
    n7022, n7027, n7032, n7037, n7042, n7047, n7052, n7057, n7062, n7067,
    n7072, n7077, n7082, n7087, n7092, n7097, n7102, n7107, n7112, n7117,
    n7122, n7127, n7132, n7137, n7142, n7147, n7152, n7157, n7161, n7164,
    n7168, n7173, n7177, n7181, n7185, n7189, n7193, n7197, n7201, n7205,
    n7210, n7214, n7219, n7223, n7227, n7231, n7235, n7239, n7243, n7247,
    n7251, n7256, n7261;
  assign n4522_1 = ~Ng3191 & ~Ng3126;
  assign n4523 = ~Ng3110 & n4522_1;
  assign n4524 = ~Ng3147 & n4523;
  assign n4525 = Ng3120 & ~Ng3139;
  assign n4526 = Ng3135 & n4525;
  assign n4527_1 = n4524 & n4526;
  assign n4528 = ~Ng185 & n4527_1;
  assign n4529 = ~Ng2992 & ~Ng2991;
  assign n4530 = ~Ng3139 & ~n4529;
  assign n4531 = Ng3110 & n4522_1;
  assign n4532_1 = Ng3147 & n4531;
  assign n4533 = ~n4530 & n4532_1;
  assign n4534 = ~n4524 & ~n4533;
  assign n4535 = ~Ng3120 & Ng3135;
  assign n4536 = ~n4534 & n4535;
  assign n4537_1 = ~n4528 & ~n4536;
  assign n4538 = Ng185 & ~n4524;
  assign n4539 = Ng3139 & n4538;
  assign n4540 = ~n4537_1 & ~n4539;
  assign n4541 = ~Ng3120 & ~Ng3139;
  assign n4542_1 = ~Ng3135 & n4524;
  assign n4543 = n4541 & n4542_1;
  assign Pg25442 = ~Pg3233 | Pg3230;
  assign n4545 = ~n4543 & ~Pg25442;
  assign n894_1 = ~n4540 & n4545;
  assign n4547_1 = ~Ng3135 & n4532_1;
  assign n4548 = n4541 & n4547_1;
  assign n4549 = Ng3167 & n4548;
  assign n4550 = ~Ng3120 & Ng3139;
  assign n4551_1 = n4547_1 & n4550;
  assign n4552 = Ng3170 & n4551_1;
  assign n4553 = ~n4549 & ~n4552;
  assign n4554 = Ng3147 & n4523;
  assign n4555 = n4541 & n4554;
  assign n4556_1 = Ng3135 & n4555;
  assign n4557 = ~n4527_1 & ~n4556_1;
  assign n4558 = n4553 & n4557;
  assign n4559 = ~Ng3147 & n4531;
  assign n4560_1 = ~Ng3135 & n4559;
  assign n4561 = n4525 & n4560_1;
  assign n4562 = Ng3161 & n4561;
  assign n4563 = Ng3135 & n4559;
  assign n4564 = Ng3120 & Ng3139;
  assign n4565_1 = n4563 & n4564;
  assign n4566 = Ng3088 & n4565_1;
  assign n4567 = ~n4562 & ~n4566;
  assign n4568 = n4525 & n4547_1;
  assign n4569_1 = Ng3173 & n4568;
  assign n4570 = n4567 & ~n4569_1;
  assign n4571 = n4558 & n4570;
  assign n4572 = n4541 & n4560_1;
  assign n4573 = Ng3155 & n4572;
  assign n4574_1 = n4526 & n4559;
  assign n4575 = Ng3185 & n4574_1;
  assign n4576 = ~Pg25442 & ~n4575;
  assign n4577 = ~n4573 & n4576;
  assign n4578_1 = n4550 & n4560_1;
  assign n4579 = Ng3158 & n4578_1;
  assign n4580 = n4577 & ~n4579;
  assign n4581 = n4550 & n4563;
  assign n4582 = Ng3182 & n4581;
  assign n4583_1 = n4560_1 & n4564;
  assign n4584 = Ng3164 & n4583_1;
  assign n4585 = ~n4582 & ~n4584;
  assign n4586 = n4541 & n4563;
  assign n4587_1 = Ng3179 & n4586;
  assign n4588 = n4547_1 & n4564;
  assign n4589 = Ng3176 & n4588;
  assign n4590 = ~n4587_1 & ~n4589;
  assign n4591 = n4585 & n4590;
  assign n4592_1 = n4580 & n4591;
  assign Pg26149 = ~n4571 | ~n4592_1;
  assign n4594 = Ng3102 & n4551_1;
  assign n4595 = Ng3106 & n4581;
  assign n4596_1 = ~n4529 & n4543;
  assign n4597 = ~n4595 & ~n4596_1;
  assign n4598 = ~n4594 & n4597;
  assign n4599 = Ng3098 & n4578_1;
  assign n4600 = ~Ng3128 & n4527_1;
  assign n4601_1 = ~n4599 & ~n4600;
  assign n4602 = Ng3107 & n4574_1;
  assign n4603 = ~Pg25442 & ~n4602;
  assign n4604 = Ng3099 & n4561;
  assign n4605_1 = n4603 & ~n4604;
  assign n4606 = n4601_1 & n4605_1;
  assign n4607 = Ng3105 & n4586;
  assign n4608 = n4526 & n4554;
  assign n4609 = ~n4555 & ~n4608;
  assign n4610_1 = ~n4607 & n4609;
  assign n4611 = n4606 & n4610_1;
  assign n4612 = n4598 & n4611;
  assign n4613 = Ng3103 & n4568;
  assign n4614_1 = Ng3097 & n4572;
  assign n4615 = Ng3101 & n4548;
  assign n4616 = Ng3104 & n4588;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618_1 = Ng3100 & n4583_1;
  assign n4619 = Ng3108 & n4565_1;
  assign n4620 = ~n4618_1 & ~n4619;
  assign n4621 = n4617 & n4620;
  assign n4622_1 = ~n4614_1 & n4621;
  assign n4623 = ~n4613 & n4622_1;
  assign n854_1 = n4612 & n4623;
  assign n4625 = Ng3092 & n4588;
  assign n4626 = Ng3086 & n4548;
  assign n4627_1 = Ng3084 & n4561;
  assign n4628 = ~n4626 & ~n4627_1;
  assign n4629 = Ng3094 & n4581;
  assign n4630 = n4628 & ~n4629;
  assign n4631 = ~n4625 & n4630;
  assign n4632_1 = Ng3087 & n4551_1;
  assign n4633 = Ng3210 & n4572;
  assign n4634 = Ng3091 & n4568;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = Ng3096 & n4565_1;
  assign n4637_1 = Ng3085 & n4583_1;
  assign n4638 = ~n4636 & ~n4637_1;
  assign n4639 = n4635 & n4638;
  assign n4640 = ~n4632_1 & n4639;
  assign n4641_1 = n4631 & n4640;
  assign n4642 = ~n4527_1 & n4609;
  assign n4643 = Ng3120 & ~n4642;
  assign n4644 = Ng3093 & n4586;
  assign n4645_1 = ~Ng2984 & ~Ng2985;
  assign n4646 = n4543 & ~n4645_1;
  assign n4647 = ~n4644 & ~n4646;
  assign n4648 = Ng3095 & n4574_1;
  assign n4649_1 = Ng3211 & n4578_1;
  assign n4650 = ~n4648 & ~n4649_1;
  assign n4651 = n4647 & n4650;
  assign n4652 = ~n4643 & n4651;
  assign n4653_1 = ~Pg25442 & n4652;
  assign Pg26104 = ~n4641_1 | ~n4653_1;
  assign n4655 = ~Ng3120 & ~n4645_1;
  assign n4656 = ~n4530 & ~n4541;
  assign n4657_1 = ~n4655 & n4656;
  assign n4658 = ~Ng3147 & ~n4657_1;
  assign n4659 = Ng3147 & n4564;
  assign n4660 = Ng3097 & n4659;
  assign Pg25489 = n4658 | n4660;
  assign n4662 = ~Ng3125 & n4527_1;
  assign n864_1 = ~Pg25442 & ~n4662;
  assign n4664 = ~Ng3123 & n4527_1;
  assign n869_1 = ~Pg25442 & ~n4664;
  assign n4666 = Pg5388 & ~Ng2986;
  assign Pg16496 = ~Ng2987 | n4666;
  assign n275_1 = ~Pg51 & Ng13457;
  assign n280 = ~Pg51 & Ng2817;
  assign n285_1 = Pg51 | Ng2933;
  assign n4671 = ~Ng13457 & Ng2883;
  assign n4672 = Ng13457 & ~Ng2883;
  assign n4673_1 = ~Pg8021 & ~n4672;
  assign n290_1 = n4671 | ~n4673_1;
  assign n4675 = Ng2888 & n4672;
  assign n4676 = ~Ng2896 & ~Ng2900;
  assign n4677_1 = Ng2892 & Ng2903;
  assign n4678 = n4676 & n4677_1;
  assign n4679 = n4675 & n4678;
  assign n4680 = Ng2908 & n4679;
  assign n4681_1 = ~Pg8021 & ~n4680;
  assign n4682 = Ng13457 & Ng2883;
  assign n4683 = ~Ng2888 & ~n4682;
  assign n4684 = Ng2888 & n4682;
  assign n4685_1 = ~n4683 & ~n4684;
  assign n295_1 = n4681_1 & n4685_1;
  assign n4687 = ~Ng2896 & ~n4684;
  assign n4688 = Ng2896 & n4684;
  assign n4689_1 = ~n4687 & ~n4688;
  assign n300_1 = n4681_1 & n4689_1;
  assign n4691 = Ng2892 & n4688;
  assign n4692 = ~Ng2892 & ~n4688;
  assign n4693_1 = ~n4691 & ~n4692;
  assign n305_1 = n4681_1 & n4693_1;
  assign n4695 = Ng2903 & n4691;
  assign n4696 = ~Ng2903 & ~n4691;
  assign n4697_1 = n4681_1 & ~n4696;
  assign n310_1 = ~n4695 & n4697_1;
  assign n4699 = Ng2900 & n4695;
  assign n4700 = ~Ng2900 & ~n4695;
  assign n4701_1 = n4681_1 & ~n4700;
  assign n315 = ~n4699 & n4701_1;
  assign n4703 = ~Ng2908 & ~n4699;
  assign n4704 = Ng2908 & n4699;
  assign n4705_1 = ~n4703 & ~n4704;
  assign n320_1 = n4681_1 & n4705_1;
  assign n4707 = Ng2912 & n4680;
  assign n4708 = ~Ng2912 & ~n4680;
  assign n4709_1 = ~n4707 & ~n4708;
  assign n4710 = ~Ng2917 & ~Ng2924;
  assign n4711 = Ng2920 & n4707;
  assign n4712 = n4710 & n4711;
  assign n4713_1 = ~Pg8021 & ~n4712;
  assign n325_1 = n4709_1 | ~n4713_1;
  assign n4715 = ~Ng2917 & ~n4707;
  assign n4716 = Ng2917 & n4707;
  assign n4717_1 = ~n4715 & ~n4716;
  assign n330_1 = n4713_1 & n4717_1;
  assign n4719 = Ng2924 & n4716;
  assign n4720 = ~Ng2924 & ~n4716;
  assign n4721_1 = ~n4719 & ~n4720;
  assign n335_1 = n4713_1 & n4721_1;
  assign n4723 = ~Ng2920 & ~n4719;
  assign n4724 = Ng2920 & n4719;
  assign n4725_1 = ~n4723 & ~n4724;
  assign n340_1 = n4713_1 & n4725_1;
  assign n4727 = ~Ng2956 & Ng2959;
  assign n4728 = Ng2956 & ~Ng2959;
  assign n4729_1 = ~n4727 & ~n4728;
  assign n4730 = Ng2935 & Ng2938;
  assign n4731 = ~Ng2935 & ~Ng2938;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733_1 = n4729_1 & n4732;
  assign n4734 = ~n4729_1 & ~n4732;
  assign n4735 = ~n4733_1 & ~n4734;
  assign n4736 = ~Ng2947 & Ng2953;
  assign n4737 = Ng2947 & ~Ng2953;
  assign n4738_1 = ~n4736 & ~n4737;
  assign n4739 = Ng2941 & Ng2944;
  assign n4740 = ~Ng2941 & ~Ng2944;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = ~n4738_1 & n4741;
  assign n4743_1 = n4738_1 & ~n4741;
  assign n4744 = ~n4742 & ~n4743_1;
  assign n4745 = n4735 & n4744;
  assign n4746 = ~n4735 & ~n4744;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748_1 = Ng2934 & ~n4747;
  assign n4749 = ~Ng2934 & n4747;
  assign n345_1 = ~n4748_1 & ~n4749;
  assign n4751 = ~Ng2981 & Ng2874;
  assign n4752 = Ng2981 & ~Ng2874;
  assign n4753_1 = ~n4751 & ~n4752;
  assign n4754 = Ng2963 & Ng2966;
  assign n4755 = ~Ng2963 & ~Ng2966;
  assign n4756 = ~n4754 & ~n4755;
  assign n4757_1 = n4753_1 & n4756;
  assign n4758 = ~n4753_1 & ~n4756;
  assign n4759 = ~n4757_1 & ~n4758;
  assign n4760 = ~Ng2975 & Ng2978;
  assign n4761_1 = Ng2975 & ~Ng2978;
  assign n4762 = ~n4760 & ~n4761_1;
  assign n4763 = Ng2969 & Ng2972;
  assign n4764 = ~Ng2969 & ~Ng2972;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766_1 = ~n4762 & n4765;
  assign n4767 = n4762 & ~n4765;
  assign n4768 = ~n4766_1 & ~n4767;
  assign n4769 = n4759 & n4768;
  assign n4770_1 = ~n4759 & ~n4768;
  assign n4771 = ~n4769 & ~n4770_1;
  assign n4772 = Ng2962 & ~n4771;
  assign n4773 = ~Ng2962 & n4771;
  assign n350_1 = ~n4772 & ~n4773;
  assign n4775_1 = Pg8021 & ~Ng2929;
  assign n359_1 = ~Ng2879 | n4775_1;
  assign n4777 = Ng2879 & Ng2959;
  assign n4778 = ~Ng2879 & Ng1506;
  assign n436 = n4777 | n4778;
  assign n4780 = Ng2879 & Ng2956;
  assign n4781 = ~Ng2879 & Ng1501;
  assign n441_1 = n4780 | n4781;
  assign n4783 = Ng2879 & Ng2953;
  assign n4784_1 = ~Ng2879 & Ng1496;
  assign n446_1 = n4783 | n4784_1;
  assign n4786 = Ng2879 & Ng2947;
  assign n4787 = ~Ng2879 & Ng1491;
  assign n451 = n4786 | n4787;
  assign n4789 = Ng2879 & Ng2944;
  assign n4790 = ~Ng2879 & Ng1486;
  assign n456 = n4789 | n4790;
  assign n4792 = Ng2879 & Ng2941;
  assign n4793_1 = ~Ng2879 & Ng1481;
  assign n461_1 = n4792 | n4793_1;
  assign n4795 = Ng2879 & Ng2938;
  assign n4796 = ~Ng2879 & Ng1476;
  assign n466_1 = n4795 | n4796;
  assign n4798 = Ng2879 & Ng2935;
  assign n4799 = ~Ng2879 & Ng1471;
  assign n471_1 = n4798 | n4799;
  assign n4801 = ~Ng2879 & ~Ng13439;
  assign n4802_1 = ~Pg3231 & Ng3139;
  assign n4803 = ~n4747 & ~n4802_1;
  assign n4804 = n4747 & n4802_1;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806_1 = Ng2879 & ~n4805;
  assign n476_1 = ~n4801 & ~n4806_1;
  assign n4808 = Ng2879 & Pg8251;
  assign n4809 = ~Ng2879 & Ng2874;
  assign n481 = n4808 | n4809;
  assign n4811_1 = Ng2879 & Pg4090;
  assign n4812 = ~Ng2879 & Ng2981;
  assign n489 = n4811_1 | n4812;
  assign n4814 = Ng2879 & Pg4323;
  assign n4815_1 = ~Ng2879 & Ng2978;
  assign n497_1 = n4814 | n4815_1;
  assign n4817 = Ng2879 & Pg4590;
  assign n4818 = ~Ng2879 & Ng2975;
  assign n505_1 = n4817 | n4818;
  assign n4820_1 = Ng2879 & Pg6225;
  assign n4821 = ~Ng2879 & Ng2972;
  assign n513_1 = n4820_1 | n4821;
  assign n4823 = Ng2879 & Pg6442;
  assign n4824 = ~Ng2879 & Ng2969;
  assign n521_1 = n4823 | n4824;
  assign n4826 = Ng2879 & Pg6895;
  assign n4827 = ~Ng2879 & Ng2966;
  assign n529_1 = n4826 | n4827;
  assign n4829 = Ng2879 & Pg7334;
  assign n4830_1 = ~Ng2879 & Ng2963;
  assign n537_1 = n4829 | n4830_1;
  assign n4832 = Ng2879 & Pg7519;
  assign n4833 = ~n4771 & n4802_1;
  assign n4834 = n4771 & ~n4802_1;
  assign n4835_1 = ~n4833 & ~n4834;
  assign n4836 = ~Ng2879 & ~n4835_1;
  assign n545_1 = n4832 | n4836;
  assign n4838 = Ng2879 & Pg8249;
  assign n4839_1 = ~Ng2879 & Ng2959;
  assign n553_1 = n4838 | n4839_1;
  assign n4841 = Ng2879 & Pg4088;
  assign n4842 = ~Ng2879 & Ng2956;
  assign n561_1 = n4841 | n4842;
  assign n4844 = Ng2879 & Pg4321;
  assign n4845 = ~Ng2879 & Ng2953;
  assign n569_1 = n4844 | n4845;
  assign n4847_1 = Ng2879 & Pg8023;
  assign n4848 = ~Ng2879 & Ng2947;
  assign n577_1 = n4847_1 | n4848;
  assign n4850 = Ng2879 & Pg8175;
  assign n4851 = ~Ng2879 & Ng2944;
  assign n585_1 = n4850 | n4851;
  assign n4853 = Ng2879 & Pg3993;
  assign n4854 = ~Ng2879 & Ng2941;
  assign n593 = n4853 | n4854;
  assign n4856 = Ng2879 & Pg4200;
  assign n4857_1 = ~Ng2879 & Ng2938;
  assign n601_1 = n4856 | n4857_1;
  assign n4859 = Ng2879 & Pg4450;
  assign n4860 = ~Ng2879 & Ng2935;
  assign n609_1 = n4859 | n4860;
  assign n4862_1 = Ng2879 & ~Pg8096;
  assign n4863 = ~Ng2879 & ~n4805;
  assign n617_1 = ~n4862_1 & ~n4863;
  assign n4865 = Ng2879 & Ng2874;
  assign n4866 = ~Ng2879 & Ng2200;
  assign n625_1 = n4865 | n4866;
  assign n4868 = Ng2879 & Ng2981;
  assign n4869 = ~Ng2879 & Ng2195;
  assign n630 = n4868 | n4869;
  assign n4871 = Ng2879 & Ng2978;
  assign n4872 = ~Ng2879 & Ng2190;
  assign n635_1 = n4871 | n4872;
  assign n4874 = Ng2879 & Ng2975;
  assign n4875 = ~Ng2879 & Ng2185;
  assign n640_1 = n4874 | n4875;
  assign n4877_1 = Ng2879 & Ng2972;
  assign n4878 = ~Ng2879 & Ng2180;
  assign n645_1 = n4877_1 | n4878;
  assign n4880 = Ng2879 & Ng2969;
  assign n4881_1 = ~Ng2879 & Ng2175;
  assign n650 = n4880 | n4881_1;
  assign n4883 = Ng2879 & Ng2966;
  assign n4884 = ~Ng2879 & Ng2170;
  assign n655 = n4883 | n4884;
  assign n4886 = Ng2879 & Ng2963;
  assign n4887 = ~Ng2879 & Ng2165;
  assign n660 = n4886 | n4887;
  assign n4889_1 = ~Ng2879 & Ng13455;
  assign n4890 = Ng2879 & ~n4835_1;
  assign n665_1 = n4889_1 | n4890;
  assign n4892 = Ng559 & \[1605] ;
  assign n4893 = Ng3210 & ~\[1605] ;
  assign n670 = n4892 | n4893;
  assign n4895 = Ng559 & \[1603] ;
  assign n4896 = Ng3211 & ~\[1603] ;
  assign n675_1 = n4895 | n4896;
  assign n4898 = Ng559 & Ng1315;
  assign n4899 = Ng3084 & ~Ng1315;
  assign n680 = n4898 | n4899;
  assign n4901 = Ng1245 & \[1605] ;
  assign n4902_1 = Ng3085 & ~\[1605] ;
  assign n685_1 = n4901 | n4902_1;
  assign n4904 = Ng1245 & \[1603] ;
  assign n4905 = Ng3086 & ~\[1603] ;
  assign n690 = n4904 | n4905;
  assign n4907 = Ng1245 & Ng1315;
  assign n4908 = Ng3087 & ~Ng1315;
  assign n695_1 = n4907 | n4908;
  assign n4910 = \[1605]  & Ng1939;
  assign n4911_1 = Ng3091 & ~\[1605] ;
  assign n700_1 = n4910 | n4911_1;
  assign n4913 = \[1603]  & Ng1939;
  assign n4914 = Ng3092 & ~\[1603] ;
  assign n705_1 = n4913 | n4914;
  assign n4916_1 = Ng1315 & Ng1939;
  assign n4917 = Ng3093 & ~Ng1315;
  assign n710_1 = n4916_1 | n4917;
  assign n4919 = \[1605]  & Ng2633;
  assign n4920_1 = Ng3094 & ~\[1605] ;
  assign n715_1 = n4919 | n4920_1;
  assign n4922 = \[1603]  & Ng2633;
  assign n4923 = Ng3095 & ~\[1603] ;
  assign n720 = n4922 | n4923;
  assign n4925_1 = Ng1315 & Ng2633;
  assign n4926 = Ng3096 & ~Ng1315;
  assign n725 = n4925_1 | n4926;
  assign n4928 = Ng544 & Ng8284;
  assign n4929_1 = \[1605]  & n4928;
  assign n4930 = Ng3097 & ~\[1605] ;
  assign n730_1 = n4929_1 | n4930;
  assign n4932 = Ng3098 & ~\[1603] ;
  assign n4933 = Ng548 & ~Ng8284;
  assign n4934_1 = ~\[1605]  & n4933;
  assign n1898_1 = n4928 | n4934_1;
  assign n4936 = \[1603]  & n1898_1;
  assign n735_1 = n4932 | n4936;
  assign n4938 = Ng3099 & ~Ng1315;
  assign n4939_1 = Ng1315 & n1898_1;
  assign n740_1 = n4938 | n4939_1;
  assign n4941 = Ng1234 & ~\[1605] ;
  assign n4942 = ~Ng8293 & ~n4941;
  assign n4943 = ~n4929_1 & n4942;
  assign n4944_1 = ~Ng1230 & Ng8293;
  assign n3404_1 = ~n4943 & ~n4944_1;
  assign n4946 = \[1605]  & ~n3404_1;
  assign n4947 = ~Ng3100 & ~\[1605] ;
  assign n745_1 = ~n4946 & ~n4947;
  assign n4949_1 = ~Ng3101 & ~\[1603] ;
  assign n4950 = \[1603]  & ~n3404_1;
  assign n750_1 = ~n4949_1 & ~n4950;
  assign n4952 = ~Ng3102 & ~Ng1315;
  assign n4953 = Ng1315 & ~n3404_1;
  assign n755_1 = ~n4952 & ~n4953;
  assign n4955 = ~\[1605]  & ~Ng1928;
  assign n4956 = ~Ng8302 & ~n4955;
  assign n4957 = ~n4946 & n4956;
  assign n4958 = Ng1924 & Ng8302;
  assign n4911 = n4957 | n4958;
  assign n4960 = \[1605]  & n4911;
  assign n4961 = Ng3103 & ~\[1605] ;
  assign n760_1 = n4960 | n4961;
  assign n4963 = Ng3104 & ~\[1603] ;
  assign n4964_1 = \[1603]  & n4911;
  assign n765_1 = n4963 | n4964_1;
  assign n4966 = Ng3105 & ~Ng1315;
  assign n4967 = Ng1315 & n4911;
  assign n770_1 = n4966 | n4967;
  assign n4969_1 = ~Ng3106 & ~\[1605] ;
  assign n4970 = ~Ng2618 & Ng8311;
  assign n4971 = ~\[1605]  & Ng2622;
  assign n4972 = ~Ng8311 & ~n4971;
  assign n4973 = ~n4960 & n4972;
  assign n6418 = ~n4970 & ~n4973;
  assign n4975 = \[1605]  & ~n6418;
  assign n775_1 = ~n4969_1 & ~n4975;
  assign n4977 = ~Ng3107 & ~\[1603] ;
  assign n4978 = \[1603]  & ~n6418;
  assign n780_1 = ~n4977 & ~n4978;
  assign n4980 = ~Ng3108 & ~Ng1315;
  assign n4981 = Ng1315 & ~n6418;
  assign n785_1 = ~n4980 & ~n4981;
  assign n4983 = ~Ng3155 & ~\[1605] ;
  assign n4984_1 = ~Ng8284 & \[1605] ;
  assign n790_1 = ~n4983 & ~n4984_1;
  assign n4986 = Ng8284 & \[1603] ;
  assign n4987 = Ng3158 & ~\[1603] ;
  assign n795_1 = n4986 | n4987;
  assign n4989_1 = Ng8284 & Ng1315;
  assign n4990 = Ng3161 & ~Ng1315;
  assign n800_1 = n4989_1 | n4990;
  assign n4992 = Ng8293 & \[1605] ;
  assign n4993 = Ng3164 & ~\[1605] ;
  assign n805_1 = n4992 | n4993;
  assign n4995 = Ng8293 & \[1603] ;
  assign n4996 = Ng3167 & ~\[1603] ;
  assign n810_1 = n4995 | n4996;
  assign n4998 = Ng8293 & Ng1315;
  assign n4999_1 = Ng3170 & ~Ng1315;
  assign n815_1 = n4998 | n4999_1;
  assign n5001 = \[1605]  & Ng8302;
  assign n5002 = Ng3173 & ~\[1605] ;
  assign n820 = n5001 | n5002;
  assign n5004_1 = \[1603]  & Ng8302;
  assign n5005 = Ng3176 & ~\[1603] ;
  assign n825_1 = n5004_1 | n5005;
  assign n5007 = Ng1315 & Ng8302;
  assign n5008 = Ng3179 & ~Ng1315;
  assign n830_1 = n5007 | n5008;
  assign n5010 = \[1605]  & Ng8311;
  assign n5011 = Ng3182 & ~\[1605] ;
  assign n835_1 = n5010 | n5011;
  assign n5013 = \[1603]  & Ng8311;
  assign n5014_1 = Ng3185 & ~\[1603] ;
  assign n840_1 = n5013 | n5014_1;
  assign n5016 = Ng1315 & Ng8311;
  assign n5017 = Ng3088 & ~Ng1315;
  assign n845_1 = n5016 | n5017;
  assign n5019_1 = \[1612]  & Ng2257;
  assign n5020 = Ng130 & ~n5019_1;
  assign n5021 = ~Ng97 & n5019_1;
  assign n899_1 = n5020 | n5021;
  assign n5023 = \[1594]  & Ng2257;
  assign n5024_1 = Ng131 & ~n5023;
  assign n5025 = ~Ng97 & n5023;
  assign n904_1 = n5024_1 | n5025;
  assign n5027 = Ng853 & Ng2257;
  assign n5028 = Ng129 & ~n5027;
  assign n5029_1 = ~Ng97 & n5027;
  assign n909_1 = n5028 | n5029_1;
  assign n5031 = Ng133 & ~n5019_1;
  assign n5032 = ~Ng101 & n5019_1;
  assign n914_1 = n5031 | n5032;
  assign n5034_1 = Ng134 & ~n5023;
  assign n5035 = ~Ng101 & n5023;
  assign n919_1 = n5034_1 | n5035;
  assign n5037 = Ng132 & ~n5027;
  assign n5038 = ~Ng101 & n5027;
  assign n924_1 = n5037 | n5038;
  assign n5040 = Ng142 & ~n5019_1;
  assign n5041 = ~Ng105 & n5019_1;
  assign n929_1 = n5040 | n5041;
  assign n5043 = Ng143 & ~n5023;
  assign n5044_1 = ~Ng105 & n5023;
  assign n934 = n5043 | n5044_1;
  assign n5046 = Ng141 & ~n5027;
  assign n5047 = ~Ng105 & n5027;
  assign n939_1 = n5046 | n5047;
  assign n5049_1 = Ng145 & ~n5019_1;
  assign n5050 = ~Ng109 & n5019_1;
  assign n944_1 = n5049_1 | n5050;
  assign n5052 = Ng146 & ~n5023;
  assign n5053 = ~Ng109 & n5023;
  assign n949_1 = n5052 | n5053;
  assign n5055 = Ng144 & ~n5027;
  assign n5056 = ~Ng109 & n5027;
  assign n954_1 = n5055 | n5056;
  assign n5058 = Ng148 & ~n5019_1;
  assign n5059_1 = ~Ng113 & n5019_1;
  assign n959_1 = n5058 | n5059_1;
  assign n5061 = Ng149 & ~n5023;
  assign n5062 = ~Ng113 & n5023;
  assign n964_1 = n5061 | n5062;
  assign n5064_1 = Ng147 & ~n5027;
  assign n5065 = ~Ng113 & n5027;
  assign n969_1 = n5064_1 | n5065;
  assign n5067 = Ng151 & ~n5019_1;
  assign n5068_1 = ~Ng117 & n5019_1;
  assign n974_1 = n5067 | n5068_1;
  assign n5070 = Ng152 & ~n5023;
  assign n5071 = ~Ng117 & n5023;
  assign n979_1 = n5070 | n5071;
  assign n5073_1 = Ng150 & ~n5027;
  assign n5074 = ~Ng117 & n5027;
  assign n984_1 = n5073_1 | n5074;
  assign n5076 = Ng154 & ~n5019_1;
  assign n5077 = ~Ng121 & n5019_1;
  assign n989_1 = n5076 | n5077;
  assign n5079 = Ng155 & ~n5023;
  assign n5080 = ~Ng121 & n5023;
  assign n994_1 = n5079 | n5080;
  assign n5082 = Ng153 & ~n5027;
  assign n5083 = ~Ng121 & n5027;
  assign n999_1 = n5082 | n5083;
  assign n5085 = Ng157 & ~n5019_1;
  assign n5086_1 = ~Ng125 & n5019_1;
  assign n1004_1 = n5085 | n5086_1;
  assign n5088 = Ng158 & ~n5023;
  assign n5089 = ~Ng125 & n5023;
  assign n1009_1 = n5088 | n5089;
  assign n5091_1 = Ng156 & ~n5027;
  assign n5092 = ~Ng125 & n5027;
  assign n1014 = n5091_1 | n5092;
  assign n5094 = ~Ng160 & ~n5019_1;
  assign n5095 = ~Ng174 & Ng853;
  assign n5096_1 = ~Ng175 & \[1612] ;
  assign n5097 = ~Ng176 & \[1594] ;
  assign n5098 = ~n5096_1 & ~n5097;
  assign n5099 = ~n5095 & n5098;
  assign n5100 = n5019_1 & ~n5099;
  assign n1019_1 = ~n5094 & ~n5100;
  assign n5102 = n5023 & n5099;
  assign n5103 = Ng161 & ~n5023;
  assign n1024_1 = n5102 | n5103;
  assign n5105 = ~Ng159 & ~n5027;
  assign n5106_1 = n5027 & ~n5099;
  assign n1029 = ~n5105 & ~n5106_1;
  assign n5108 = ~Ng163 & ~n5019_1;
  assign n5109 = ~Ng171 & Ng853;
  assign n5110 = ~Ng173 & \[1594] ;
  assign n5111_1 = ~Ng172 & \[1612] ;
  assign n5112 = ~n5110 & ~n5111_1;
  assign n5113 = ~n5109 & n5112;
  assign n5114 = n5019_1 & ~n5113;
  assign n1034_1 = ~n5108 & ~n5114;
  assign n5116_1 = n5023 & n5113;
  assign n5117 = Ng164 & ~n5023;
  assign n1039_1 = n5116_1 | n5117;
  assign n5119 = ~Ng162 & ~n5027;
  assign n5120 = n5027 & ~n5113;
  assign n1044 = ~n5119 & ~n5120;
  assign n5122 = ~Ng2892 & ~Ng2908;
  assign n5123 = n4676 & n5122;
  assign n5124 = ~Ng2903 & n5123;
  assign n5125 = ~Ng2912 & ~Ng2917;
  assign n5126_1 = Ng2924 & ~Ng2920;
  assign n5127 = n5125 & n5126_1;
  assign n5128 = Ng2883 & ~Ng2888;
  assign n5129 = n5127 & n5128;
  assign n5816 = n5124 & n5129;
  assign n5131_1 = \[1612]  & n5816;
  assign n5132 = Ng125 & Ng113;
  assign n5133 = ~Ng117 & n5132;
  assign n5134 = ~Ng121 & n5133;
  assign n5135 = n5131_1 & n5134;
  assign n5136_1 = Ng169 & ~n5131_1;
  assign n1049 = n5135 | n5136_1;
  assign n5138 = \[1594]  & n5816;
  assign n5139 = n5134 & n5138;
  assign n5140 = Ng170 & ~n5138;
  assign n1054_1 = n5139 | n5140;
  assign n5142 = Ng853 & n5816;
  assign n5143 = n5134 & n5142;
  assign n5144 = Ng168 & ~n5142;
  assign n1059_1 = n5143 | n5144;
  assign n5146_1 = Ng172 & ~n5131_1;
  assign n5147 = ~Ng101 & n5131_1;
  assign n1064_1 = n5146_1 | n5147;
  assign n5149 = Ng173 & ~n5138;
  assign n5150 = ~Ng101 & n5138;
  assign n1069 = n5149 | n5150;
  assign n5152 = Ng171 & ~n5142;
  assign n5153 = ~Ng101 & n5142;
  assign n1074_1 = n5152 | n5153;
  assign n5155 = Ng175 & ~n5131_1;
  assign n5156_1 = ~Ng97 & n5131_1;
  assign n1079 = n5155 | n5156_1;
  assign n5158 = Ng176 & ~n5138;
  assign n5159 = ~Ng97 & n5138;
  assign n1084_1 = n5158 | n5159;
  assign n5161_1 = Ng174 & ~n5142;
  assign n5162 = ~Ng97 & n5142;
  assign n1089_1 = n5161_1 | n5162;
  assign n5164 = Ng178 & ~n5131_1;
  assign n5165 = Ng101 & Ng97;
  assign n5166_1 = Ng109 & Ng105;
  assign n5167 = n5165 & n5166_1;
  assign n5168 = Ng121 & Ng117;
  assign n5169 = n5132 & n5168;
  assign n5170 = n5167 & n5169;
  assign n5171_1 = n5131_1 & ~n5170;
  assign n1094_1 = n5164 | n5171_1;
  assign n5173 = Ng179 & ~n5138;
  assign n5174 = n5138 & ~n5170;
  assign n1099_1 = n5173 | n5174;
  assign n5176_1 = Ng177 & ~n5142;
  assign n5177 = n5142 & ~n5170;
  assign n1104_1 = n5176_1 | n5177;
  assign n5179 = ~Ng186 & ~\[1612] ;
  assign n5180 = Ng192 & Ng853;
  assign n5181_1 = Ng186 & \[1612] ;
  assign n5182 = Ng189 & \[1594] ;
  assign n5183 = ~n5181_1 & ~n5182;
  assign n5184 = ~n5180 & n5183;
  assign n5185 = ~Ng320 & Ng853;
  assign n5186_1 = ~Ng318 & \[1612] ;
  assign n5187 = ~Ng319 & \[1594] ;
  assign n5188 = ~n5186_1 & ~n5187;
  assign n5189 = ~n5185 & n5188;
  assign n5190 = ~Ng314 & Ng853;
  assign n5191_1 = ~Ng312 & \[1612] ;
  assign n5192 = ~Ng313 & \[1594] ;
  assign n5193 = ~n5191_1 & ~n5192;
  assign n5194 = ~n5190 & n5193;
  assign n5195 = n5189 & n5194;
  assign n5196_1 = n5184 & n5195;
  assign n5197 = Ng264 & Ng853;
  assign n5198 = Ng258 & \[1612] ;
  assign n5199 = Ng261 & \[1594] ;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201_1 = ~n5197 & n5200;
  assign n5202 = Ng216 & \[1594] ;
  assign n5203 = Ng219 & Ng853;
  assign n5204 = Ng213 & \[1612] ;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206_1 = ~n5202 & n5205;
  assign n5207 = n5201_1 & n5206_1;
  assign n5208 = Ng210 & Ng853;
  assign n5209 = Ng204 & \[1612] ;
  assign n5210 = Ng207 & \[1594] ;
  assign n5211_1 = ~n5209 & ~n5210;
  assign n5212 = ~n5208 & n5211_1;
  assign n5213 = Ng255 & Ng853;
  assign n5214 = Ng249 & \[1612] ;
  assign n5215 = Ng252 & \[1594] ;
  assign n5216_1 = ~n5214 & ~n5215;
  assign n5217 = ~n5213 & n5216_1;
  assign n5218 = n5212 & n5217;
  assign n5219 = n5207 & n5218;
  assign n5220 = n5196_1 & n5219;
  assign n5221_1 = ~Ng317 & Ng853;
  assign n5222 = ~Ng315 & \[1612] ;
  assign n5223 = ~Ng316 & \[1594] ;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5221_1 & n5224;
  assign n5226_1 = Ng201 & Ng853;
  assign n5227 = Ng195 & \[1612] ;
  assign n5228 = Ng198 & \[1594] ;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = ~n5226_1 & n5229;
  assign n5231_1 = n5225 & n5230;
  assign n5232 = Ng222 & \[1612] ;
  assign n5233 = Ng225 & \[1594] ;
  assign n5234 = Ng228 & Ng853;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236_1 = ~n5232 & n5235;
  assign n5237 = Ng273 & Ng853;
  assign n5238 = Ng267 & \[1612] ;
  assign n5239 = Ng270 & \[1594] ;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241_1 = ~n5237 & n5240;
  assign n5242 = n5236_1 & n5241_1;
  assign n5243 = n5231_1 & n5242;
  assign n5244 = Ng237 & Ng853;
  assign n5245 = Ng231 & \[1612] ;
  assign n5246_1 = Ng234 & \[1594] ;
  assign n5247 = ~n5245 & ~n5246_1;
  assign n5248 = ~n5244 & n5247;
  assign n5249 = Ng246 & Ng853;
  assign n5250 = Ng240 & \[1612] ;
  assign n5251_1 = Ng243 & \[1594] ;
  assign n5252 = ~n5250 & ~n5251_1;
  assign n5253 = ~n5249 & n5252;
  assign n5254 = n5248 & n5253;
  assign n5255 = n5243 & n5254;
  assign n5256_1 = n5220 & n5255;
  assign n5257 = ~n5194 & n5225;
  assign n5258 = ~n5189 & n5257;
  assign n5259 = n5189 & ~n5194;
  assign n5260 = ~Ng168 & Ng853;
  assign n5261_1 = ~Ng170 & \[1594] ;
  assign n5262 = ~Ng169 & \[1612] ;
  assign n5263 = ~n5261_1 & ~n5262;
  assign n5264 = ~n5260 & n5263;
  assign n5265 = Ng2257 & ~n5264;
  assign n5266_1 = ~Ng101 & ~n5248;
  assign n5267 = Ng101 & n5248;
  assign n5268 = ~n5266_1 & ~n5267;
  assign n5269 = ~Ng109 & ~n5253;
  assign n5270 = Ng109 & n5253;
  assign n5271_1 = ~n5269 & ~n5270;
  assign n5272 = n5268 & n5271_1;
  assign n5273 = ~Ng125 & ~n5201_1;
  assign n5274 = Ng125 & n5201_1;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276_1 = ~Ng117 & ~n5217;
  assign n5277 = Ng117 & n5217;
  assign n5278 = ~n5276_1 & ~n5277;
  assign n5279 = n5275 & n5278;
  assign n5280 = ~n5113 & ~n5241_1;
  assign n5281_1 = n5113 & n5241_1;
  assign n5282 = ~n5280 & ~n5281_1;
  assign n5283 = ~n5279 & n5282;
  assign n5284 = ~n5272 & n5283;
  assign n5285 = n5275 & ~n5282;
  assign n5286_1 = ~n5268 & ~n5285;
  assign n5287 = n5271_1 & ~n5282;
  assign n5288 = ~n5278 & ~n5287;
  assign n5289 = ~n5286_1 & ~n5288;
  assign n5290 = n5271_1 & n5278;
  assign n5291_1 = n5268 & n5275;
  assign n5292 = ~n5290 & ~n5291_1;
  assign n5293 = ~n5289 & n5292;
  assign n5294 = ~n5284 & ~n5293;
  assign n5295 = n5265 & ~n5294;
  assign n5296_1 = ~Ng97 & ~n5184;
  assign n5297 = Ng97 & n5184;
  assign n5298 = ~n5296_1 & ~n5297;
  assign n5299 = ~Ng105 & ~n5230;
  assign n5300 = Ng105 & n5230;
  assign n5301_1 = ~n5299 & ~n5300;
  assign n5302 = ~n5298 & ~n5301_1;
  assign n5303 = ~Ng113 & ~n5212;
  assign n5304 = Ng113 & n5212;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306_1 = ~n5302 & n5305;
  assign n5307 = n5302 & ~n5305;
  assign n5308 = n5099 & ~n5236_1;
  assign n5309 = ~n5099 & n5236_1;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311_1 = ~n5298 & ~n5310;
  assign n5312 = ~Ng121 & ~n5206_1;
  assign n5313 = Ng121 & n5206_1;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = ~n5311_1 & n5314;
  assign n5316_1 = ~n5307 & n5315;
  assign n5317 = n5298 & n5301_1;
  assign n5318 = n5310 & n5317;
  assign n5319 = ~n5316_1 & ~n5318;
  assign n5320 = ~n5306_1 & n5319;
  assign n5321_1 = n5305 & n5314;
  assign n5322 = ~n5310 & ~n5321_1;
  assign n5323 = ~n5317 & n5322;
  assign n5324 = ~n5320 & ~n5323;
  assign n5325 = n5265 & ~n5324;
  assign n5326_1 = ~n5295 & ~n5325;
  assign n5327 = n5259 & n5326_1;
  assign n5328 = ~n5258 & ~n5327;
  assign n5329 = ~Ng147 & Ng853;
  assign n5330 = ~Ng149 & \[1594] ;
  assign n5331_1 = ~Ng148 & \[1612] ;
  assign n5332 = ~n5330 & ~n5331_1;
  assign n5333 = ~n5329 & n5332;
  assign n5334 = ~Ng113 & ~n5333;
  assign n5335 = ~Ng129 & Ng853;
  assign n5336_1 = ~Ng130 & \[1612] ;
  assign n5337 = ~Ng131 & \[1594] ;
  assign n5338 = ~n5336_1 & ~n5337;
  assign n5339 = ~n5335 & n5338;
  assign n5340 = Ng97 & n5339;
  assign n5341_1 = ~n5334 & ~n5340;
  assign n5342 = ~Ng156 & Ng853;
  assign n5343 = ~Ng157 & \[1612] ;
  assign n5344 = ~Ng158 & \[1594] ;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346_1 = ~n5342 & n5345;
  assign n5347 = Ng125 & n5346_1;
  assign n5348 = ~Ng125 & ~n5346_1;
  assign n5349 = ~n5347 & ~n5348;
  assign n5350 = n5341_1 & n5349;
  assign n5351_1 = ~Ng150 & Ng853;
  assign n5352 = ~Ng152 & \[1594] ;
  assign n5353 = ~Ng151 & \[1612] ;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~n5351_1 & n5354;
  assign n5356_1 = Ng117 & n5355;
  assign n5357 = ~Ng97 & ~n5339;
  assign n5358 = ~n5356_1 & ~n5357;
  assign n5359 = n5265 & n5358;
  assign n5360 = n5350 & n5359;
  assign n5361_1 = ~Ng153 & Ng853;
  assign n5362 = ~Ng154 & \[1612] ;
  assign n5363 = ~Ng155 & \[1594] ;
  assign n5364 = ~n5362 & ~n5363;
  assign n5365 = ~n5361_1 & n5364;
  assign n5366_1 = ~Ng121 & ~n5365;
  assign n5367 = ~Ng132 & Ng853;
  assign n5368 = ~Ng133 & \[1612] ;
  assign n5369 = ~Ng134 & \[1594] ;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371_1 = ~n5367 & n5370;
  assign n5372 = Ng101 & n5371_1;
  assign n5373 = ~Ng141 & Ng853;
  assign n5374 = ~Ng143 & \[1594] ;
  assign n5375 = ~Ng142 & \[1612] ;
  assign n5376_1 = ~n5374 & ~n5375;
  assign n5377 = ~n5373 & n5376_1;
  assign n5378 = ~Ng105 & ~n5377;
  assign n5379 = ~n5372 & ~n5378;
  assign n5380 = ~n5366_1 & n5379;
  assign n5381_1 = n5360 & n5380;
  assign n5382 = ~Ng101 & ~n5371_1;
  assign n5383 = ~Ng159 & Ng853;
  assign n5384 = ~Ng160 & \[1612] ;
  assign n5385 = ~Ng161 & \[1594] ;
  assign n5386_1 = ~n5384 & ~n5385;
  assign n5387 = ~n5383 & n5386_1;
  assign n5388 = n5099 & n5387;
  assign n5389 = ~n5099 & ~n5387;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391_1 = ~n5382 & ~n5390;
  assign n5392 = ~Ng144 & Ng853;
  assign n5393 = ~Ng146 & \[1594] ;
  assign n5394 = ~Ng145 & \[1612] ;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396_1 = ~n5392 & n5395;
  assign n5397 = ~Ng109 & n5396_1;
  assign n5398 = Ng109 & ~n5396_1;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = n5391_1 & ~n5399;
  assign n5401_1 = ~Ng162 & Ng853;
  assign n5402 = ~Ng163 & \[1612] ;
  assign n5403 = ~Ng164 & \[1594] ;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = ~n5401_1 & n5404;
  assign n5406_1 = n5113 & ~n5405;
  assign n5407 = Ng113 & n5333;
  assign n5408 = ~n5406_1 & ~n5407;
  assign n5409 = Ng105 & n5377;
  assign n5410 = n5408 & ~n5409;
  assign n5411_1 = Ng121 & n5365;
  assign n5412 = ~Ng117 & ~n5355;
  assign n5413 = ~n5113 & n5405;
  assign n5414 = ~n5412 & ~n5413;
  assign n5415 = ~n5411_1 & n5414;
  assign n5416_1 = n5410 & n5415;
  assign n5417 = n5400 & n5416_1;
  assign n5418 = n5381_1 & n5417;
  assign n5419 = ~Ng323 & \[1594] ;
  assign n5420 = ~Ng321 & Ng853;
  assign n5421_1 = ~Ng322 & \[1612] ;
  assign n5422 = ~n5420 & ~n5421_1;
  assign n5423 = ~n5419 & n5422;
  assign n5424 = n5418 & ~n5423;
  assign n5425 = n5225 & n5424;
  assign n5426_1 = ~n5328 & n5425;
  assign n5427 = ~Ng402 & Ng853;
  assign n5428 = ~Ng403 & \[1612] ;
  assign n5429 = ~Ng404 & \[1594] ;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431_1 = ~n5427 & n5430;
  assign n5432 = n5418 & ~n5431_1;
  assign n5433 = Ng2257 & n5264;
  assign n5434 = ~n5194 & n5433;
  assign n5435 = ~n5432 & ~n5434;
  assign n5436_1 = ~n5426_1 & n5435;
  assign n5437 = n5195 & ~n5225;
  assign n5438 = ~n5236_1 & n5437;
  assign n5439 = ~n5241_1 & ~n5248;
  assign n5440 = ~n5253 & n5439;
  assign n5441_1 = n5184 & ~n5230;
  assign n5442 = n5440 & n5441_1;
  assign n5443 = n5438 & n5442;
  assign n5444 = n5219 & n5443;
  assign n5445 = n5436_1 & ~n5444;
  assign n5446_1 = ~n5256_1 & n5445;
  assign n5447 = Ng97 & ~n5436_1;
  assign n5448 = ~n5446_1 & ~n5447;
  assign n5449 = ~n5184 & ~n5195;
  assign n5450 = ~n5196_1 & ~n5449;
  assign n5451_1 = n5445 & n5450;
  assign n5452 = ~n5448 & ~n5451_1;
  assign n5453 = \[1612]  & ~n5452;
  assign n1109_1 = ~n5179 & ~n5453;
  assign n5455 = ~Ng189 & ~\[1594] ;
  assign n5456_1 = \[1594]  & ~n5452;
  assign n1114 = ~n5455 & ~n5456_1;
  assign n5458 = ~Ng192 & ~Ng853;
  assign n5459 = Ng853 & ~n5452;
  assign n1119_1 = ~n5458 & ~n5459;
  assign n5461_1 = ~Ng231 & ~\[1612] ;
  assign n5462 = Ng101 & ~n5436_1;
  assign n5463 = ~n5445 & ~n5462;
  assign n5464 = n5184 & n5225;
  assign n5465 = ~n5184 & ~n5225;
  assign n5466_1 = ~n5464 & ~n5465;
  assign n5467 = n5195 & ~n5466_1;
  assign n5468 = ~n5248 & n5467;
  assign n5469 = n5248 & ~n5467;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471_1 = n5446_1 & ~n5470;
  assign n5472 = ~n5463 & ~n5471_1;
  assign n5473 = \[1612]  & ~n5472;
  assign n1124_1 = ~n5461_1 & ~n5473;
  assign n5475 = ~Ng234 & ~\[1594] ;
  assign n5476_1 = \[1594]  & ~n5472;
  assign n1129_1 = ~n5475 & ~n5476_1;
  assign n5478 = ~Ng237 & ~Ng853;
  assign n5479 = Ng853 & ~n5472;
  assign n1134_1 = ~n5478 & ~n5479;
  assign n5481_1 = ~Ng195 & ~\[1612] ;
  assign n5482 = Ng105 & ~n5436_1;
  assign n5483 = ~n5445 & ~n5482;
  assign n5484 = ~n5248 & n5465;
  assign n5485 = n5248 & n5464;
  assign n5486_1 = ~n5484 & ~n5485;
  assign n5487 = n5195 & ~n5486_1;
  assign n5488 = n5230 & n5487;
  assign n5489 = ~n5230 & ~n5487;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491_1 = n5446_1 & n5490;
  assign n5492 = ~n5483 & ~n5491_1;
  assign n5493 = \[1612]  & ~n5492;
  assign n1139_1 = ~n5481_1 & ~n5493;
  assign n5495 = ~Ng198 & ~\[1594] ;
  assign n5496_1 = \[1594]  & ~n5492;
  assign n1144_1 = ~n5495 & ~n5496_1;
  assign n5498 = ~Ng201 & ~Ng853;
  assign n5499 = Ng853 & ~n5492;
  assign n1149_1 = ~n5498 & ~n5499;
  assign n5501_1 = ~Ng240 & ~\[1612] ;
  assign n5502 = Ng109 & ~n5436_1;
  assign n5503 = ~n5445 & ~n5502;
  assign n5504 = ~n5225 & ~n5230;
  assign n5505 = ~n5231_1 & ~n5504;
  assign n5506_1 = n5487 & ~n5505;
  assign n5507 = ~n5253 & n5506_1;
  assign n5508 = n5253 & ~n5506_1;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = n5446_1 & ~n5509;
  assign n5511_1 = ~n5503 & ~n5510;
  assign n5512 = \[1612]  & ~n5511_1;
  assign n1154_1 = ~n5501_1 & ~n5512;
  assign n5514 = ~Ng243 & ~\[1594] ;
  assign n5515 = \[1594]  & ~n5511_1;
  assign n1159_1 = ~n5514 & ~n5515;
  assign n5517 = ~Ng246 & ~Ng853;
  assign n5518 = Ng853 & ~n5511_1;
  assign n1164 = ~n5517 & ~n5518;
  assign n5520 = Ng113 & ~n5436_1;
  assign n5521_1 = ~n5253 & ~n5437;
  assign n5522 = n5253 & n5437;
  assign n5523 = ~n5521_1 & ~n5522;
  assign n5524 = n5506_1 & n5523;
  assign n5525 = ~n5212 & n5524;
  assign n5526_1 = n5212 & ~n5524;
  assign n5527 = ~n5525 & ~n5526_1;
  assign n5528 = n5446_1 & n5527;
  assign n5529 = ~n5520 & ~n5528;
  assign n5530 = \[1612]  & n5529;
  assign n5531_1 = ~Ng204 & ~\[1612] ;
  assign n1169_1 = ~n5530 & ~n5531_1;
  assign n5533 = \[1594]  & n5529;
  assign n5534 = ~Ng207 & ~\[1594] ;
  assign n1174_1 = ~n5533 & ~n5534;
  assign n5536_1 = Ng853 & n5529;
  assign n5537 = ~Ng210 & ~Ng853;
  assign n1179_1 = ~n5536_1 & ~n5537;
  assign n5539 = Ng249 & ~\[1612] ;
  assign n5540 = Ng117 & ~n5436_1;
  assign n5541_1 = ~n5212 & n5437;
  assign n5542 = n5212 & ~n5437;
  assign n5543 = ~n5541_1 & ~n5542;
  assign n5544 = n5524 & ~n5543;
  assign n5545 = n5217 & n5544;
  assign n5546_1 = ~n5217 & ~n5544;
  assign n5547 = ~n5545 & ~n5546_1;
  assign n5548 = n5446_1 & ~n5547;
  assign n5549 = ~n5540 & ~n5548;
  assign n5550 = \[1612]  & ~n5549;
  assign n1184_1 = n5539 | n5550;
  assign n5552 = Ng252 & ~\[1594] ;
  assign n5553 = \[1594]  & ~n5549;
  assign n1189_1 = n5552 | n5553;
  assign n5555 = Ng255 & ~Ng853;
  assign n5556_1 = Ng853 & ~n5549;
  assign n1194 = n5555 | n5556_1;
  assign n5558 = Ng121 & ~n5436_1;
  assign n5559 = n5217 & n5437;
  assign n5560 = n5507 & n5541_1;
  assign n5561_1 = ~n5545 & ~n5560;
  assign n5562 = ~n5559 & ~n5561_1;
  assign n5563 = n5206_1 & n5562;
  assign n5564 = ~n5206_1 & ~n5562;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566_1 = n5446_1 & ~n5565;
  assign n5567 = ~n5558 & ~n5566_1;
  assign n5568 = \[1612]  & n5567;
  assign n5569 = ~Ng213 & ~\[1612] ;
  assign n1199_1 = ~n5568 & ~n5569;
  assign n5571_1 = \[1594]  & n5567;
  assign n5572 = ~Ng216 & ~\[1594] ;
  assign n1204_1 = ~n5571_1 & ~n5572;
  assign n5574 = Ng853 & n5567;
  assign n5575 = ~Ng219 & ~Ng853;
  assign n1209_1 = ~n5574 & ~n5575;
  assign n5577 = Ng125 & ~n5436_1;
  assign n5578 = n5206_1 & ~n5437;
  assign n5579 = ~n5206_1 & n5437;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581_1 = n5562 & ~n5580;
  assign n5582 = ~n5201_1 & n5581_1;
  assign n5583 = n5201_1 & ~n5581_1;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = n5446_1 & n5584;
  assign n5586_1 = ~n5577 & ~n5585;
  assign n5587 = \[1612]  & n5586_1;
  assign n5588 = ~Ng258 & ~\[1612] ;
  assign n1214_1 = ~n5587 & ~n5588;
  assign n5590 = \[1594]  & n5586_1;
  assign n5591_1 = ~Ng261 & ~\[1594] ;
  assign n1219_1 = ~n5590 & ~n5591_1;
  assign n5593 = Ng853 & n5586_1;
  assign n5594 = ~Ng264 & ~Ng853;
  assign n1224_1 = ~n5593 & ~n5594;
  assign n5596_1 = ~Ng222 & ~\[1612] ;
  assign n5597 = ~n5099 & ~n5436_1;
  assign n5598 = ~n5445 & ~n5597;
  assign n5599 = ~n5201_1 & ~n5217;
  assign n5600 = ~n5207 & ~n5599;
  assign n5601_1 = ~n5580 & ~n5600;
  assign n5602 = ~n5561_1 & n5601_1;
  assign n5603 = ~n5236_1 & n5602;
  assign n5604 = n5236_1 & ~n5602;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606_1 = n5446_1 & ~n5605;
  assign n5607 = ~n5598 & ~n5606_1;
  assign n5608 = \[1612]  & ~n5607;
  assign n1229_1 = ~n5596_1 & ~n5608;
  assign n5610 = ~Ng225 & ~\[1594] ;
  assign n5611_1 = \[1594]  & ~n5607;
  assign n1234_1 = ~n5610 & ~n5611_1;
  assign n5613 = ~Ng228 & ~Ng853;
  assign n5614 = Ng853 & ~n5607;
  assign n1239_1 = ~n5613 & ~n5614;
  assign n5616_1 = ~Ng267 & ~\[1612] ;
  assign n5617 = ~n5113 & ~n5436_1;
  assign n5618 = ~n5445 & ~n5617;
  assign n5619 = n5236_1 & ~n5437;
  assign n5620 = ~n5438 & ~n5619;
  assign n5621_1 = n5602 & ~n5620;
  assign n5622 = ~n5241_1 & n5621_1;
  assign n5623 = n5241_1 & ~n5621_1;
  assign n5624 = ~n5622 & ~n5623;
  assign n5625 = n5446_1 & ~n5624;
  assign n5626_1 = ~n5618 & ~n5625;
  assign n5627 = \[1612]  & ~n5626_1;
  assign n1244_1 = ~n5616_1 & ~n5627;
  assign n5629 = ~Ng270 & ~\[1594] ;
  assign n5630 = \[1594]  & ~n5626_1;
  assign n1249_1 = ~n5629 & ~n5630;
  assign n5632 = ~Ng273 & ~Ng853;
  assign n5633 = Ng853 & ~n5626_1;
  assign n1254_1 = ~n5632 & ~n5633;
  assign n5635 = Ng853 & ~n5124;
  assign n5636_1 = Ng92 & n5635;
  assign n5637 = Ng92 & ~n5027;
  assign n5638 = ~n5635 & ~n5637;
  assign n1259_1 = ~n5636_1 & ~n5638;
  assign n5640 = ~Ng88 & ~n5636_1;
  assign n5641_1 = Ng88 & n5636_1;
  assign n5642 = n5027 & n5124;
  assign n5643 = ~n5641_1 & ~n5642;
  assign n1264_1 = ~n5640 & n5643;
  assign n5645 = Ng83 & n5641_1;
  assign n5646_1 = ~Ng83 & ~n5641_1;
  assign n5647 = ~n5642 & ~n5646_1;
  assign n1269 = ~n5645 & n5647;
  assign n5649 = Ng79 & n5645;
  assign n5650 = ~Ng79 & ~n5645;
  assign n5651_1 = ~n5642 & ~n5650;
  assign n1274 = ~n5649 & n5651_1;
  assign n5653 = Ng74 & n5649;
  assign n5654 = ~Ng74 & ~n5649;
  assign n5655 = ~n5642 & ~n5654;
  assign n1279 = ~n5653 & n5655;
  assign n5657 = Ng70 & n5653;
  assign n5658 = ~Ng70 & ~n5653;
  assign n5659 = ~n5642 & ~n5658;
  assign n1284_1 = ~n5657 & n5659;
  assign n5661_1 = Ng65 & n5657;
  assign n5662 = ~Ng65 & ~n5657;
  assign n5663 = ~n5642 & ~n5662;
  assign n1289 = ~n5661_1 & n5663;
  assign n5665 = Ng61 & n5661_1;
  assign n5666_1 = ~Ng61 & ~n5661_1;
  assign n5667 = ~n5642 & ~n5666_1;
  assign n1294 = ~n5665 & n5667;
  assign n5669 = Ng56 & n5665;
  assign n5670 = ~Ng56 & ~n5665;
  assign n5671_1 = ~n5642 & ~n5670;
  assign n1299 = ~n5669 & n5671_1;
  assign n5673 = Ng52 & n5669;
  assign n5674 = ~Ng52 & ~n5669;
  assign n5675 = ~n5673 & ~n5674;
  assign n1304 = ~n5642 & n5675;
  assign n5677 = n5195 & n5225;
  assign n5678 = n5194 & ~n5225;
  assign n5679 = ~n5189 & n5678;
  assign n5680 = ~n5124 & ~n5679;
  assign n5681_1 = ~n5677 & ~n5680;
  assign n5682 = \[1612]  & ~n5681_1;
  assign n5683 = ~Ng11499 & Ng853;
  assign n5684 = ~Ng11497 & \[1612] ;
  assign n5685 = ~Ng11498 & \[1594] ;
  assign n5686_1 = ~n5684 & ~n5685;
  assign n5687 = ~n5683 & n5686_1;
  assign n5688 = ~Ng11505 & Ng853;
  assign n5689 = ~Ng11503 & \[1612] ;
  assign n5690 = ~Ng11504 & \[1594] ;
  assign n5691_1 = ~n5689 & ~n5690;
  assign n5692 = ~n5688 & n5691_1;
  assign n5693 = ~Ng11502 & Ng853;
  assign n5694 = ~Ng11500 & \[1612] ;
  assign n5695 = ~Ng11501 & \[1594] ;
  assign n5696_1 = ~n5694 & ~n5695;
  assign n5697 = ~n5693 & n5696_1;
  assign n5698 = n5692 & ~n5697;
  assign n5699 = ~Ng11508 & Ng853;
  assign n5700 = ~Ng11506 & \[1612] ;
  assign n5701_1 = ~Ng11507 & \[1594] ;
  assign n5702 = ~n5700 & ~n5701_1;
  assign n5703 = ~n5699 & n5702;
  assign n5704 = ~n5698 & n5703;
  assign n5705 = ~n5687 & n5704;
  assign n5706_1 = ~Pg3229 & n5698;
  assign n5707 = Pg3229 & ~n5703;
  assign n5708 = ~n5706_1 & ~n5707;
  assign n5709 = ~n5705 & n5708;
  assign n5710 = n5682 & ~n5709;
  assign n5711_1 = ~Ng11497 & ~n5682;
  assign n1309 = ~n5710 & ~n5711_1;
  assign n5713 = \[1594]  & ~n5681_1;
  assign n5714 = ~n5709 & n5713;
  assign n5715 = ~Ng11498 & ~n5713;
  assign n1314_1 = ~n5714 & ~n5715;
  assign n5717 = Ng853 & ~n5681_1;
  assign n5718 = ~n5709 & n5717;
  assign n5719 = ~Ng11499 & ~n5717;
  assign n1319 = ~n5718 & ~n5719;
  assign n5721_1 = ~Ng11500 & ~n5682;
  assign n5722 = ~Pg3229 & ~n5687;
  assign n5723 = Pg3229 & n5687;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = ~n5692 & n5724;
  assign n5726_1 = ~n5698 & ~n5725;
  assign n5727 = n5682 & ~n5726_1;
  assign n1324_1 = ~n5721_1 & ~n5727;
  assign n5729 = n5713 & n5726_1;
  assign n5730 = Ng11501 & ~n5713;
  assign n1329_1 = n5729 | n5730;
  assign n5732 = n5717 & n5726_1;
  assign n5733 = Ng11502 & ~n5717;
  assign n1334_1 = n5732 | n5733;
  assign n5735 = n5697 & n5703;
  assign n5736_1 = n5724 & ~n5735;
  assign n5737 = n5697 & ~n5724;
  assign n5738 = ~n5736_1 & ~n5737;
  assign n5739 = n5682 & n5738;
  assign n5740 = ~Ng11503 & ~n5682;
  assign n1339_1 = ~n5739 & ~n5740;
  assign n5742 = Ng11504 & ~n5713;
  assign n5743 = n5713 & ~n5738;
  assign n1344_1 = n5742 | n5743;
  assign n5745 = n5717 & n5738;
  assign n5746_1 = ~Ng11505 & ~n5717;
  assign n1349_1 = ~n5745 & ~n5746_1;
  assign n5748 = n5692 & n5737;
  assign n5749 = n5682 & ~n5748;
  assign n5750 = Ng11506 & ~n5682;
  assign n1354 = n5749 | n5750;
  assign n5752 = n5713 & ~n5748;
  assign n5753 = Ng11507 & ~n5713;
  assign n1359 = n5752 | n5753;
  assign n5755 = n5717 & ~n5748;
  assign n5756_1 = Ng11508 & ~n5717;
  assign n1364 = n5755 | n5756_1;
  assign n5758 = ~n5113 & n5170;
  assign n5759 = ~n5099 & n5758;
  assign n5760 = Ng423 & Ng853;
  assign n5761_1 = Ng417 & \[1612] ;
  assign n5762 = Ng420 & \[1594] ;
  assign n5763 = ~n5761_1 & ~n5762;
  assign n1614_1 = n5760 | ~n5763;
  assign n5765 = ~n5759 & ~n1614_1;
  assign n5766_1 = ~n5433 & ~n1614_1;
  assign n5767 = n5759 & ~n5766_1;
  assign n5768 = ~n5765 & ~n5767;
  assign n5769 = Ng414 & Ng853;
  assign n5770 = Ng408 & \[1612] ;
  assign n5771_1 = Ng411 & \[1594] ;
  assign n5772 = ~n5770 & ~n5771_1;
  assign n5773 = ~n5769 & n5772;
  assign n5774 = Ng2257 & n5773;
  assign n5775 = n5768 & n5774;
  assign n5776_1 = ~Ng426 & Ng853;
  assign n5777 = ~Ng427 & \[1612] ;
  assign n5778 = ~Ng428 & \[1594] ;
  assign n5779 = ~n5777 & ~n5778;
  assign n5780 = ~n5776_1 & n5779;
  assign n5781_1 = n5768 & n5780;
  assign n5782 = Ng2257 & ~n5781_1;
  assign n5783 = ~n5773 & ~n5782;
  assign n5784 = ~n5775 & ~n5783;
  assign n5785 = \[1612]  & n5784;
  assign n5786_1 = ~Ng408 & ~\[1612] ;
  assign n1369 = ~n5785 & ~n5786_1;
  assign n5788 = \[1594]  & n5784;
  assign n5789 = ~Ng411 & ~\[1594] ;
  assign n1374_1 = ~n5788 & ~n5789;
  assign n5791_1 = Ng853 & n5784;
  assign n5792 = ~Ng414 & ~Ng853;
  assign n1379 = ~n5791_1 & ~n5792;
  assign n5794 = Ng2257 & ~n5773;
  assign n5795 = ~n5780 & n5794;
  assign n5796_1 = n5766_1 & ~n5795;
  assign n5797 = n1614_1 & ~n5795;
  assign n5798 = ~n5759 & ~n5797;
  assign n5799 = ~n5796_1 & ~n5798;
  assign n5800 = \[1612]  & n5799;
  assign n5801_1 = Ng417 & ~\[1612] ;
  assign n1384_1 = n5800 | n5801_1;
  assign n5803 = \[1594]  & n5799;
  assign n5804 = Ng420 & ~\[1594] ;
  assign n1389_1 = n5803 | n5804;
  assign n5806_1 = Ng853 & n5799;
  assign n5807 = Ng423 & ~Ng853;
  assign n1394_1 = n5806_1 | n5807;
  assign n5809 = n5781_1 & n5794;
  assign n5810 = \[1612]  & n5809;
  assign n5811_1 = \[1612]  & n5775;
  assign n5812 = ~Ng427 & ~n5811_1;
  assign n1399_1 = ~n5810 & ~n5812;
  assign n5814 = \[1594]  & n5809;
  assign n5815 = \[1594]  & n5775;
  assign n5816_1 = ~Ng428 & ~n5815;
  assign n1404_1 = ~n5814 & ~n5816_1;
  assign n5818 = Ng853 & n5809;
  assign n5819 = Ng853 & n5775;
  assign n5820_1 = ~Ng426 & ~n5819;
  assign n1409_1 = ~n5818 & ~n5820_1;
  assign n5822 = Ng429 & ~\[1612] ;
  assign n5823 = ~Ng177 & Ng853;
  assign n5824_1 = ~Ng178 & \[1612] ;
  assign n5825 = ~Ng179 & \[1594] ;
  assign n5826 = ~n5824_1 & ~n5825;
  assign n5827 = ~n5823 & n5826;
  assign n5828 = n5170 & ~n5827;
  assign n5829_1 = Ng2257 & n5828;
  assign n5830 = Ng435 & Ng853;
  assign n5831 = Ng429 & \[1612] ;
  assign n5832 = Ng432 & \[1594] ;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834_1 = ~n5830 & n5833;
  assign n5835 = ~Ng2257 & ~n5834_1;
  assign n5836 = ~n5829_1 & ~n5835;
  assign n5837 = \[1612]  & ~n5836;
  assign n1414 = n5822 | n5837;
  assign n5839_1 = Ng432 & ~\[1594] ;
  assign n5840 = \[1594]  & ~n5836;
  assign n1419 = n5839_1 | n5840;
  assign n5842 = Ng435 & ~Ng853;
  assign n5843 = Ng853 & ~n5836;
  assign n1424_1 = n5842 | n5843;
  assign n5845 = ~Ng438 & ~\[1612] ;
  assign n5846 = Ng444 & Ng853;
  assign n5847 = Ng438 & \[1612] ;
  assign n5848 = Ng441 & \[1594] ;
  assign n5849_1 = ~n5847 & ~n5848;
  assign n5850 = ~n5846 & n5849_1;
  assign n5851 = ~Ng447 & Ng853;
  assign n5852 = ~Ng448 & \[1612] ;
  assign n5853 = ~Ng449 & \[1594] ;
  assign n5854_1 = ~n5852 & ~n5853;
  assign n5855 = ~n5851 & n5854_1;
  assign n5856 = ~n5828 & ~n5850;
  assign n5857 = n5834_1 & ~n5856;
  assign n5858 = n5828 & n5850;
  assign n5859_1 = ~n5834_1 & ~n5858;
  assign n5860 = Ng2257 & ~n5859_1;
  assign n5861 = ~n5857 & n5860;
  assign n5862 = ~n5855 & n5861;
  assign n5863 = n5850 & n5862;
  assign n5864_1 = ~n5850 & ~n5862;
  assign n5865 = ~n5863 & ~n5864_1;
  assign n5866 = \[1612]  & n5865;
  assign n1429_1 = ~n5845 & ~n5866;
  assign n5868 = ~Ng441 & ~\[1594] ;
  assign n5869_1 = \[1594]  & n5865;
  assign n1434 = ~n5868 & ~n5869_1;
  assign n5871 = ~Ng444 & ~Ng853;
  assign n5872 = Ng853 & n5865;
  assign n1439_1 = ~n5871 & ~n5872;
  assign n5874_1 = n5855 & n5861;
  assign n5875 = \[1612]  & n5874_1;
  assign n5876 = n5834_1 & ~n5858;
  assign n5877 = ~n5834_1 & ~n5856;
  assign n5878 = Ng2257 & ~n5877;
  assign n5879_1 = ~n5876 & n5878;
  assign n5880 = \[1612]  & n5879_1;
  assign n5881 = ~Ng448 & ~n5880;
  assign n1444_1 = ~n5875 & ~n5881;
  assign n5883 = \[1594]  & n5874_1;
  assign n5884_1 = \[1594]  & n5879_1;
  assign n5885 = ~Ng449 & ~n5884_1;
  assign n1449 = ~n5883 & ~n5885;
  assign n5887 = Ng853 & n5874_1;
  assign n5888 = Ng853 & n5879_1;
  assign n5889_1 = ~Ng447 & ~n5888;
  assign n1454 = ~n5887 & ~n5889_1;
  assign n5891 = ~Ng312 & ~\[1612] ;
  assign n5892 = ~n5194 & ~n5225;
  assign n5893 = ~n5259 & ~n5892;
  assign n5894_1 = ~n5326_1 & ~n5893;
  assign n5895 = ~n5437 & ~n5894_1;
  assign n5896 = ~n5432 & ~n5895;
  assign n5897 = \[1612]  & ~n5896;
  assign n1459_1 = ~n5891 & ~n5897;
  assign n5899_1 = ~Ng313 & ~\[1594] ;
  assign n5900 = \[1594]  & ~n5896;
  assign n1464 = ~n5899_1 & ~n5900;
  assign n5902 = ~Ng314 & ~Ng853;
  assign n5903 = Ng853 & ~n5896;
  assign n1469_1 = ~n5902 & ~n5903;
  assign n5905 = ~Ng315 & ~\[1612] ;
  assign n5906 = n5326_1 & n5424;
  assign n5907 = n5189 & ~n5295;
  assign n5908 = n5268 & n5285;
  assign n5909_1 = n5318 & n5321_1;
  assign n5910 = n5290 & n5909_1;
  assign n5911 = n5908 & n5910;
  assign n5912 = ~n5264 & ~n5911;
  assign n5913 = Ng2257 & ~n5912;
  assign n5914_1 = n5907 & ~n5913;
  assign n5915 = ~n5424 & ~n5433;
  assign n5916 = ~n5189 & n5915;
  assign n5917 = ~n5914_1 & ~n5916;
  assign n5918 = ~n5906 & ~n5917;
  assign n5919_1 = n5257 & ~n5918;
  assign n5920 = n5265 & ~n5911;
  assign n5921 = n5907 & n5920;
  assign n5922 = ~n5225 & ~n5325;
  assign n5923 = ~n5921 & n5922;
  assign n5924_1 = ~n5195 & ~n5432;
  assign n5925 = ~n5678 & n5924_1;
  assign n5926 = ~n5923 & n5925;
  assign n5927 = ~n5919_1 & n5926;
  assign n5928 = \[1612]  & ~n5927;
  assign n1474_1 = ~n5905 & ~n5928;
  assign n5930 = ~Ng316 & ~\[1594] ;
  assign n5931 = \[1594]  & ~n5927;
  assign n1479_1 = ~n5930 & ~n5931;
  assign n5933 = ~Ng317 & ~Ng853;
  assign n5934_1 = Ng853 & ~n5927;
  assign n1484_1 = ~n5933 & ~n5934_1;
  assign n5936 = ~Ng318 & ~\[1612] ;
  assign n5937 = Ng2257 & n5225;
  assign n5938 = n5326_1 & n5937;
  assign n5939_1 = ~n5225 & n5913;
  assign n5940 = n5259 & ~n5939_1;
  assign n5941 = ~n5938 & n5940;
  assign n5942 = ~n5189 & n5920;
  assign n5943 = n5892 & n5942;
  assign n5944_1 = ~n5941 & ~n5943;
  assign n5945 = ~n5432 & ~n5944_1;
  assign n5946 = \[1612]  & ~n5945;
  assign n1489 = ~n5936 & ~n5946;
  assign n5948 = ~Ng319 & ~\[1594] ;
  assign n5949_1 = \[1594]  & ~n5945;
  assign n1494_1 = ~n5948 & ~n5949_1;
  assign n5951 = ~Ng320 & ~Ng853;
  assign n5952 = Ng853 & ~n5945;
  assign n1499 = ~n5951 & ~n5952;
  assign n5954_1 = ~n5258 & ~n5912;
  assign n5955 = n5019_1 & ~n5954_1;
  assign n5956 = Ng322 & ~n5955;
  assign n5957 = ~n5328 & n5418;
  assign n5958 = n5955 & ~n5957;
  assign n1504 = n5956 | n5958;
  assign n5960 = n5023 & ~n5954_1;
  assign n5961 = n5957 & n5960;
  assign n5962 = ~Ng323 & ~n5960;
  assign n1509_1 = ~n5961 & ~n5962;
  assign n5964_1 = n5027 & ~n5954_1;
  assign n5965 = Ng321 & ~n5964_1;
  assign n5966 = ~n5957 & n5964_1;
  assign n1514_1 = n5965 | n5966;
  assign n5968 = n5418 & n5431_1;
  assign n5969_1 = n5019_1 & ~n5968;
  assign n5970 = Ng403 & ~n5019_1;
  assign n1519_1 = n5969_1 | n5970;
  assign n5972 = n5023 & ~n5968;
  assign n5973 = Ng404 & ~n5023;
  assign n1524_1 = n5972 | n5973;
  assign n5975 = n5027 & ~n5968;
  assign n5976 = Ng402 & ~n5027;
  assign n1529_1 = n5975 | n5976;
  assign n5978 = ~Ng299 & ~Ng298;
  assign n5979_1 = Ng299 & Ng305;
  assign n5980 = ~\[1594]  & n5979_1;
  assign n1619_1 = n5978 | n5980;
  assign n5982 = ~Ng65 & ~n5206_1;
  assign n5983 = Ng88 & ~n5248;
  assign n5984_1 = ~Ng88 & n5248;
  assign n5985 = ~n5983 & ~n5984_1;
  assign n5986 = ~n5982 & ~n5985;
  assign n5987 = Ng70 & n5217;
  assign n5988 = Ng61 & n5201_1;
  assign n5989_1 = ~Ng61 & ~n5201_1;
  assign n5990 = ~n5988 & ~n5989_1;
  assign n5991 = ~n5987 & n5990;
  assign n5992 = n5986 & n5991;
  assign n5993 = ~Ng83 & n5230;
  assign n5994_1 = Ng83 & ~n5230;
  assign n5995 = ~n5993 & ~n5994_1;
  assign n5996 = n5992 & ~n5995;
  assign n5997 = ~Ng70 & ~n5217;
  assign n5998 = n5680 & ~n5997;
  assign n5999_1 = ~Ng74 & ~n5212;
  assign n6000 = Ng74 & n5212;
  assign n6001 = ~n5999_1 & ~n6000;
  assign n6002 = ~Ng92 & n5184;
  assign n6003 = Ng92 & ~n5184;
  assign n6004_1 = ~n6002 & ~n6003;
  assign n6005 = n6001 & ~n6004_1;
  assign n6006 = Ng65 & n5206_1;
  assign n6007 = ~Ng52 & n5241_1;
  assign n6008 = Ng52 & ~n5241_1;
  assign n6009_1 = ~n6007 & ~n6008;
  assign n6010 = ~n6006 & ~n6009_1;
  assign n6011 = n6005 & n6010;
  assign n6012 = n5998 & n6011;
  assign n6013 = ~Ng79 & ~n5253;
  assign n6014_1 = Ng79 & n5253;
  assign n6015 = ~n6013 & ~n6014_1;
  assign n6016 = Ng56 & ~n5236_1;
  assign n6017 = ~Ng56 & n5236_1;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019_1 = n6015 & ~n6018;
  assign n6020 = n6012 & n6019_1;
  assign n6021 = n5996 & n6020;
  assign n1624_1 = ~n5256_1 & ~n6021;
  assign n6023 = ~Ng3006 & ~Ng3010;
  assign n6024_1 = Ng2998 & n6023;
  assign n6025 = ~Ng2993 & Ng3002;
  assign n6026 = Ng3013 & Ng3024;
  assign n6027 = n6025 & n6026;
  assign n6028 = n6024_1 & n6027;
  assign n6029_1 = Ng3028 & ~Ng3032;
  assign n6030 = ~Ng3036 & n6029_1;
  assign n6031 = Ng3018 & n6030;
  assign n6032 = n6028 & n6031;
  assign n6033 = Ng1315 & ~n6032;
  assign n6034_1 = Ng554 & ~Ng1315;
  assign n1725 = n6033 | n6034_1;
  assign n6036 = Ng554 & Ng1315;
  assign n6037 = ~Ng557 & ~Ng1315;
  assign n1730 = ~n6036 & ~n6037;
  assign n6039_1 = Ng557 & Ng1315;
  assign n6040 = Ng510 & ~Ng1315;
  assign n1735_1 = n6039_1 | n6040;
  assign n6042 = Ng573 & Ng1315;
  assign n6043 = Ng569 & \[1605] ;
  assign n6044_1 = Ng571 & \[1603] ;
  assign n6045 = ~n6043 & ~n6044_1;
  assign n1740 = ~n6042 & n6045;
  assign n6047 = Ng486 & ~\[1612] ;
  assign n6048 = \[1612]  & ~n5850;
  assign n1807_1 = n6047 | n6048;
  assign n6050 = Ng487 & ~\[1594] ;
  assign n6051 = \[1594]  & ~n5850;
  assign n1812_1 = n6050 | n6051;
  assign n6053 = Ng488 & ~Ng853;
  assign n6054_1 = Ng853 & ~n5850;
  assign n1817_1 = n6053 | n6054_1;
  assign n6056 = ~Ng11512 & ~\[1612] ;
  assign n6057 = \[1612]  & ~n5679;
  assign n1822_1 = ~n6056 & ~n6057;
  assign n6059 = ~Ng11515 & ~\[1594] ;
  assign n6060 = \[1594]  & ~n5679;
  assign n1826_1 = ~n6059 & ~n6060;
  assign n6062 = ~Ng11516 & ~Ng853;
  assign n6063_1 = Ng853 & ~n5679;
  assign n1830_1 = ~n6062 & ~n6063_1;
  assign n6065 = ~Ng477 & ~\[1612] ;
  assign n6066 = \[1612]  & ~n5258;
  assign n1834_1 = ~n6065 & ~n6066;
  assign n6068 = ~Ng478 & ~\[1594] ;
  assign n6069 = \[1594]  & ~n5258;
  assign n1839 = ~n6068 & ~n6069;
  assign n6071 = ~Ng479 & ~Ng853;
  assign n6072_1 = Ng853 & ~n5258;
  assign n1844_1 = ~n6071 & ~n6072_1;
  assign n6074 = ~Ng480 & ~\[1612] ;
  assign n6075 = \[1612]  & n1614_1;
  assign n1849_1 = ~n6074 & ~n6075;
  assign n6077 = ~Ng484 & ~\[1594] ;
  assign n6078 = \[1594]  & n1614_1;
  assign n1854 = ~n6077 & ~n6078;
  assign n6080 = ~Ng464 & ~Ng853;
  assign n6081_1 = Ng853 & n1614_1;
  assign n1859_1 = ~n6080 & ~n6081_1;
  assign n6083 = ~Ng11517 & ~\[1612] ;
  assign n6084 = \[1612]  & ~n5677;
  assign n1864_1 = ~n6083 & ~n6084;
  assign n6086 = ~Ng11513 & ~\[1594] ;
  assign n6087 = \[1594]  & ~n5677;
  assign n1868_1 = ~n6086 & ~n6087;
  assign n6089 = ~Ng11514 & ~Ng853;
  assign n6090_1 = Ng853 & ~n5677;
  assign n1872_1 = ~n6089 & ~n6090_1;
  assign n6092 = Ng489 & Ng1315;
  assign n6093 = Ng565 & \[1605] ;
  assign n6094_1 = Ng567 & \[1603] ;
  assign n6095 = ~n6093 & ~n6094_1;
  assign n1876_1 = ~n6092 & n6095;
  assign n6097 = ~Ng479 & \[1605] ;
  assign n6098 = ~Ng477 & \[1603] ;
  assign n6099_1 = ~Ng478 & Ng1315;
  assign n6100 = ~n6098 & ~n6099_1;
  assign n1889_1 = ~n6097 & n6100;
  assign n6102 = ~Ng464 & \[1605] ;
  assign n6103_1 = ~Ng480 & \[1603] ;
  assign n6104 = ~Ng484 & Ng1315;
  assign n6105 = ~n6103_1 & ~n6104;
  assign n1903 = ~n6102 & n6105;
  assign n6107 = ~Ng488 & \[1605] ;
  assign n6108_1 = ~Ng486 & \[1603] ;
  assign n6109 = ~Ng487 & Ng1315;
  assign n6110 = ~n6108_1 & ~n6109;
  assign n1912_1 = ~n6107 & n6110;
  assign n6112_1 = Ng620 & Ng1315;
  assign n6113 = Ng614 & \[1605] ;
  assign n6114 = Ng617 & \[1603] ;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~n6112_1 & n6115;
  assign n6117_1 = Ng496 & Ng1315;
  assign n6118 = Ng490 & \[1605] ;
  assign n6119 = Ng493 & \[1603] ;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121_1 = ~n6117_1 & n6120;
  assign n6122 = Ng510 & n6121_1;
  assign n6123 = ~n6116 & n6122;
  assign n6124 = ~Ng3002 & ~Ng3024;
  assign n6125_1 = n6023 & n6124;
  assign n6126 = ~Ng3013 & n6125_1;
  assign n6127 = Ng611 & Ng1315;
  assign n6128 = Ng605 & \[1605] ;
  assign n6129_1 = Ng608 & \[1603] ;
  assign n6130 = ~n6128 & ~n6129_1;
  assign n6131 = ~n6127 & n6130;
  assign n6132 = ~n6121_1 & ~n6131;
  assign n6133 = ~n6126 & ~n6132;
  assign n2060_1 = n6123 | n6133;
  assign n6135 = \[1605]  & n2060_1;
  assign n6136 = ~Ng576 & ~n6135;
  assign n6137 = ~Ng584 & Ng1315;
  assign n6138 = ~Ng585 & \[1605] ;
  assign n6139_1 = ~Ng586 & \[1603] ;
  assign n6140 = ~n6138 & ~n6139_1;
  assign n6141 = ~n6137 & n6140;
  assign n6142 = Pg3229 & ~n6141;
  assign n6143 = ~Ng581 & Ng1315;
  assign n6144_1 = ~Ng582 & \[1605] ;
  assign n6145 = ~Ng583 & \[1603] ;
  assign n6146 = ~n6144_1 & ~n6145;
  assign n6147 = ~n6143 & n6146;
  assign n6148_1 = ~Ng578 & Ng1315;
  assign n6149 = ~Ng579 & \[1605] ;
  assign n6150 = ~Ng580 & \[1603] ;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152_1 = ~n6148_1 & n6151;
  assign n6153 = n6147 & ~n6152_1;
  assign n6154 = ~Ng575 & Ng1315;
  assign n6155 = ~Ng576 & \[1605] ;
  assign n6156_1 = ~Ng577 & \[1603] ;
  assign n6157 = ~n6155 & ~n6156_1;
  assign n6158 = ~n6154 & n6157;
  assign n6159 = n6141 & ~n6158;
  assign n6160_1 = ~n6153 & n6159;
  assign n6161 = ~Pg3229 & n6153;
  assign n6162 = ~n6160_1 & ~n6161;
  assign n6163 = ~n6142 & n6162;
  assign n6164_1 = n6135 & ~n6163;
  assign n1921 = ~n6136 & ~n6164_1;
  assign n6166 = \[1603]  & n2060_1;
  assign n6167 = ~n6163 & n6166;
  assign n6168_1 = ~Ng577 & ~n6166;
  assign n1926_1 = ~n6167 & ~n6168_1;
  assign n6170 = Ng1315 & n2060_1;
  assign n6171 = ~Ng575 & ~n6170;
  assign n6172_1 = ~n6163 & n6170;
  assign n1931 = ~n6171 & ~n6172_1;
  assign n6174 = ~Pg3229 & ~n6158;
  assign n6175 = Pg3229 & n6158;
  assign n6176_1 = ~n6174 & ~n6175;
  assign n6177 = ~n6147 & n6176_1;
  assign n6178 = ~n6153 & ~n6177;
  assign n6179 = n6135 & n6178;
  assign n6180_1 = Ng579 & ~n6135;
  assign n1936_1 = n6179 | n6180_1;
  assign n6182 = n6166 & n6178;
  assign n6183 = Ng580 & ~n6166;
  assign n1941_1 = n6182 | n6183;
  assign n6185 = n6170 & n6178;
  assign n6186 = Ng578 & ~n6170;
  assign n1946_1 = n6185 | n6186;
  assign n6188_1 = n6141 & n6152_1;
  assign n6189 = n6176_1 & ~n6188_1;
  assign n6190 = n6152_1 & ~n6176_1;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192_1 = n6135 & ~n6191;
  assign n6193 = Ng582 & ~n6135;
  assign n1951_1 = n6192_1 | n6193;
  assign n6195 = n6166 & ~n6191;
  assign n6196_1 = Ng583 & ~n6166;
  assign n1956_1 = n6195 | n6196_1;
  assign n6198 = n6170 & ~n6191;
  assign n6199 = Ng581 & ~n6170;
  assign n1961 = n6198 | n6199;
  assign n6201 = Ng585 & ~n6135;
  assign n6202 = n6147 & n6152_1;
  assign n6203 = ~n6176_1 & n6202;
  assign n6204_1 = n6135 & ~n6203;
  assign n1966_1 = n6201 | n6204_1;
  assign n6206 = Ng586 & ~n6166;
  assign n6207 = n6166 & ~n6203;
  assign n1971 = n6206 | n6207;
  assign n6209 = Ng584 & ~n6170;
  assign n6210 = n6170 & ~n6203;
  assign n1976_1 = n6209 | n6210;
  assign n6212_1 = ~Ng587 & ~\[1605] ;
  assign n6213 = Ng185 & Ng524;
  assign n6214 = ~n1740 & n6213;
  assign n6215 = Ng590 & \[1603] ;
  assign n6216_1 = Ng593 & Ng1315;
  assign n6217 = Ng587 & \[1605] ;
  assign n6218 = ~n6216_1 & ~n6217;
  assign n6219 = ~n6215 & n6218;
  assign n6220_1 = ~n6214 & n6219;
  assign n6221 = ~n6032 & ~n6220_1;
  assign n6222 = \[1605]  & ~n6221;
  assign n1981 = ~n6212_1 & ~n6222;
  assign n6224_1 = ~Ng590 & ~\[1603] ;
  assign n6225 = \[1603]  & ~n6221;
  assign n1986 = ~n6224_1 & ~n6225;
  assign n6227 = Ng593 & ~Ng1315;
  assign n6228_1 = n6033 & ~n6220_1;
  assign n1991_1 = n6227 | n6228_1;
  assign n6230 = ~Ng596 & ~\[1605] ;
  assign n6231 = Ng185 & Ng542;
  assign n6232_1 = ~n1876_1 & n6231;
  assign n6233 = Ng602 & Ng1315;
  assign n6234 = Ng599 & \[1603] ;
  assign n6235 = Ng596 & \[1605] ;
  assign n6236_1 = ~n6234 & ~n6235;
  assign n6237 = ~n6233 & n6236_1;
  assign n6238 = ~n6232_1 & n6237;
  assign n6239 = ~n6032 & ~n6238;
  assign n6240_1 = \[1605]  & ~n6239;
  assign n1996_1 = ~n6230 & ~n6240_1;
  assign n6242 = ~Ng599 & ~\[1603] ;
  assign n6243 = \[1603]  & ~n6239;
  assign n2001 = ~n6242 & ~n6243;
  assign n6245_1 = Ng602 & ~Ng1315;
  assign n6246 = n6033 & ~n6238;
  assign n2006_1 = n6245_1 | n6246;
  assign n6248 = Ng614 & ~\[1605] ;
  assign n6249 = ~n6032 & ~n6116;
  assign n6250_1 = ~n6220_1 & ~n6238;
  assign n6251 = n6032 & ~n6250_1;
  assign n6252 = Ng353 & Ng1315;
  assign n6253 = Ng349 & \[1605] ;
  assign n6254 = Ng351 & \[1603] ;
  assign n6255_1 = ~n6253 & ~n6254;
  assign n6256 = ~n6252 & n6255_1;
  assign n6257 = Ng383 & Ng1315;
  assign n6258 = Ng379 & \[1605] ;
  assign n6259 = Ng381 & \[1603] ;
  assign n6260_1 = ~n6258 & ~n6259;
  assign n6261 = ~n6257 & n6260_1;
  assign n6262 = Ng368 & Ng1315;
  assign n6263 = Ng364 & \[1605] ;
  assign n6264_1 = Ng366 & \[1603] ;
  assign n6265 = ~n6263 & ~n6264_1;
  assign n6266 = ~n6262 & n6265;
  assign n6267 = ~n6261 & ~n6266;
  assign n6268_1 = ~n6141 & n6267;
  assign n6269 = ~n6147 & n6266;
  assign n6270 = n6188_1 & n6261;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = Ng324 & Ng1315;
  assign n6273_1 = Ng394 & \[1605] ;
  assign n6274 = Ng396 & \[1603] ;
  assign n6275 = ~n6273_1 & ~n6274;
  assign n6276 = ~n6272 & n6275;
  assign n6277_1 = ~n6266 & ~n6276;
  assign n6278 = n6147 & n6277_1;
  assign n6279 = n6152_1 & n6278;
  assign n6280 = n6271 & ~n6279;
  assign n6281 = n6158 & ~n6280;
  assign n6282_1 = ~n6268_1 & ~n6281;
  assign n6283 = ~n6256 & ~n6282_1;
  assign n6284 = n6188_1 & n6267;
  assign n6285 = ~n6147 & n6277_1;
  assign n6286_1 = ~n6284 & ~n6285;
  assign n6287 = n6256 & ~n6286_1;
  assign n6288 = ~n6152_1 & n6256;
  assign n6289 = n6261 & n6288;
  assign n6290 = n6202 & n6276;
  assign n6291_1 = ~n6289 & ~n6290;
  assign n6292 = ~n6287 & n6291_1;
  assign n6293 = ~n6158 & ~n6292;
  assign n6294 = n6147 & n6256;
  assign n6295_1 = n6158 & ~n6261;
  assign n6296 = ~n6294 & ~n6295_1;
  assign n6297 = n6266 & ~n6296;
  assign n6298 = ~n6152_1 & n6297;
  assign n6299 = ~n6293 & ~n6298;
  assign n6300_1 = ~n6283 & n6299;
  assign n6301 = n6141 & ~n6256;
  assign n6302 = n6147 & ~n6301;
  assign n6303 = n6276 & ~n6302;
  assign n6304_1 = n6147 & ~n6256;
  assign n6305 = ~n6288 & ~n6304_1;
  assign n6306 = n6267 & n6305;
  assign n6307 = ~n6303 & ~n6306;
  assign n6308 = n6158 & ~n6307;
  assign n6309_1 = n6202 & ~n6266;
  assign n6310 = n6141 & ~n6309_1;
  assign n6311 = ~n6141 & ~n6276;
  assign n6312 = ~n6261 & ~n6311;
  assign n6313_1 = ~n6295_1 & ~n6312;
  assign n6314 = n6256 & n6313_1;
  assign n6315 = ~n6310 & n6314;
  assign n6316 = ~n6308 & ~n6315;
  assign n6317 = ~n6261 & ~n6278;
  assign n6318_1 = ~n6152_1 & ~n6269;
  assign n6319 = ~n6256 & n6318_1;
  assign n6320 = ~n6317 & n6319;
  assign n6321 = ~n6261 & ~n6302;
  assign n6322_1 = ~n6305 & ~n6321;
  assign n6323 = ~n6158 & n6266;
  assign n6324 = ~n6322_1 & n6323;
  assign n6325 = ~n6320 & ~n6324;
  assign n6326 = n6316 & n6325;
  assign n6327_1 = n6238 & n6326;
  assign n6328 = n6300_1 & ~n6327_1;
  assign n6329 = n6251 & n6328;
  assign n6330 = ~n6249 & ~n6329;
  assign n6331 = \[1605]  & ~n6330;
  assign n2011_1 = n6248 | n6331;
  assign n6333 = Ng617 & ~\[1603] ;
  assign n6334 = \[1603]  & ~n6330;
  assign n2016 = n6333 | n6334;
  assign n6336 = Ng620 & ~Ng1315;
  assign n6337_1 = Ng1315 & ~n6330;
  assign n2021_1 = n6336 | n6337_1;
  assign n6339 = Ng605 & ~\[1605] ;
  assign n6340 = ~n6032 & ~n6131;
  assign n6341 = n6220_1 & n6300_1;
  assign n6342_1 = n6251 & ~n6341;
  assign n6343 = n6326 & n6342_1;
  assign n6344 = ~n6340 & ~n6343;
  assign n6345 = \[1605]  & ~n6344;
  assign n2026_1 = n6339 | n6345;
  assign n6347 = Ng608 & ~\[1603] ;
  assign n6348 = \[1603]  & ~n6344;
  assign n2031_1 = n6347 | n6348;
  assign n6350_1 = Ng611 & ~Ng1315;
  assign n6351 = Ng1315 & ~n6344;
  assign n2036_1 = n6350_1 | n6351;
  assign n6353 = ~Ng490 & ~\[1605] ;
  assign n6354_1 = n6116 & n6122;
  assign n6355 = \[1605]  & ~n6354_1;
  assign n2041_1 = ~n6353 & ~n6355;
  assign n6357 = ~Ng493 & ~\[1603] ;
  assign n6358 = \[1603]  & ~n6354_1;
  assign n2046 = ~n6357 & ~n6358;
  assign n6360 = ~Ng496 & ~Ng1315;
  assign n6361 = Ng1315 & ~n6354_1;
  assign n2051_1 = ~n6360 & ~n6361;
  assign n6363 = Ng506 & ~Ng507;
  assign n6364_1 = \[1603]  & ~n6363;
  assign n6365 = ~Ng506 & ~Pg16297;
  assign n6366 = ~n6363 & ~n6365;
  assign n2065 = n6364_1 | n6366;
  assign n6368 = Pg3229 & Ng291;
  assign n6369_1 = ~Pg3229 & ~Ng305;
  assign n2113_1 = ~n6368 & ~n6369_1;
  assign n6371 = Ng510 & Ng1315;
  assign n6372 = Ng630 & ~Ng1315;
  assign n2123_1 = n6371 | n6372;
  assign n6374_1 = Ng1315 & ~n6126;
  assign n6375 = ~Ng659 & ~Ng1315;
  assign n2128 = ~n6374_1 & ~n6375;
  assign n6377 = Ng630 & \[1603] ;
  assign n6378 = ~Ng659 & Ng1315;
  assign n6379_1 = Ng640 & n6378;
  assign n6380 = ~Ng640 & ~n6378;
  assign n6381 = ~n6379_1 & ~n6380;
  assign n2133 = ~n6377 & n6381;
  assign n6383 = Ng633 & n6379_1;
  assign n6384_1 = ~Ng633 & ~n6379_1;
  assign n6385 = ~n6377 & ~n6384_1;
  assign n2138_1 = ~n6383 & n6385;
  assign n6387 = Ng653 & n6383;
  assign n6388_1 = ~Ng653 & ~n6383;
  assign n6389 = ~n6377 & ~n6388_1;
  assign n2143_1 = ~n6387 & n6389;
  assign n6391 = Ng646 & n6387;
  assign n6392_1 = ~Ng646 & ~n6387;
  assign n6393 = ~n6377 & ~n6392_1;
  assign n2148_1 = ~n6391 & n6393;
  assign n6395 = Ng660 & n6391;
  assign n6396_1 = ~Ng660 & ~n6391;
  assign n6397 = ~n6377 & ~n6396_1;
  assign n2153_1 = ~n6395 & n6397;
  assign n6399 = Ng672 & n6395;
  assign n6400_1 = ~Ng672 & ~n6395;
  assign n6401 = ~n6377 & ~n6400_1;
  assign n2158_1 = ~n6399 & n6401;
  assign n6403 = Ng666 & n6399;
  assign n6404_1 = ~Ng666 & ~n6399;
  assign n6405 = ~n6377 & ~n6404_1;
  assign n2163_1 = ~n6403 & n6405;
  assign n6407 = Ng679 & n6403;
  assign n6408 = ~Ng679 & ~n6403;
  assign n6409_1 = ~n6377 & ~n6408;
  assign n2168_1 = ~n6407 & n6409_1;
  assign n6411 = Ng686 & n6407;
  assign n6412 = ~Ng686 & ~n6407;
  assign n6413_1 = ~n6377 & ~n6412;
  assign n2173_1 = ~n6411 & n6413_1;
  assign n6415 = Ng692 & n6411;
  assign n6416 = ~Ng692 & ~n6411;
  assign n6417 = ~n6415 & ~n6416;
  assign n2178_1 = ~n6377 & n6417;
  assign n6419 = Ng525 & ~Ng659;
  assign n6420 = Ng538 & n6419;
  assign n6421 = \[1605]  & n6420;
  assign n6422 = Ng699 & ~n6421;
  assign n6423_1 = ~Ng640 & n6421;
  assign n2183_1 = n6422 | n6423_1;
  assign n6425 = \[1603]  & n6420;
  assign n6426 = Ng700 & ~n6425;
  assign n6427_1 = ~Ng640 & n6425;
  assign n2188 = n6426 | n6427_1;
  assign n6429 = Ng1315 & n6420;
  assign n6430 = Ng698 & ~n6429;
  assign n6431 = ~Ng640 & n6429;
  assign n2193 = n6430 | n6431;
  assign n6433 = Ng702 & ~n6421;
  assign n6434 = ~Ng633 & n6421;
  assign n2198_1 = n6433 | n6434;
  assign n6436_1 = Ng703 & ~n6425;
  assign n6437 = ~Ng633 & n6425;
  assign n2203_1 = n6436_1 | n6437;
  assign n6439 = Ng701 & ~n6429;
  assign n6440 = ~Ng633 & n6429;
  assign n2208_1 = n6439 | n6440;
  assign n6442 = Ng705 & ~n6421;
  assign n6443 = ~Ng653 & n6421;
  assign n2213 = n6442 | n6443;
  assign n6445 = Ng706 & ~n6425;
  assign n6446_1 = ~Ng653 & n6425;
  assign n2218 = n6445 | n6446_1;
  assign n6448 = Ng704 & ~n6429;
  assign n6449 = ~Ng653 & n6429;
  assign n2223_1 = n6448 | n6449;
  assign n6451_1 = Ng708 & ~n6421;
  assign n6452 = ~Ng646 & n6421;
  assign n2228 = n6451_1 | n6452;
  assign n6454 = Ng709 & ~n6425;
  assign n6455 = ~Ng646 & n6425;
  assign n2233_1 = n6454 | n6455;
  assign n6457 = Ng707 & ~n6429;
  assign n6458 = ~Ng646 & n6429;
  assign n2238 = n6457 | n6458;
  assign n6460 = Ng711 & ~n6421;
  assign n6461_1 = ~Ng660 & n6421;
  assign n2243_1 = n6460 | n6461_1;
  assign n6463 = Ng712 & ~n6425;
  assign n6464 = ~Ng660 & n6425;
  assign n2248 = n6463 | n6464;
  assign n6466_1 = Ng710 & ~n6429;
  assign n6467 = ~Ng660 & n6429;
  assign n2253_1 = n6466_1 | n6467;
  assign n6469 = Ng714 & ~n6421;
  assign n6470 = ~Ng672 & n6421;
  assign n2258 = n6469 | n6470;
  assign n6472 = Ng715 & ~n6425;
  assign n6473 = ~Ng672 & n6425;
  assign n2263 = n6472 | n6473;
  assign n6475 = Ng713 & ~n6429;
  assign n6476_1 = ~Ng672 & n6429;
  assign n2268 = n6475 | n6476_1;
  assign n6478 = Ng717 & ~n6421;
  assign n6479 = ~Ng666 & n6421;
  assign n2273 = n6478 | n6479;
  assign n6481_1 = Ng718 & ~n6425;
  assign n6482 = ~Ng666 & n6425;
  assign n2278_1 = n6481_1 | n6482;
  assign n6484 = Ng716 & ~n6429;
  assign n6485 = ~Ng666 & n6429;
  assign n2283 = n6484 | n6485;
  assign n6487 = Ng720 & ~n6421;
  assign n6488 = ~Ng679 & n6421;
  assign n2288 = n6487 | n6488;
  assign n6490 = Ng721 & ~n6425;
  assign n6491_1 = ~Ng679 & n6425;
  assign n2293 = n6490 | n6491_1;
  assign n6493 = Ng719 & ~n6429;
  assign n6494 = ~Ng679 & n6429;
  assign n2298 = n6493 | n6494;
  assign n6496_1 = Ng723 & ~n6421;
  assign n6497 = ~Ng686 & n6421;
  assign n2303 = n6496_1 | n6497;
  assign n6499 = Ng724 & ~n6425;
  assign n6500 = ~Ng686 & n6425;
  assign n2308 = n6499 | n6500;
  assign n6502 = Ng722 & ~n6429;
  assign n6503 = ~Ng686 & n6429;
  assign n2313 = n6502 | n6503;
  assign n6505 = Ng726 & ~n6421;
  assign n6506_1 = ~Ng692 & n6421;
  assign n2318 = n6505 | n6506_1;
  assign n6508 = Ng727 & ~n6425;
  assign n6509 = ~Ng692 & n6425;
  assign n2323_1 = n6508 | n6509;
  assign n6511_1 = Ng725 & ~n6429;
  assign n6512 = ~Ng692 & n6429;
  assign n2328 = n6511_1 | n6512;
  assign n6514 = Ng630 & \[1605] ;
  assign n6515 = ~n6116 & n6514;
  assign n6516_1 = ~Ng729 & ~n6514;
  assign n2333 = ~n6515 & ~n6516_1;
  assign n6518 = ~Ng730 & ~n6377;
  assign n6519 = ~n6116 & n6377;
  assign n2338 = ~n6518 & ~n6519;
  assign n6521_1 = Ng630 & Ng1315;
  assign n6522 = ~Ng728 & ~n6521_1;
  assign n6523 = ~n6116 & n6521_1;
  assign n2343 = ~n6522 & ~n6523;
  assign n6525 = ~n6131 & n6514;
  assign n6526_1 = ~Ng732 & ~n6514;
  assign n2348 = ~n6525 & ~n6526_1;
  assign n6528 = ~Ng733 & ~n6377;
  assign n6529 = ~n6131 & n6377;
  assign n2353 = ~n6528 & ~n6529;
  assign n6531_1 = ~Ng731 & ~n6521_1;
  assign n6532 = ~n6131 & n6521_1;
  assign n2358_1 = ~n6531_1 & ~n6532;
  assign n6534 = ~Ng716 & Ng1315;
  assign n6535 = ~Ng717 & \[1605] ;
  assign n6536_1 = ~Ng718 & \[1603] ;
  assign n6537 = ~n6535 & ~n6536_1;
  assign n6538 = ~n6534 & n6537;
  assign n6539 = ~Ng666 & ~n6538;
  assign n6540 = ~Ng725 & Ng1315;
  assign n6541_1 = ~Ng726 & \[1605] ;
  assign n6542 = ~Ng727 & \[1603] ;
  assign n6543 = ~n6541_1 & ~n6542;
  assign n6544 = ~n6540 & n6543;
  assign n6545 = Ng692 & n6544;
  assign n6546_1 = ~Ng692 & ~n6544;
  assign n6547 = ~n6545 & ~n6546_1;
  assign n6548 = ~n6539 & n6547;
  assign n6549 = ~Ng722 & Ng1315;
  assign n6550 = ~Ng723 & \[1605] ;
  assign n6551_1 = ~Ng724 & \[1603] ;
  assign n6552 = ~n6550 & ~n6551_1;
  assign n6553 = ~n6549 & n6552;
  assign n6554 = ~Ng686 & n6553;
  assign n6555 = Ng686 & ~n6553;
  assign n6556_1 = ~n6554 & ~n6555;
  assign n6557 = n6548 & ~n6556_1;
  assign n6558 = ~Ng704 & Ng1315;
  assign n6559 = ~Ng705 & \[1605] ;
  assign n6560 = ~Ng706 & \[1603] ;
  assign n6561_1 = ~n6559 & ~n6560;
  assign n6562 = ~n6558 & n6561_1;
  assign n6563 = Ng653 & ~n6562;
  assign n6564 = ~Ng653 & n6562;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566_1 = ~Ng707 & Ng1315;
  assign n6567 = ~Ng708 & \[1605] ;
  assign n6568 = ~Ng709 & \[1603] ;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = ~n6566_1 & n6569;
  assign n6571_1 = ~Ng646 & n6570;
  assign n6572 = Ng646 & ~n6570;
  assign n6573 = ~n6571_1 & ~n6572;
  assign n6574 = ~n6565 & ~n6573;
  assign n6575_1 = ~Ng713 & Ng1315;
  assign n6576 = ~Ng714 & \[1605] ;
  assign n6577 = ~Ng715 & \[1603] ;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = ~n6575_1 & n6578;
  assign n6580_1 = Ng672 & n6579;
  assign n6581 = ~Ng719 & Ng1315;
  assign n6582 = ~Ng720 & \[1605] ;
  assign n6583 = ~Ng721 & \[1603] ;
  assign n6584 = ~n6582 & ~n6583;
  assign n6585_1 = ~n6581 & n6584;
  assign n6586 = Ng679 & n6585_1;
  assign n6587 = ~Ng679 & ~n6585_1;
  assign n6588_1 = ~n6586 & ~n6587;
  assign n6589 = ~n6580_1 & n6588_1;
  assign n6590 = n6574 & n6589;
  assign n6591 = n6557 & n6590;
  assign n6592 = ~Ng672 & ~n6579;
  assign n6593_1 = ~Ng710 & Ng1315;
  assign n6594 = ~Ng711 & \[1605] ;
  assign n6595 = ~Ng712 & \[1603] ;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = ~n6593_1 & n6596;
  assign n6598_1 = Ng660 & n6597;
  assign n6599 = ~Ng660 & ~n6597;
  assign n6600 = ~n6598_1 & ~n6599;
  assign n6601 = ~n6592 & n6600;
  assign n6602 = Ng666 & n6538;
  assign n6603_1 = ~Ng701 & Ng1315;
  assign n6604 = ~Ng702 & \[1605] ;
  assign n6605 = ~Ng703 & \[1603] ;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~n6603_1 & n6606;
  assign n6608_1 = ~Ng633 & ~n6607;
  assign n6609 = ~n6602 & ~n6608_1;
  assign n6610 = Ng633 & n6607;
  assign n6611 = n6609 & ~n6610;
  assign n6612 = ~Ng698 & Ng1315;
  assign n6613_1 = ~Ng699 & \[1605] ;
  assign n6614 = ~Ng700 & \[1603] ;
  assign n6615 = ~n6613_1 & ~n6614;
  assign n6616 = ~n6612 & n6615;
  assign n6617 = Ng640 & ~n6616;
  assign n6618_1 = ~Ng640 & n6616;
  assign n6619 = ~n6617 & ~n6618_1;
  assign n6620 = n6611 & ~n6619;
  assign n6621 = n6601 & n6620;
  assign n6622 = n6591 & n6621;
  assign n6623_1 = ~Ng728 & Ng1315;
  assign n6624 = ~Ng731 & Ng1315;
  assign n6625 = ~Ng732 & \[1605] ;
  assign n6626 = ~Ng733 & \[1603] ;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628_1 = ~n6624 & n6627;
  assign n6629 = ~Ng729 & \[1605] ;
  assign n6630 = ~Ng730 & \[1603] ;
  assign n6631 = ~n6629 & ~n6630;
  assign n6632 = n6628_1 & n6631;
  assign n6633_1 = ~n6623_1 & n6632;
  assign n6634 = ~n6622 & n6633_1;
  assign n6635 = n6421 & n6634;
  assign n6636 = Ng735 & ~n6421;
  assign n2363 = n6635 | n6636;
  assign n6638_1 = n6425 & n6634;
  assign n6639 = Ng736 & ~n6425;
  assign n2368 = n6638_1 | n6639;
  assign n6641 = n6429 & n6634;
  assign n6642 = Ng734 & ~n6429;
  assign n2373 = n6641 | n6642;
  assign n6644 = ~Ng738 & ~n6421;
  assign n2378 = ~n6514 & ~n6644;
  assign n6646 = ~Ng739 & ~n6425;
  assign n2383 = ~n6377 & ~n6646;
  assign n6648_1 = ~Ng737 & ~n6429;
  assign n2388 = ~n6521_1 & ~n6648_1;
  assign n6650 = Ng818 & ~n5019_1;
  assign n6651 = ~Ng785 & n5019_1;
  assign n2405 = n6650 | n6651;
  assign n6653_1 = Ng819 & ~n5023;
  assign n6654 = ~Ng785 & n5023;
  assign n2410 = n6653_1 | n6654;
  assign n6656 = Ng817 & ~n5027;
  assign n6657 = ~Ng785 & n5027;
  assign n2415 = n6656 | n6657;
  assign n6659 = Ng821 & ~n5019_1;
  assign n6660 = ~Ng789 & n5019_1;
  assign n2420 = n6659 | n6660;
  assign n6662 = Ng822 & ~n5023;
  assign n6663_1 = ~Ng789 & n5023;
  assign n2425_1 = n6662 | n6663_1;
  assign n6665 = Ng820 & ~n5027;
  assign n6666 = ~Ng789 & n5027;
  assign n2430_1 = n6665 | n6666;
  assign n6668_1 = Ng830 & ~n5019_1;
  assign n6669 = ~Ng793 & n5019_1;
  assign n2435 = n6668_1 | n6669;
  assign n6671 = Ng831 & ~n5023;
  assign n6672 = ~Ng793 & n5023;
  assign n2440 = n6671 | n6672;
  assign n6674 = Ng829 & ~n5027;
  assign n6675 = ~Ng793 & n5027;
  assign n2445 = n6674 | n6675;
  assign n6677 = Ng833 & ~n5019_1;
  assign n6678_1 = ~Ng797 & n5019_1;
  assign n2450_1 = n6677 | n6678_1;
  assign n6680 = Ng834 & ~n5023;
  assign n6681 = ~Ng797 & n5023;
  assign n2455_1 = n6680 | n6681;
  assign n6683_1 = Ng832 & ~n5027;
  assign n6684 = ~Ng797 & n5027;
  assign n2460_1 = n6683_1 | n6684;
  assign n6686 = Ng836 & ~n5019_1;
  assign n6687 = ~Ng801 & n5019_1;
  assign n2465 = n6686 | n6687;
  assign n6689 = Ng837 & ~n5023;
  assign n6690 = ~Ng801 & n5023;
  assign n2470 = n6689 | n6690;
  assign n6692 = Ng835 & ~n5027;
  assign n6693_1 = ~Ng801 & n5027;
  assign n2475 = n6692 | n6693_1;
  assign n6695 = Ng839 & ~n5019_1;
  assign n6696 = ~Ng805 & n5019_1;
  assign n2480 = n6695 | n6696;
  assign n6698_1 = Ng840 & ~n5023;
  assign n6699 = ~Ng805 & n5023;
  assign n2485 = n6698_1 | n6699;
  assign n6701 = Ng838 & ~n5027;
  assign n6702 = ~Ng805 & n5027;
  assign n2490 = n6701 | n6702;
  assign n6704 = Ng842 & ~n5019_1;
  assign n6705 = ~Ng809 & n5019_1;
  assign n2495_1 = n6704 | n6705;
  assign n6707 = Ng843 & ~n5023;
  assign n6708_1 = ~Ng809 & n5023;
  assign n2500_1 = n6707 | n6708_1;
  assign n6710 = Ng841 & ~n5027;
  assign n6711 = ~Ng809 & n5027;
  assign n2505_1 = n6710 | n6711;
  assign n6713_1 = Ng845 & ~n5019_1;
  assign n6714 = ~Ng813 & n5019_1;
  assign n2510_1 = n6713_1 | n6714;
  assign n6716 = Ng846 & ~n5023;
  assign n6717 = ~Ng813 & n5023;
  assign n2515_1 = n6716 | n6717;
  assign n6719 = Ng844 & ~n5027;
  assign n6720 = ~Ng813 & n5027;
  assign n2520_1 = n6719 | n6720;
  assign n6722 = ~Ng848 & ~n5019_1;
  assign n6723_1 = Ng853 & ~Ng862;
  assign n6724 = \[1612]  & ~Ng863;
  assign n6725 = \[1594]  & ~Ng864;
  assign n6726 = ~n6724 & ~n6725;
  assign n6727 = ~n6723_1 & n6726;
  assign n6728_1 = n5019_1 & ~n6727;
  assign n2525 = ~n6722 & ~n6728_1;
  assign n6730 = n5023 & n6727;
  assign n6731 = Ng849 & ~n5023;
  assign n2530 = n6730 | n6731;
  assign n6733_1 = ~Ng847 & ~n5027;
  assign n6734 = n5027 & ~n6727;
  assign n2535 = ~n6733_1 & ~n6734;
  assign n6736 = ~Ng851 & ~n5019_1;
  assign n6737 = Ng853 & ~Ng859;
  assign n6738_1 = \[1612]  & ~Ng860;
  assign n6739 = \[1594]  & ~Ng861;
  assign n6740 = ~n6738_1 & ~n6739;
  assign n6741 = ~n6737 & n6740;
  assign n6742 = n5019_1 & ~n6741;
  assign n2540 = ~n6736 & ~n6742;
  assign n6744 = n5023 & n6741;
  assign n6745 = Ng852 & ~n5023;
  assign n2545_1 = n6744 | n6745;
  assign n6747 = ~Ng850 & ~n5027;
  assign n6748_1 = n5027 & ~n6741;
  assign n2550 = ~n6747 & ~n6748_1;
  assign n6750 = Ng813 & Ng801;
  assign n6751 = ~Ng805 & n6750;
  assign n6752 = ~Ng809 & n6751;
  assign n6753_1 = n5131_1 & n6752;
  assign n6754 = Ng857 & ~n5131_1;
  assign n2555 = n6753_1 | n6754;
  assign n6756 = n5138 & n6752;
  assign n6757 = Ng858 & ~n5138;
  assign n2560_1 = n6756 | n6757;
  assign n6759 = n5142 & n6752;
  assign n6760 = Ng856 & ~n5142;
  assign n2565 = n6759 | n6760;
  assign n6762 = Ng860 & ~n5131_1;
  assign n6763_1 = ~Ng789 & n5131_1;
  assign n2570 = n6762 | n6763_1;
  assign n6765 = Ng861 & ~n5138;
  assign n6766 = ~Ng789 & n5138;
  assign n2575_1 = n6765 | n6766;
  assign n6768_1 = Ng859 & ~n5142;
  assign n6769 = ~Ng789 & n5142;
  assign n2580 = n6768_1 | n6769;
  assign n6771 = Ng863 & ~n5131_1;
  assign n6772 = ~Ng785 & n5131_1;
  assign n2585 = n6771 | n6772;
  assign n6774 = Ng864 & ~n5138;
  assign n6775 = ~Ng785 & n5138;
  assign n2590 = n6774 | n6775;
  assign n6777 = Ng862 & ~n5142;
  assign n6778_1 = ~Ng785 & n5142;
  assign n2595_1 = n6777 | n6778_1;
  assign n6780 = Ng866 & ~n5131_1;
  assign n6781 = Ng789 & Ng785;
  assign n6782 = Ng797 & Ng793;
  assign n6783_1 = n6781 & n6782;
  assign n6784 = Ng809 & Ng805;
  assign n6785 = n6750 & n6784;
  assign n6786 = n6783_1 & n6785;
  assign n6787 = n5131_1 & ~n6786;
  assign n2600 = n6780 | n6787;
  assign n6789 = Ng867 & ~n5138;
  assign n6790 = n5138 & ~n6786;
  assign n2605 = n6789 | n6790;
  assign n6792 = Ng865 & ~n5142;
  assign n6793_1 = n5142 & ~n6786;
  assign n2610 = n6792 | n6793_1;
  assign n6795 = ~\[1612]  & ~Ng873;
  assign n6796 = Ng853 & Ng879;
  assign n6797 = \[1612]  & Ng873;
  assign n6798_1 = \[1594]  & Ng876;
  assign n6799 = ~n6797 & ~n6798_1;
  assign n6800 = ~n6796 & n6799;
  assign n6801 = Ng853 & ~Ng1007;
  assign n6802 = \[1612]  & ~Ng1005;
  assign n6803_1 = \[1594]  & ~Ng1006;
  assign n6804 = ~n6802 & ~n6803_1;
  assign n6805 = ~n6801 & n6804;
  assign n6806 = Ng853 & ~Ng1001;
  assign n6807 = \[1612]  & ~Ng999;
  assign n6808_1 = \[1594]  & ~Ng1000;
  assign n6809 = ~n6807 & ~n6808_1;
  assign n6810 = ~n6806 & n6809;
  assign n6811 = n6805 & n6810;
  assign n6812 = n6800 & n6811;
  assign n6813_1 = Ng853 & Ng951;
  assign n6814 = \[1612]  & Ng945;
  assign n6815 = \[1594]  & Ng948;
  assign n6816 = ~n6814 & ~n6815;
  assign n6817 = ~n6813_1 & n6816;
  assign n6818_1 = \[1612]  & Ng900;
  assign n6819 = \[1594]  & Ng903;
  assign n6820 = Ng853 & Ng906;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = ~n6818_1 & n6821;
  assign n6823_1 = n6817 & n6822;
  assign n6824 = Ng853 & Ng942;
  assign n6825 = \[1612]  & Ng936;
  assign n6826 = \[1594]  & Ng939;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828_1 = ~n6824 & n6827;
  assign n6829 = Ng853 & Ng897;
  assign n6830 = \[1612]  & Ng891;
  assign n6831 = \[1594]  & Ng894;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833_1 = ~n6829 & n6832;
  assign n6834 = n6828_1 & n6833_1;
  assign n6835 = n6823_1 & n6834;
  assign n6836 = n6812 & n6835;
  assign n6837 = Ng853 & ~Ng1004;
  assign n6838_1 = \[1612]  & ~Ng1002;
  assign n6839 = \[1594]  & ~Ng1003;
  assign n6840 = ~n6838_1 & ~n6839;
  assign n6841 = ~n6837 & n6840;
  assign n6842 = Ng853 & Ng888;
  assign n6843_1 = \[1612]  & Ng882;
  assign n6844 = \[1594]  & Ng885;
  assign n6845 = ~n6843_1 & ~n6844;
  assign n6846 = ~n6842 & n6845;
  assign n6847 = n6841 & n6846;
  assign n6848_1 = Ng853 & Ng960;
  assign n6849 = \[1612]  & Ng954;
  assign n6850 = \[1594]  & Ng957;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = ~n6848_1 & n6851;
  assign n6853_1 = Ng853 & Ng924;
  assign n6854 = \[1612]  & Ng918;
  assign n6855 = \[1594]  & Ng921;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = ~n6853_1 & n6856;
  assign n6858_1 = n6852 & n6857;
  assign n6859 = n6847 & n6858_1;
  assign n6860 = Ng853 & Ng933;
  assign n6861 = \[1612]  & Ng927;
  assign n6862 = \[1594]  & Ng930;
  assign n6863_1 = ~n6861 & ~n6862;
  assign n6864 = ~n6860 & n6863_1;
  assign n6865 = Ng853 & Ng915;
  assign n6866 = \[1612]  & Ng909;
  assign n6867 = \[1594]  & Ng912;
  assign n6868_1 = ~n6866 & ~n6867;
  assign n6869 = ~n6865 & n6868_1;
  assign n6870 = n6864 & n6869;
  assign n6871 = n6859 & n6870;
  assign n6872 = n6836 & n6871;
  assign n6873_1 = ~n6810 & n6841;
  assign n6874 = ~n6805 & n6873_1;
  assign n6875 = n6805 & ~n6810;
  assign n6876 = Ng853 & ~Ng856;
  assign n6877 = \[1594]  & ~Ng858;
  assign n6878_1 = \[1612]  & ~Ng857;
  assign n6879 = ~n6877 & ~n6878_1;
  assign n6880 = ~n6876 & n6879;
  assign n6881 = Ng2257 & ~n6880;
  assign n6882 = ~Ng797 & ~n6864;
  assign n6883_1 = Ng797 & n6864;
  assign n6884 = ~n6882 & ~n6883_1;
  assign n6885 = ~Ng805 & ~n6828_1;
  assign n6886 = Ng805 & n6828_1;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888_1 = n6884 & n6887;
  assign n6889 = ~n6741 & ~n6852;
  assign n6890 = n6741 & n6852;
  assign n6891 = ~n6889 & ~n6890;
  assign n6892 = ~Ng813 & ~n6817;
  assign n6893_1 = Ng813 & n6817;
  assign n6894 = ~n6892 & ~n6893_1;
  assign n6895 = ~n6891 & n6894;
  assign n6896 = ~Ng789 & ~n6857;
  assign n6897 = Ng789 & n6857;
  assign n6898_1 = ~n6896 & ~n6897;
  assign n6899 = ~n6895 & ~n6898_1;
  assign n6900 = n6884 & ~n6891;
  assign n6901 = n6894 & n6898_1;
  assign n6902 = ~n6887 & ~n6901;
  assign n6903_1 = ~n6900 & n6902;
  assign n6904 = ~n6899 & ~n6903_1;
  assign n6905 = ~n6888_1 & ~n6904;
  assign n6906 = n6887 & n6894;
  assign n6907 = n6884 & n6898_1;
  assign n6908_1 = n6891 & ~n6907;
  assign n6909 = ~n6906 & n6908_1;
  assign n6910 = ~n6905 & ~n6909;
  assign n6911 = n6881 & ~n6910;
  assign n6912 = n6727 & ~n6869;
  assign n6913_1 = ~n6727 & n6869;
  assign n6914 = ~n6912 & ~n6913_1;
  assign n6915 = ~Ng809 & ~n6822;
  assign n6916 = Ng809 & n6822;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918_1 = ~Ng801 & ~n6833_1;
  assign n6919 = Ng801 & n6833_1;
  assign n6920 = ~n6918_1 & ~n6919;
  assign n6921 = n6917 & n6920;
  assign n6922 = ~Ng785 & ~n6800;
  assign n6923_1 = Ng785 & n6800;
  assign n6924 = ~n6922 & ~n6923_1;
  assign n6925 = ~Ng793 & ~n6846;
  assign n6926 = Ng793 & n6846;
  assign n6927_1 = ~n6925 & ~n6926;
  assign n6928 = n6924 & n6927_1;
  assign n6929 = ~n6921 & ~n6928;
  assign n6930 = ~n6914 & n6929;
  assign n6931 = n6920 & n6927_1;
  assign n6932_1 = n6914 & n6917;
  assign n6933 = ~n6924 & ~n6932_1;
  assign n6934 = ~n6931 & n6933;
  assign n6935 = n6917 & n6924;
  assign n6936 = n6914 & n6927_1;
  assign n6937_1 = ~n6920 & ~n6936;
  assign n6938 = ~n6935 & n6937_1;
  assign n6939 = ~n6934 & ~n6938;
  assign n6940 = ~n6930 & n6939;
  assign n6941 = n6881 & ~n6940;
  assign n6942_1 = ~n6911 & ~n6941;
  assign n6943 = n6875 & n6942_1;
  assign n6944 = ~n6874 & ~n6943;
  assign n6945 = Ng853 & ~Ng838;
  assign n6946 = \[1612]  & ~Ng839;
  assign n6947_1 = \[1594]  & ~Ng840;
  assign n6948 = ~n6946 & ~n6947_1;
  assign n6949 = ~n6945 & n6948;
  assign n6950 = ~Ng805 & ~n6949;
  assign n6951 = Ng853 & ~Ng844;
  assign n6952_1 = \[1612]  & ~Ng845;
  assign n6953 = \[1594]  & ~Ng846;
  assign n6954 = ~n6952_1 & ~n6953;
  assign n6955 = ~n6951 & n6954;
  assign n6956 = ~Ng813 & ~n6955;
  assign n6957_1 = Ng853 & ~Ng850;
  assign n6958 = \[1612]  & ~Ng851;
  assign n6959 = \[1594]  & ~Ng852;
  assign n6960 = ~n6958 & ~n6959;
  assign n6961 = ~n6957_1 & n6960;
  assign n6962_1 = ~n6741 & n6961;
  assign n6963 = ~n6956 & ~n6962_1;
  assign n6964 = ~n6950 & n6963;
  assign n6965 = Ng813 & n6955;
  assign n6966 = Ng805 & n6949;
  assign n6967_1 = n6881 & ~n6966;
  assign n6968 = ~n6965 & n6967_1;
  assign n6969 = n6964 & n6968;
  assign n6970 = Ng853 & ~Ng841;
  assign n6971 = \[1612]  & ~Ng842;
  assign n6972_1 = \[1594]  & ~Ng843;
  assign n6973 = ~n6971 & ~n6972_1;
  assign n6974 = ~n6970 & n6973;
  assign n6975 = Ng809 & n6974;
  assign n6976 = Ng853 & ~Ng829;
  assign n6977_1 = \[1594]  & ~Ng831;
  assign n6978 = \[1612]  & ~Ng830;
  assign n6979 = ~n6977_1 & ~n6978;
  assign n6980 = ~n6976 & n6979;
  assign n6981 = ~Ng793 & ~n6980;
  assign n6982_1 = ~n6975 & ~n6981;
  assign n6983 = Ng793 & n6980;
  assign n6984 = n6982_1 & ~n6983;
  assign n6985 = n6969 & n6984;
  assign n6986 = Ng853 & ~Ng832;
  assign n6987_1 = \[1594]  & ~Ng834;
  assign n6988 = \[1612]  & ~Ng833;
  assign n6989 = ~n6987_1 & ~n6988;
  assign n6990 = ~n6986 & n6989;
  assign n6991 = Ng797 & n6990;
  assign n6992_1 = ~Ng797 & ~n6990;
  assign n6993 = ~n6991 & ~n6992_1;
  assign n6994 = Ng853 & ~Ng847;
  assign n6995 = \[1612]  & ~Ng848;
  assign n6996 = \[1594]  & ~Ng849;
  assign n6997_1 = ~n6995 & ~n6996;
  assign n6998 = ~n6994 & n6997_1;
  assign n6999 = n6727 & n6998;
  assign n7000 = ~n6727 & ~n6998;
  assign n7001 = ~n6999 & ~n7000;
  assign n7002_1 = Ng853 & ~Ng820;
  assign n7003 = \[1612]  & ~Ng821;
  assign n7004 = \[1594]  & ~Ng822;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n7002_1 & n7005;
  assign n7007_1 = ~Ng789 & n7006;
  assign n7008 = Ng789 & ~n7006;
  assign n7009 = ~n7007_1 & ~n7008;
  assign n7010 = ~n7001 & ~n7009;
  assign n7011 = n6993 & n7010;
  assign n7012_1 = n6741 & ~n6961;
  assign n7013 = ~Ng809 & ~n6974;
  assign n7014 = ~n7012_1 & ~n7013;
  assign n7015 = Ng853 & ~Ng835;
  assign n7016 = \[1594]  & ~Ng837;
  assign n7017_1 = \[1612]  & ~Ng836;
  assign n7018 = ~n7016 & ~n7017_1;
  assign n7019 = ~n7015 & n7018;
  assign n7020 = ~Ng801 & n7019;
  assign n7021 = Ng801 & ~n7019;
  assign n7022_1 = ~n7020 & ~n7021;
  assign n7023 = n7014 & ~n7022_1;
  assign n7024 = Ng853 & ~Ng817;
  assign n7025 = \[1612]  & ~Ng818;
  assign n7026 = \[1594]  & ~Ng819;
  assign n7027_1 = ~n7025 & ~n7026;
  assign n7028 = ~n7024 & n7027_1;
  assign n7029 = ~Ng785 & n7028;
  assign n7030 = Ng785 & ~n7028;
  assign n7031 = ~n7029 & ~n7030;
  assign n7032_1 = n7023 & ~n7031;
  assign n7033 = n7011 & n7032_1;
  assign n7034 = n6985 & n7033;
  assign n7035 = \[1594]  & ~Ng1010;
  assign n7036 = Ng853 & ~Ng1008;
  assign n7037_1 = \[1612]  & ~Ng1009;
  assign n7038 = ~n7036 & ~n7037_1;
  assign n7039 = ~n7035 & n7038;
  assign n7040 = n7034 & ~n7039;
  assign n7041 = n6841 & n7040;
  assign n7042_1 = ~n6944 & n7041;
  assign n7043 = Ng853 & ~Ng1089;
  assign n7044 = \[1612]  & ~Ng1090;
  assign n7045 = \[1594]  & ~Ng1091;
  assign n7046 = ~n7044 & ~n7045;
  assign n7047_1 = ~n7043 & n7046;
  assign n7048 = n7034 & ~n7047_1;
  assign n7049 = Ng2257 & n6880;
  assign n7050 = ~n6810 & n7049;
  assign n7051 = ~n7048 & ~n7050;
  assign n7052_1 = ~n7042_1 & n7051;
  assign n7053 = ~n6852 & ~n6864;
  assign n7054 = ~n6846 & n7053;
  assign n7055 = n6811 & ~n6841;
  assign n7056 = ~n6869 & n7055;
  assign n7057_1 = n6800 & n6835;
  assign n7058 = n7056 & n7057_1;
  assign n7059 = n7054 & n7058;
  assign n7060 = ~n6857 & n7059;
  assign n7061 = n7052_1 & ~n7060;
  assign n7062_1 = ~n6872 & n7061;
  assign n7063 = Ng785 & ~n7052_1;
  assign n7064 = ~n7062_1 & ~n7063;
  assign n7065 = ~n6800 & ~n6811;
  assign n7066 = ~n6812 & ~n7065;
  assign n7067_1 = n7061 & n7066;
  assign n7068 = ~n7064 & ~n7067_1;
  assign n7069 = \[1612]  & ~n7068;
  assign n2615 = ~n6795 & ~n7069;
  assign n7071 = ~\[1594]  & ~Ng876;
  assign n7072_1 = \[1594]  & ~n7068;
  assign n2620_1 = ~n7071 & ~n7072_1;
  assign n7074 = ~Ng853 & ~Ng879;
  assign n7075 = Ng853 & ~n7068;
  assign n2625 = ~n7074 & ~n7075;
  assign n7077_1 = ~\[1612]  & ~Ng918;
  assign n7078 = Ng789 & ~n7052_1;
  assign n7079 = ~n7061 & ~n7078;
  assign n7080 = n6800 & n6841;
  assign n7081 = ~n6800 & ~n6841;
  assign n7082_1 = ~n7080 & ~n7081;
  assign n7083 = n6811 & ~n7082_1;
  assign n7084 = ~n6857 & n7083;
  assign n7085 = n6857 & ~n7083;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087_1 = n7062_1 & ~n7086;
  assign n7088 = ~n7079 & ~n7087_1;
  assign n7089 = \[1612]  & ~n7088;
  assign n2630 = ~n7077_1 & ~n7089;
  assign n7091 = ~\[1594]  & ~Ng921;
  assign n7092_1 = \[1594]  & ~n7088;
  assign n2635 = ~n7091 & ~n7092_1;
  assign n7094 = ~Ng853 & ~Ng924;
  assign n7095 = Ng853 & ~n7088;
  assign n2640 = ~n7094 & ~n7095;
  assign n7097_1 = ~\[1612]  & ~Ng882;
  assign n7098 = Ng793 & ~n7052_1;
  assign n7099 = ~n7061 & ~n7098;
  assign n7100 = n6857 & n7080;
  assign n7101 = ~n6857 & n7081;
  assign n7102_1 = ~n7100 & ~n7101;
  assign n7103 = n6811 & ~n7102_1;
  assign n7104 = n6846 & n7103;
  assign n7105 = ~n6846 & ~n7103;
  assign n7106 = ~n7104 & ~n7105;
  assign n7107_1 = n7062_1 & n7106;
  assign n7108 = ~n7099 & ~n7107_1;
  assign n7109 = \[1612]  & ~n7108;
  assign n2645 = ~n7097_1 & ~n7109;
  assign n7111 = ~\[1594]  & ~Ng885;
  assign n7112_1 = \[1594]  & ~n7108;
  assign n2650 = ~n7111 & ~n7112_1;
  assign n7114 = ~Ng853 & ~Ng888;
  assign n7115 = Ng853 & ~n7108;
  assign n2655 = ~n7114 & ~n7115;
  assign n7117_1 = ~\[1612]  & ~Ng927;
  assign n7118 = Ng797 & ~n7052_1;
  assign n7119 = ~n7061 & ~n7118;
  assign n7120 = ~n6841 & ~n6846;
  assign n7121 = ~n6847 & ~n7120;
  assign n7122_1 = n7103 & ~n7121;
  assign n7123 = ~n6864 & n7122_1;
  assign n7124 = n6864 & ~n7122_1;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = n7062_1 & ~n7125;
  assign n7127_1 = ~n7119 & ~n7126;
  assign n7128 = \[1612]  & ~n7127_1;
  assign n2660 = ~n7117_1 & ~n7128;
  assign n7130 = ~\[1594]  & ~Ng930;
  assign n7131 = \[1594]  & ~n7127_1;
  assign n2665 = ~n7130 & ~n7131;
  assign n7133 = ~Ng853 & ~Ng933;
  assign n7134 = Ng853 & ~n7127_1;
  assign n2670 = ~n7133 & ~n7134;
  assign n7136 = Ng801 & ~n7052_1;
  assign n7137_1 = ~n6864 & ~n7055;
  assign n7138 = n6864 & n7055;
  assign n7139 = ~n7137_1 & ~n7138;
  assign n7140 = n7122_1 & n7139;
  assign n7141 = n6833_1 & n7140;
  assign n7142_1 = ~n6833_1 & ~n7140;
  assign n7143 = ~n7141 & ~n7142_1;
  assign n7144 = n7062_1 & ~n7143;
  assign n7145 = ~n7136 & ~n7144;
  assign n7146 = \[1612]  & n7145;
  assign n7147_1 = ~\[1612]  & ~Ng891;
  assign n2675 = ~n7146 & ~n7147_1;
  assign n7149 = \[1594]  & n7145;
  assign n7150 = ~\[1594]  & ~Ng894;
  assign n2680_1 = ~n7149 & ~n7150;
  assign n7152_1 = Ng853 & n7145;
  assign n7153 = ~Ng853 & ~Ng897;
  assign n2685 = ~n7152_1 & ~n7153;
  assign n7155 = ~\[1612]  & Ng936;
  assign n7156 = Ng805 & ~n7052_1;
  assign n7157_1 = ~n6833_1 & n7055;
  assign n7158 = n6833_1 & ~n7055;
  assign n7159 = ~n7157_1 & ~n7158;
  assign n7160 = n7140 & ~n7159;
  assign n7161_1 = n6828_1 & n7160;
  assign n7162 = ~n6828_1 & ~n7160;
  assign n7163 = ~n7161_1 & ~n7162;
  assign n7164_1 = n7062_1 & ~n7163;
  assign n7165 = ~n7156 & ~n7164_1;
  assign n7166 = \[1612]  & ~n7165;
  assign n2690 = n7155 | n7166;
  assign n7168_1 = ~\[1594]  & Ng939;
  assign n7169 = \[1594]  & ~n7165;
  assign n2695_1 = n7168_1 | n7169;
  assign n7171 = ~Ng853 & Ng942;
  assign n7172 = Ng853 & ~n7165;
  assign n2700 = n7171 | n7172;
  assign n7174 = Ng809 & ~n7052_1;
  assign n7175 = n6828_1 & n7055;
  assign n7176 = n7123 & n7157_1;
  assign n7177_1 = ~n7161_1 & ~n7176;
  assign n7178 = ~n7175 & ~n7177_1;
  assign n7179 = n6822 & n7178;
  assign n7180 = ~n6822 & ~n7178;
  assign n7181_1 = ~n7179 & ~n7180;
  assign n7182 = n7062_1 & ~n7181_1;
  assign n7183 = ~n7174 & ~n7182;
  assign n7184 = \[1612]  & n7183;
  assign n7185_1 = ~\[1612]  & ~Ng900;
  assign n2705_1 = ~n7184 & ~n7185_1;
  assign n7187 = \[1594]  & n7183;
  assign n7188 = ~\[1594]  & ~Ng903;
  assign n2710_1 = ~n7187 & ~n7188;
  assign n7190 = Ng853 & n7183;
  assign n7191 = ~Ng853 & ~Ng906;
  assign n2715_1 = ~n7190 & ~n7191;
  assign n7193_1 = Ng813 & ~n7052_1;
  assign n7194 = n6822 & ~n7055;
  assign n7195 = ~n6822 & n7055;
  assign n7196 = ~n7194 & ~n7195;
  assign n7197_1 = n7178 & ~n7196;
  assign n7198 = ~n6817 & n7197_1;
  assign n7199 = n6817 & ~n7197_1;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201_1 = n7062_1 & n7200;
  assign n7202 = ~n7193_1 & ~n7201_1;
  assign n7203 = \[1612]  & n7202;
  assign n7204 = ~\[1612]  & ~Ng945;
  assign n2720 = ~n7203 & ~n7204;
  assign n7206 = \[1594]  & n7202;
  assign n7207 = ~\[1594]  & ~Ng948;
  assign n2725_1 = ~n7206 & ~n7207;
  assign n7209 = Ng853 & n7202;
  assign n7210_1 = ~Ng853 & ~Ng951;
  assign n2730_1 = ~n7209 & ~n7210_1;
  assign n7212 = ~\[1612]  & ~Ng909;
  assign n7213 = ~n6727 & ~n7052_1;
  assign n7214_1 = ~n7061 & ~n7213;
  assign n7215 = ~n6817 & ~n6828_1;
  assign n7216 = ~n6823_1 & ~n7215;
  assign n7217 = ~n7196 & ~n7216;
  assign n7218 = ~n7177_1 & n7217;
  assign n7219_1 = ~n6869 & n7218;
  assign n7220 = n6869 & ~n7218;
  assign n7221 = ~n7219_1 & ~n7220;
  assign n7222 = n7062_1 & ~n7221;
  assign n7223_1 = ~n7214_1 & ~n7222;
  assign n7224 = \[1612]  & ~n7223_1;
  assign n2735_1 = ~n7212 & ~n7224;
  assign n7226 = ~\[1594]  & ~Ng912;
  assign n7227_1 = \[1594]  & ~n7223_1;
  assign n2740_1 = ~n7226 & ~n7227_1;
  assign n7229 = ~Ng853 & ~Ng915;
  assign n7230 = Ng853 & ~n7223_1;
  assign n2745_1 = ~n7229 & ~n7230;
  assign n7232 = ~\[1612]  & ~Ng954;
  assign n7233 = ~n6741 & ~n7052_1;
  assign n7234 = ~n7061 & ~n7233;
  assign n7235_1 = n6869 & ~n7055;
  assign n7236 = ~n7056 & ~n7235_1;
  assign n7237 = n7218 & ~n7236;
  assign n7238 = ~n6852 & n7237;
  assign n7239_1 = n6852 & ~n7237;
  assign n7240 = ~n7238 & ~n7239_1;
  assign n7241 = n7062_1 & ~n7240;
  assign n7242 = ~n7234 & ~n7241;
  assign n7243_1 = \[1612]  & ~n7242;
  assign n2750_1 = ~n7232 & ~n7243_1;
  assign n7245 = ~\[1594]  & ~Ng957;
  assign n7246 = \[1594]  & ~n7242;
  assign n2755_1 = ~n7245 & ~n7246;
  assign n7248 = ~Ng853 & ~Ng960;
  assign n7249 = Ng853 & ~n7242;
  assign n2760_1 = ~n7248 & ~n7249;
  assign n7251_1 = Ng780 & n5635;
  assign n7252 = Ng780 & ~n5027;
  assign n7253 = ~n5635 & ~n7252;
  assign n2765_1 = ~n7251_1 & ~n7253;
  assign n7255 = Ng776 & n7251_1;
  assign n7256_1 = ~Ng776 & ~n7251_1;
  assign n7257 = ~n5642 & ~n7256_1;
  assign n2770_1 = ~n7255 & n7257;
  assign n7259 = Ng771 & n7255;
  assign n7260 = ~Ng771 & ~n7255;
  assign n7261_1 = ~n5642 & ~n7260;
  assign n2775_1 = ~n7259 & n7261_1;
  assign n7263 = Ng767 & n7259;
  assign n7264 = ~Ng767 & ~n7259;
  assign n7265 = ~n5642 & ~n7264;
  assign n2780_1 = ~n7263 & n7265;
  assign n7267 = Ng762 & n7263;
  assign n7268 = ~Ng762 & ~n7263;
  assign n7269 = ~n5642 & ~n7268;
  assign n2785_1 = ~n7267 & n7269;
  assign n7271 = Ng758 & n7267;
  assign n7272 = ~Ng758 & ~n7267;
  assign n7273 = ~n5642 & ~n7272;
  assign n2790_1 = ~n7271 & n7273;
  assign n7275 = Ng753 & n7271;
  assign n7276 = ~Ng753 & ~n7271;
  assign n7277 = ~n5642 & ~n7276;
  assign n2795_1 = ~n7275 & n7277;
  assign n7279 = Ng749 & n7275;
  assign n7280 = ~Ng749 & ~n7275;
  assign n7281 = ~n5642 & ~n7280;
  assign n2800_1 = ~n7279 & n7281;
  assign n7283 = Ng744 & n7279;
  assign n7284 = ~Ng744 & ~n7279;
  assign n7285 = ~n5642 & ~n7284;
  assign n2805_1 = ~n7283 & n7285;
  assign n7287 = Ng740 & n7283;
  assign n7288 = ~Ng740 & ~n7283;
  assign n7289 = ~n7287 & ~n7288;
  assign n2810_1 = ~n5642 & n7289;
  assign n7291 = n6811 & n6841;
  assign n7292 = n6810 & ~n6841;
  assign n7293 = ~n6805 & n7292;
  assign n7294 = ~n5124 & ~n7293;
  assign n7295 = ~n7291 & ~n7294;
  assign n7296 = \[1612]  & ~n7295;
  assign n7297 = Ng853 & ~Ng11526;
  assign n7298 = \[1612]  & ~Ng11524;
  assign n7299 = \[1594]  & ~Ng11525;
  assign n7300 = ~n7298 & ~n7299;
  assign n7301 = ~n7297 & n7300;
  assign n7302 = Ng853 & ~Ng11532;
  assign n7303 = \[1612]  & ~Ng11530;
  assign n7304 = \[1594]  & ~Ng11531;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~n7302 & n7305;
  assign n7307 = Ng853 & ~Ng11529;
  assign n7308 = \[1612]  & ~Ng11527;
  assign n7309 = \[1594]  & ~Ng11528;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~n7307 & n7310;
  assign n7312 = n7306 & ~n7311;
  assign n7313 = Ng853 & ~Ng11535;
  assign n7314 = \[1612]  & ~Ng11533;
  assign n7315 = \[1594]  & ~Ng11534;
  assign n7316 = ~n7314 & ~n7315;
  assign n7317 = ~n7313 & n7316;
  assign n7318 = ~n7312 & n7317;
  assign n7319 = ~n7301 & n7318;
  assign n7320 = ~Pg3229 & n7312;
  assign n7321 = Pg3229 & ~n7317;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = ~n7319 & n7322;
  assign n7324 = n7296 & ~n7323;
  assign n7325 = ~Ng11524 & ~n7296;
  assign n2815_1 = ~n7324 & ~n7325;
  assign n7327 = \[1594]  & ~n7295;
  assign n7328 = ~n7323 & n7327;
  assign n7329 = ~Ng11525 & ~n7327;
  assign n2820_1 = ~n7328 & ~n7329;
  assign n7331 = Ng853 & ~n7295;
  assign n7332 = ~n7323 & n7331;
  assign n7333 = ~Ng11526 & ~n7331;
  assign n2825_1 = ~n7332 & ~n7333;
  assign n7335 = ~Ng11527 & ~n7296;
  assign n7336 = ~Pg3229 & ~n7301;
  assign n7337 = Pg3229 & n7301;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~n7306 & n7338;
  assign n7340 = ~n7312 & ~n7339;
  assign n7341 = n7296 & ~n7340;
  assign n2830_1 = ~n7335 & ~n7341;
  assign n7343 = n7327 & n7340;
  assign n7344 = Ng11528 & ~n7327;
  assign n2835 = n7343 | n7344;
  assign n7346 = ~Ng11529 & ~n7331;
  assign n7347 = n7331 & ~n7340;
  assign n2840_1 = ~n7346 & ~n7347;
  assign n7349 = n7311 & ~n7338;
  assign n7350 = n7311 & n7317;
  assign n7351 = n7338 & ~n7350;
  assign n7352 = ~n7349 & ~n7351;
  assign n7353 = n7296 & n7352;
  assign n7354 = ~Ng11530 & ~n7296;
  assign n2845_1 = ~n7353 & ~n7354;
  assign n7356 = n7327 & ~n7352;
  assign n7357 = Ng11531 & ~n7327;
  assign n2850_1 = n7356 | n7357;
  assign n7359 = n7331 & n7352;
  assign n7360 = ~Ng11532 & ~n7331;
  assign n2855_1 = ~n7359 & ~n7360;
  assign n7362 = n7306 & n7349;
  assign n7363 = n7296 & ~n7362;
  assign n7364 = Ng11533 & ~n7296;
  assign n2860_1 = n7363 | n7364;
  assign n7366 = n7327 & ~n7362;
  assign n7367 = Ng11534 & ~n7327;
  assign n2865_1 = n7366 | n7367;
  assign n7369 = n7331 & ~n7362;
  assign n7370 = Ng11535 & ~n7331;
  assign n2870_1 = n7369 | n7370;
  assign n7372 = ~n6741 & n6786;
  assign n7373 = ~n6727 & n7372;
  assign n7374 = Ng853 & Ng1110;
  assign n7375 = \[1612]  & Ng1104;
  assign n7376 = \[1594]  & Ng1107;
  assign n7377 = ~n7375 & ~n7376;
  assign n3120_1 = n7374 | ~n7377;
  assign n7379 = ~n7049 & ~n3120_1;
  assign n7380 = n7373 & n7379;
  assign n7381 = ~n7373 & n3120_1;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = Ng853 & Ng1101;
  assign n7384 = \[1612]  & Ng1095;
  assign n7385 = \[1594]  & Ng1098;
  assign n7386 = ~n7384 & ~n7385;
  assign n7387 = ~n7383 & n7386;
  assign n7388 = Ng2257 & n7387;
  assign n7389 = ~n7382 & n7388;
  assign n7390 = Ng853 & ~Ng1113;
  assign n7391 = \[1612]  & ~Ng1114;
  assign n7392 = \[1594]  & ~Ng1115;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 = ~n7390 & n7393;
  assign n7395 = ~n7382 & n7394;
  assign n7396 = Ng2257 & ~n7395;
  assign n7397 = ~n7387 & ~n7396;
  assign n7398 = ~n7389 & ~n7397;
  assign n7399 = \[1612]  & n7398;
  assign n7400 = ~\[1612]  & ~Ng1095;
  assign n2875_1 = ~n7399 & ~n7400;
  assign n7402 = \[1594]  & n7398;
  assign n7403 = ~\[1594]  & ~Ng1098;
  assign n2880_1 = ~n7402 & ~n7403;
  assign n7405 = Ng853 & n7398;
  assign n7406 = ~Ng853 & ~Ng1101;
  assign n2885_1 = ~n7405 & ~n7406;
  assign n7408 = ~\[1612]  & Ng1104;
  assign n7409 = Ng2257 & ~n7387;
  assign n7410 = ~n7394 & n7409;
  assign n7411 = n3120_1 & ~n7410;
  assign n7412 = ~n7049 & ~n7410;
  assign n7413 = n7373 & ~n7412;
  assign n7414 = ~n7411 & ~n7413;
  assign n7415 = \[1612]  & ~n7414;
  assign n2890_1 = n7408 | n7415;
  assign n7417 = ~\[1594]  & Ng1107;
  assign n7418 = \[1594]  & ~n7414;
  assign n2895_1 = n7417 | n7418;
  assign n7420 = ~Ng853 & Ng1110;
  assign n7421 = Ng853 & ~n7414;
  assign n2900_1 = n7420 | n7421;
  assign n7423 = n7395 & n7409;
  assign n7424 = \[1612]  & n7423;
  assign n7425 = \[1612]  & n7389;
  assign n7426 = ~Ng1114 & ~n7425;
  assign n2905_1 = ~n7424 & ~n7426;
  assign n7428 = \[1594]  & n7423;
  assign n7429 = \[1594]  & n7389;
  assign n7430 = ~Ng1115 & ~n7429;
  assign n2910_1 = ~n7428 & ~n7430;
  assign n7432 = Ng853 & n7423;
  assign n7433 = Ng853 & n7389;
  assign n7434 = ~Ng1113 & ~n7433;
  assign n2915_1 = ~n7432 & ~n7434;
  assign n7436 = ~\[1612]  & Ng1116;
  assign n7437 = Ng853 & ~Ng865;
  assign n7438 = \[1612]  & ~Ng866;
  assign n7439 = \[1594]  & ~Ng867;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = ~n7437 & n7440;
  assign n7442 = n6786 & ~n7441;
  assign n7443 = Ng2257 & n7442;
  assign n7444 = Ng853 & Ng1122;
  assign n7445 = \[1612]  & Ng1116;
  assign n7446 = \[1594]  & Ng1119;
  assign n7447 = ~n7445 & ~n7446;
  assign n7448 = ~n7444 & n7447;
  assign n7449 = ~Ng2257 & ~n7448;
  assign n7450 = ~n7443 & ~n7449;
  assign n7451 = \[1612]  & ~n7450;
  assign n2920_1 = n7436 | n7451;
  assign n7453 = ~\[1594]  & Ng1119;
  assign n7454 = \[1594]  & ~n7450;
  assign n2925_1 = n7453 | n7454;
  assign n7456 = ~Ng853 & Ng1122;
  assign n7457 = Ng853 & ~n7450;
  assign n2930_1 = n7456 | n7457;
  assign n7459 = ~\[1612]  & ~Ng1125;
  assign n7460 = Ng853 & Ng1131;
  assign n7461 = \[1612]  & Ng1125;
  assign n7462 = \[1594]  & Ng1128;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = ~n7460 & n7463;
  assign n7465 = Ng853 & ~Ng1134;
  assign n7466 = \[1612]  & ~Ng1135;
  assign n7467 = \[1594]  & ~Ng1136;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = ~n7465 & n7468;
  assign n7470 = ~n7442 & ~n7464;
  assign n7471 = n7448 & ~n7470;
  assign n7472 = n7442 & n7464;
  assign n7473 = ~n7448 & ~n7472;
  assign n7474 = Ng2257 & ~n7473;
  assign n7475 = ~n7471 & n7474;
  assign n7476 = ~n7469 & n7475;
  assign n7477 = n7464 & n7476;
  assign n7478 = ~n7464 & ~n7476;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = \[1612]  & n7479;
  assign n2935_1 = ~n7459 & ~n7480;
  assign n7482 = ~\[1594]  & ~Ng1128;
  assign n7483 = \[1594]  & n7479;
  assign n2940_1 = ~n7482 & ~n7483;
  assign n7485 = ~Ng853 & ~Ng1131;
  assign n7486 = Ng853 & n7479;
  assign n2945_1 = ~n7485 & ~n7486;
  assign n7488 = n7469 & n7475;
  assign n7489 = \[1612]  & n7488;
  assign n7490 = n7448 & ~n7472;
  assign n7491 = ~n7448 & ~n7470;
  assign n7492 = Ng2257 & ~n7491;
  assign n7493 = ~n7490 & n7492;
  assign n7494 = \[1612]  & n7493;
  assign n7495 = ~Ng1135 & ~n7494;
  assign n2950_1 = ~n7489 & ~n7495;
  assign n7497 = \[1594]  & n7488;
  assign n7498 = \[1594]  & n7493;
  assign n7499 = ~Ng1136 & ~n7498;
  assign n2955_1 = ~n7497 & ~n7499;
  assign n7501 = Ng853 & n7488;
  assign n7502 = Ng853 & n7493;
  assign n7503 = ~Ng1134 & ~n7502;
  assign n2960_1 = ~n7501 & ~n7503;
  assign n7505 = ~\[1612]  & ~Ng999;
  assign n7506 = ~n6810 & ~n6841;
  assign n7507 = ~n6875 & ~n7506;
  assign n7508 = ~n6942_1 & ~n7507;
  assign n7509 = ~n7055 & ~n7508;
  assign n7510 = ~n7048 & ~n7509;
  assign n7511 = \[1612]  & ~n7510;
  assign n2965_1 = ~n7505 & ~n7511;
  assign n7513 = ~\[1594]  & ~Ng1000;
  assign n7514 = \[1594]  & ~n7510;
  assign n2970_1 = ~n7513 & ~n7514;
  assign n7516 = ~Ng853 & ~Ng1001;
  assign n7517 = Ng853 & ~n7510;
  assign n2975_1 = ~n7516 & ~n7517;
  assign n7519 = ~\[1612]  & ~Ng1002;
  assign n7520 = ~n6941 & n7040;
  assign n7521 = n6898_1 & n6914;
  assign n7522 = n6900 & n7521;
  assign n7523 = n6906 & n6928;
  assign n7524 = n7522 & n7523;
  assign n7525 = n6921 & n7524;
  assign n7526 = ~n6880 & ~n7525;
  assign n7527 = Ng2257 & ~n7526;
  assign n7528 = n6805 & ~n6911;
  assign n7529 = ~n7527 & n7528;
  assign n7530 = ~n7040 & ~n7049;
  assign n7531 = ~n6805 & n7530;
  assign n7532 = ~n7529 & ~n7531;
  assign n7533 = ~n7520 & ~n7532;
  assign n7534 = n6873_1 & ~n7533;
  assign n7535 = n6881 & ~n7525;
  assign n7536 = n7528 & n7535;
  assign n7537 = ~n6841 & ~n6941;
  assign n7538 = ~n7536 & n7537;
  assign n7539 = ~n6811 & ~n7048;
  assign n7540 = ~n7292 & n7539;
  assign n7541 = ~n7538 & n7540;
  assign n7542 = ~n7534 & n7541;
  assign n7543 = \[1612]  & ~n7542;
  assign n2980_1 = ~n7519 & ~n7543;
  assign n7545 = ~\[1594]  & ~Ng1003;
  assign n7546 = \[1594]  & ~n7542;
  assign n2985_1 = ~n7545 & ~n7546;
  assign n7548 = ~Ng853 & ~Ng1004;
  assign n7549 = Ng853 & ~n7542;
  assign n2990_1 = ~n7548 & ~n7549;
  assign n7551 = ~\[1612]  & ~Ng1005;
  assign n7552 = Ng2257 & n6841;
  assign n7553 = n6942_1 & n7552;
  assign n7554 = ~n6841 & n7527;
  assign n7555 = n6875 & ~n7554;
  assign n7556 = ~n7553 & n7555;
  assign n7557 = ~n6805 & n7535;
  assign n7558 = n7506 & n7557;
  assign n7559 = ~n7556 & ~n7558;
  assign n7560 = ~n7048 & ~n7559;
  assign n7561 = \[1612]  & ~n7560;
  assign n2995_1 = ~n7551 & ~n7561;
  assign n7563 = ~\[1594]  & ~Ng1006;
  assign n7564 = \[1594]  & ~n7560;
  assign n3000_1 = ~n7563 & ~n7564;
  assign n7566 = ~Ng853 & ~Ng1007;
  assign n7567 = Ng853 & ~n7560;
  assign n3005_1 = ~n7566 & ~n7567;
  assign n7569 = ~n6874 & ~n7526;
  assign n7570 = n5019_1 & ~n7569;
  assign n7571 = ~n6944 & n7034;
  assign n7572 = n7570 & ~n7571;
  assign n7573 = Ng1009 & ~n7570;
  assign n3010_1 = n7572 | n7573;
  assign n7575 = n5023 & ~n7569;
  assign n7576 = n7571 & n7575;
  assign n7577 = ~Ng1010 & ~n7575;
  assign n3015 = ~n7576 & ~n7577;
  assign n7579 = n5027 & ~n7569;
  assign n7580 = Ng1008 & ~n7579;
  assign n7581 = ~n7571 & n7579;
  assign n3020_1 = n7580 | n7581;
  assign n7583 = n7034 & n7047_1;
  assign n7584 = n5019_1 & ~n7583;
  assign n7585 = Ng1090 & ~n5019_1;
  assign n3025 = n7584 | n7585;
  assign n7587 = n5023 & ~n7583;
  assign n7588 = Ng1091 & ~n5023;
  assign n3030_1 = n7587 | n7588;
  assign n7590 = n5027 & ~n7583;
  assign n7591 = Ng1089 & ~n5027;
  assign n3035_1 = n7590 | n7591;
  assign n7593 = ~Ng986 & Ng985;
  assign n7594 = ~\[1594]  & Ng992;
  assign n7595 = \[1594]  & n5978;
  assign n7596 = Ng986 & ~n7595;
  assign n7597 = ~n7594 & n7596;
  assign n3125_1 = ~n7593 & ~n7597;
  assign n7599 = Ng780 & n6800;
  assign n7600 = Ng744 & n6869;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = ~Ng771 & ~n6846;
  assign n7603 = ~Ng776 & ~n6857;
  assign n7604 = Ng749 & n6817;
  assign n7605 = ~n7603 & ~n7604;
  assign n7606 = Ng771 & n6846;
  assign n7607 = n7605 & ~n7606;
  assign n7608 = ~n7602 & n7607;
  assign n7609 = n7601 & n7608;
  assign n7610 = Ng776 & n6857;
  assign n7611 = ~Ng780 & ~n6800;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~Ng749 & ~n6817;
  assign n7614 = n7612 & ~n7613;
  assign n7615 = ~Ng744 & ~n6869;
  assign n7616 = ~Ng767 & ~n6864;
  assign n7617 = Ng767 & n6864;
  assign n7618 = ~n7616 & ~n7617;
  assign n7619 = Ng762 & n6833_1;
  assign n7620 = ~Ng762 & ~n6833_1;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = n7618 & n7621;
  assign n7623 = ~n7615 & n7622;
  assign n7624 = Ng740 & ~n6852;
  assign n7625 = ~Ng740 & n6852;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = Ng753 & n6822;
  assign n7628 = ~Ng753 & ~n6822;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~n7626 & n7629;
  assign n7631 = ~Ng758 & n6828_1;
  assign n7632 = Ng758 & ~n6828_1;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = n7630 & ~n7633;
  assign n7635 = n7623 & n7634;
  assign n7636 = n7614 & n7635;
  assign n7637 = n7294 & n7636;
  assign n7638 = n7609 & n7637;
  assign n3130_1 = ~n6872 & ~n7638;
  assign n7640 = Ng1240 & ~Ng1315;
  assign n3231_1 = n6033 | n7640;
  assign n7642 = Ng1240 & Ng1315;
  assign n7643 = ~Ng1243 & ~Ng1315;
  assign n3236_1 = ~n7642 & ~n7643;
  assign n7645 = Ng1243 & Ng1315;
  assign n7646 = Ng1196 & ~Ng1315;
  assign n3241_1 = n7645 | n7646;
  assign n7648 = Ng1259 & Ng1315;
  assign n7649 = Ng1255 & \[1605] ;
  assign n7650 = Ng1257 & \[1603] ;
  assign n7651 = ~n7649 & ~n7650;
  assign n3246_1 = ~n7648 & n7651;
  assign n7653 = ~\[1612]  & Ng1173;
  assign n7654 = \[1612]  & ~n7464;
  assign n3313_1 = n7653 | n7654;
  assign n7656 = ~\[1594]  & Ng1174;
  assign n7657 = \[1594]  & ~n7464;
  assign n3318_1 = n7656 | n7657;
  assign n7659 = ~Ng853 & Ng1175;
  assign n7660 = Ng853 & ~n7464;
  assign n3323_1 = n7659 | n7660;
  assign n7662 = ~\[1612]  & ~Ng11539;
  assign n7663 = \[1612]  & ~n7293;
  assign n3328_1 = ~n7662 & ~n7663;
  assign n7665 = ~\[1594]  & ~Ng11542;
  assign n7666 = \[1594]  & ~n7293;
  assign n3332_1 = ~n7665 & ~n7666;
  assign n7668 = ~Ng853 & ~Ng11543;
  assign n7669 = Ng853 & ~n7293;
  assign n3336_1 = ~n7668 & ~n7669;
  assign n7671 = ~\[1612]  & ~Ng1164;
  assign n7672 = \[1612]  & ~n6874;
  assign n3340_1 = ~n7671 & ~n7672;
  assign n7674 = ~\[1594]  & ~Ng1165;
  assign n7675 = \[1594]  & ~n6874;
  assign n3345_1 = ~n7674 & ~n7675;
  assign n7677 = ~Ng853 & ~Ng1166;
  assign n7678 = Ng853 & ~n6874;
  assign n3350_1 = ~n7677 & ~n7678;
  assign n7680 = ~\[1612]  & ~Ng1167;
  assign n7681 = \[1612]  & n3120_1;
  assign n3355_1 = ~n7680 & ~n7681;
  assign n7683 = ~\[1594]  & ~Ng1171;
  assign n7684 = \[1594]  & n3120_1;
  assign n3360_1 = ~n7683 & ~n7684;
  assign n7686 = ~Ng853 & ~Ng1151;
  assign n7687 = Ng853 & n3120_1;
  assign n3365_1 = ~n7686 & ~n7687;
  assign n7689 = ~\[1612]  & ~Ng11544;
  assign n7690 = \[1612]  & ~n7291;
  assign n3370_1 = ~n7689 & ~n7690;
  assign n7692 = ~\[1594]  & ~Ng11540;
  assign n7693 = \[1594]  & ~n7291;
  assign n3374_1 = ~n7692 & ~n7693;
  assign n7695 = ~Ng853 & ~Ng11541;
  assign n7696 = Ng853 & ~n7291;
  assign n3378_1 = ~n7695 & ~n7696;
  assign n7698 = Ng1176 & Ng1315;
  assign n7699 = Ng1251 & \[1605] ;
  assign n7700 = Ng1253 & \[1603] ;
  assign n7701 = ~n7699 & ~n7700;
  assign n3382_1 = ~n7698 & n7701;
  assign n7703 = ~Ng1166 & \[1605] ;
  assign n7704 = ~Ng1164 & \[1603] ;
  assign n7705 = ~Ng1165 & Ng1315;
  assign n7706 = ~n7704 & ~n7705;
  assign n3395_1 = ~n7703 & n7706;
  assign n7708 = ~Ng1151 & \[1605] ;
  assign n7709 = ~Ng1167 & \[1603] ;
  assign n7710 = ~Ng1171 & Ng1315;
  assign n7711 = ~n7709 & ~n7710;
  assign n3409_1 = ~n7708 & n7711;
  assign n7713 = ~Ng1175 & \[1605] ;
  assign n7714 = ~Ng1173 & \[1603] ;
  assign n7715 = ~Ng1174 & Ng1315;
  assign n7716 = ~n7714 & ~n7715;
  assign n3418_1 = ~n7713 & n7716;
  assign n7718 = Ng1306 & Ng1315;
  assign n7719 = Ng1300 & \[1605] ;
  assign n7720 = Ng1303 & \[1603] ;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = ~n7718 & n7721;
  assign n7723 = Ng1183 & Ng1315;
  assign n7724 = Ng1177 & \[1605] ;
  assign n7725 = Ng1180 & \[1603] ;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = ~n7723 & n7726;
  assign n7728 = Ng1196 & n7727;
  assign n7729 = ~n7722 & n7728;
  assign n7730 = Ng1297 & Ng1315;
  assign n7731 = Ng1291 & \[1605] ;
  assign n7732 = Ng1294 & \[1603] ;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = ~n7730 & n7733;
  assign n7735 = ~n7727 & ~n7734;
  assign n7736 = ~n6126 & ~n7735;
  assign n3566_1 = n7729 | n7736;
  assign n7738 = \[1605]  & n3566_1;
  assign n7739 = ~Ng1262 & ~n7738;
  assign n7740 = ~Ng1270 & Ng1315;
  assign n7741 = ~Ng1271 & \[1605] ;
  assign n7742 = ~Ng1272 & \[1603] ;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = ~n7740 & n7743;
  assign n7745 = Pg3229 & ~n7744;
  assign n7746 = ~Ng1267 & Ng1315;
  assign n7747 = ~Ng1268 & \[1605] ;
  assign n7748 = ~Ng1269 & \[1603] ;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = ~n7746 & n7749;
  assign n7751 = ~Ng1264 & Ng1315;
  assign n7752 = ~Ng1265 & \[1605] ;
  assign n7753 = ~Ng1266 & \[1603] ;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = ~n7751 & n7754;
  assign n7756 = n7750 & ~n7755;
  assign n7757 = ~Ng1261 & Ng1315;
  assign n7758 = ~Ng1262 & \[1605] ;
  assign n7759 = ~Ng1263 & \[1603] ;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~n7757 & n7760;
  assign n7762 = n7744 & ~n7761;
  assign n7763 = ~n7756 & n7762;
  assign n7764 = ~Pg3229 & n7756;
  assign n7765 = ~n7763 & ~n7764;
  assign n7766 = ~n7745 & n7765;
  assign n7767 = n7738 & ~n7766;
  assign n3427_1 = ~n7739 & ~n7767;
  assign n7769 = \[1603]  & n3566_1;
  assign n7770 = ~n7766 & n7769;
  assign n7771 = ~Ng1263 & ~n7769;
  assign n3432_1 = ~n7770 & ~n7771;
  assign n7773 = Ng1315 & n3566_1;
  assign n7774 = ~n7766 & n7773;
  assign n7775 = ~Ng1261 & ~n7773;
  assign n3437_1 = ~n7774 & ~n7775;
  assign n7777 = ~Pg3229 & ~n7761;
  assign n7778 = Pg3229 & n7761;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~n7750 & n7779;
  assign n7781 = ~n7756 & ~n7780;
  assign n7782 = n7738 & n7781;
  assign n7783 = Ng1265 & ~n7738;
  assign n3442_1 = n7782 | n7783;
  assign n7785 = n7769 & n7781;
  assign n7786 = Ng1266 & ~n7769;
  assign n3447_1 = n7785 | n7786;
  assign n7788 = n7773 & n7781;
  assign n7789 = Ng1264 & ~n7773;
  assign n3452_1 = n7788 | n7789;
  assign n7791 = n7744 & n7755;
  assign n7792 = n7779 & ~n7791;
  assign n7793 = n7755 & ~n7779;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = n7738 & ~n7794;
  assign n7796 = Ng1268 & ~n7738;
  assign n3457_1 = n7795 | n7796;
  assign n7798 = n7769 & ~n7794;
  assign n7799 = Ng1269 & ~n7769;
  assign n3462_1 = n7798 | n7799;
  assign n7801 = n7773 & ~n7794;
  assign n7802 = Ng1267 & ~n7773;
  assign n3467_1 = n7801 | n7802;
  assign n7804 = n7750 & n7755;
  assign n7805 = ~n7779 & n7804;
  assign n7806 = n7738 & ~n7805;
  assign n7807 = Ng1271 & ~n7738;
  assign n3472_1 = n7806 | n7807;
  assign n7809 = Ng1272 & ~n7769;
  assign n7810 = n7769 & ~n7805;
  assign n3477_1 = n7809 | n7810;
  assign n7812 = n7773 & ~n7805;
  assign n7813 = Ng1270 & ~n7773;
  assign n3482_1 = n7812 | n7813;
  assign n7815 = ~Ng1273 & ~\[1605] ;
  assign n7816 = Ng185 & Ng1210;
  assign n7817 = ~n3246_1 & n7816;
  assign n7818 = Ng1276 & \[1603] ;
  assign n7819 = Ng1279 & Ng1315;
  assign n7820 = Ng1273 & \[1605] ;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~n7818 & n7821;
  assign n7823 = ~n7817 & n7822;
  assign n7824 = ~n6032 & ~n7823;
  assign n7825 = \[1605]  & ~n7824;
  assign n3487_1 = ~n7815 & ~n7825;
  assign n7827 = ~Ng1276 & ~\[1603] ;
  assign n7828 = \[1603]  & ~n7824;
  assign n3492_1 = ~n7827 & ~n7828;
  assign n7830 = Ng1279 & ~Ng1315;
  assign n7831 = n6033 & ~n7823;
  assign n3497_1 = n7830 | n7831;
  assign n7833 = ~Ng1282 & ~\[1605] ;
  assign n7834 = Ng185 & Ng1228;
  assign n7835 = ~n3382_1 & n7834;
  assign n7836 = Ng1288 & Ng1315;
  assign n7837 = Ng1285 & \[1603] ;
  assign n7838 = Ng1282 & \[1605] ;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~n7836 & n7839;
  assign n7841 = ~n7835 & n7840;
  assign n7842 = ~n6032 & ~n7841;
  assign n7843 = \[1605]  & ~n7842;
  assign n3502_1 = ~n7833 & ~n7843;
  assign n7845 = ~Ng1285 & ~\[1603] ;
  assign n7846 = \[1603]  & ~n7842;
  assign n3507_1 = ~n7845 & ~n7846;
  assign n7848 = Ng1288 & ~Ng1315;
  assign n7849 = n6033 & ~n7841;
  assign n3512_1 = n7848 | n7849;
  assign n7851 = Ng1300 & ~\[1605] ;
  assign n7852 = ~n6032 & ~n7722;
  assign n7853 = ~n7823 & ~n7841;
  assign n7854 = n6032 & ~n7853;
  assign n7855 = Ng1040 & Ng1315;
  assign n7856 = Ng1036 & \[1605] ;
  assign n7857 = Ng1038 & \[1603] ;
  assign n7858 = ~n7856 & ~n7857;
  assign n7859 = ~n7855 & n7858;
  assign n7860 = Ng1055 & Ng1315;
  assign n7861 = Ng1051 & \[1605] ;
  assign n7862 = Ng1053 & \[1603] ;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = ~n7860 & n7863;
  assign n7865 = Ng1070 & Ng1315;
  assign n7866 = Ng1066 & \[1605] ;
  assign n7867 = Ng1068 & \[1603] ;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = ~n7865 & n7868;
  assign n7870 = ~n7864 & ~n7869;
  assign n7871 = ~n7744 & n7870;
  assign n7872 = ~n7750 & n7864;
  assign n7873 = n7791 & n7869;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = Ng1011 & Ng1315;
  assign n7876 = Ng1081 & \[1605] ;
  assign n7877 = Ng1083 & \[1603] ;
  assign n7878 = ~n7876 & ~n7877;
  assign n7879 = ~n7875 & n7878;
  assign n7880 = ~n7864 & ~n7879;
  assign n7881 = n7750 & n7880;
  assign n7882 = n7755 & n7881;
  assign n7883 = n7874 & ~n7882;
  assign n7884 = n7761 & ~n7883;
  assign n7885 = ~n7871 & ~n7884;
  assign n7886 = ~n7859 & ~n7885;
  assign n7887 = n7791 & n7870;
  assign n7888 = ~n7750 & n7880;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = n7859 & ~n7889;
  assign n7891 = ~n7755 & n7859;
  assign n7892 = n7869 & n7891;
  assign n7893 = n7804 & n7879;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n7890 & n7894;
  assign n7896 = ~n7761 & ~n7895;
  assign n7897 = n7761 & ~n7869;
  assign n7898 = n7750 & n7859;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = n7864 & ~n7899;
  assign n7901 = ~n7755 & n7900;
  assign n7902 = ~n7896 & ~n7901;
  assign n7903 = ~n7886 & n7902;
  assign n7904 = n7744 & ~n7859;
  assign n7905 = n7750 & ~n7904;
  assign n7906 = n7879 & ~n7905;
  assign n7907 = n7750 & ~n7859;
  assign n7908 = ~n7891 & ~n7907;
  assign n7909 = n7870 & n7908;
  assign n7910 = ~n7906 & ~n7909;
  assign n7911 = n7761 & ~n7910;
  assign n7912 = n7804 & ~n7864;
  assign n7913 = n7744 & ~n7912;
  assign n7914 = ~n7744 & ~n7879;
  assign n7915 = ~n7869 & ~n7914;
  assign n7916 = ~n7897 & ~n7915;
  assign n7917 = ~n7913 & n7916;
  assign n7918 = n7859 & n7917;
  assign n7919 = ~n7911 & ~n7918;
  assign n7920 = ~n7869 & ~n7905;
  assign n7921 = ~n7908 & ~n7920;
  assign n7922 = ~n7761 & n7864;
  assign n7923 = ~n7921 & n7922;
  assign n7924 = ~n7869 & ~n7881;
  assign n7925 = ~n7755 & ~n7872;
  assign n7926 = ~n7924 & n7925;
  assign n7927 = ~n7859 & n7926;
  assign n7928 = ~n7923 & ~n7927;
  assign n7929 = n7919 & n7928;
  assign n7930 = n7841 & n7929;
  assign n7931 = n7903 & ~n7930;
  assign n7932 = n7854 & n7931;
  assign n7933 = ~n7852 & ~n7932;
  assign n7934 = \[1605]  & ~n7933;
  assign n3517_1 = n7851 | n7934;
  assign n7936 = Ng1303 & ~\[1603] ;
  assign n7937 = \[1603]  & ~n7933;
  assign n3522_1 = n7936 | n7937;
  assign n7939 = Ng1306 & ~Ng1315;
  assign n7940 = Ng1315 & ~n7933;
  assign n3527_1 = n7939 | n7940;
  assign n7942 = Ng1291 & ~\[1605] ;
  assign n7943 = ~n6032 & ~n7734;
  assign n7944 = n7823 & n7903;
  assign n7945 = n7854 & n7929;
  assign n7946 = ~n7944 & n7945;
  assign n7947 = ~n7943 & ~n7946;
  assign n7948 = \[1605]  & ~n7947;
  assign n3532_1 = n7942 | n7948;
  assign n7950 = Ng1294 & ~\[1603] ;
  assign n7951 = \[1603]  & ~n7947;
  assign n3537_1 = n7950 | n7951;
  assign n7953 = Ng1297 & ~Ng1315;
  assign n7954 = Ng1315 & ~n7947;
  assign n3542_1 = n7953 | n7954;
  assign n7956 = ~Ng1177 & ~\[1605] ;
  assign n7957 = n7722 & n7728;
  assign n7958 = \[1605]  & ~n7957;
  assign n3547_1 = ~n7956 & ~n7958;
  assign n7960 = ~Ng1180 & ~\[1603] ;
  assign n7961 = \[1603]  & ~n7957;
  assign n3552_1 = ~n7960 & ~n7961;
  assign n7963 = ~Ng1183 & ~Ng1315;
  assign n7964 = Ng1315 & ~n7957;
  assign n3557_1 = ~n7963 & ~n7964;
  assign n7966 = Pg16355 & ~\[1603] ;
  assign n7967 = ~Ng1192 & ~n7966;
  assign n7968 = ~n6364_1 & n7967;
  assign n7969 = Ng1192 & ~Ng1193;
  assign n3571_1 = ~n7968 & ~n7969;
  assign n7971 = Pg3229 & Ng978;
  assign n7972 = ~Pg3229 & ~Ng992;
  assign n3619_1 = ~n7971 & ~n7972;
  assign n7974 = Ng1196 & Ng1315;
  assign n7975 = ~Ng1315 & Ng1316;
  assign n3642_1 = n7974 | n7975;
  assign n7977 = ~Ng1315 & ~Ng1345;
  assign n3647_1 = ~n6374_1 & ~n7977;
  assign n7979 = \[1603]  & Ng1316;
  assign n7980 = Ng1315 & ~Ng1345;
  assign n7981 = Ng1326 & n7980;
  assign n7982 = ~Ng1326 & ~n7980;
  assign n7983 = ~n7981 & ~n7982;
  assign n3652_1 = ~n7979 & n7983;
  assign n7985 = Ng1319 & n7981;
  assign n7986 = ~Ng1319 & ~n7981;
  assign n7987 = ~n7979 & ~n7986;
  assign n3657_1 = ~n7985 & n7987;
  assign n7989 = Ng1339 & n7985;
  assign n7990 = ~Ng1339 & ~n7985;
  assign n7991 = ~n7979 & ~n7990;
  assign n3662_1 = ~n7989 & n7991;
  assign n7993 = Ng1332 & n7989;
  assign n7994 = ~Ng1332 & ~n7989;
  assign n7995 = ~n7979 & ~n7994;
  assign n3667_1 = ~n7993 & n7995;
  assign n7997 = Ng1346 & n7993;
  assign n7998 = ~Ng1346 & ~n7993;
  assign n7999 = ~n7979 & ~n7998;
  assign n3672_1 = ~n7997 & n7999;
  assign n8001 = Ng1358 & n7997;
  assign n8002 = ~Ng1358 & ~n7997;
  assign n8003 = ~n7979 & ~n8002;
  assign n3677_1 = ~n8001 & n8003;
  assign n8005 = Ng1352 & n8001;
  assign n8006 = ~Ng1352 & ~n8001;
  assign n8007 = ~n7979 & ~n8006;
  assign n3682_1 = ~n8005 & n8007;
  assign n8009 = Ng1365 & n8005;
  assign n8010 = ~Ng1365 & ~n8005;
  assign n8011 = ~n7979 & ~n8010;
  assign n3687_1 = ~n8009 & n8011;
  assign n8013 = Ng1372 & n8009;
  assign n8014 = ~Ng1372 & ~n8009;
  assign n8015 = ~n7979 & ~n8014;
  assign n3692_1 = ~n8013 & n8015;
  assign n8017 = Ng1378 & n8013;
  assign n8018 = ~Ng1378 & ~n8013;
  assign n8019 = ~n8017 & ~n8018;
  assign n3697_1 = ~n7979 & n8019;
  assign n8021 = Ng1211 & ~Ng1345;
  assign n8022 = Ng1224 & n8021;
  assign n8023 = \[1605]  & n8022;
  assign n8024 = Ng1385 & ~n8023;
  assign n8025 = ~Ng1326 & n8023;
  assign n3702_1 = n8024 | n8025;
  assign n8027 = \[1603]  & n8022;
  assign n8028 = Ng1386 & ~n8027;
  assign n8029 = ~Ng1326 & n8027;
  assign n3707_1 = n8028 | n8029;
  assign n8031 = Ng1315 & n8022;
  assign n8032 = Ng1384 & ~n8031;
  assign n8033 = ~Ng1326 & n8031;
  assign n3712_1 = n8032 | n8033;
  assign n8035 = Ng1388 & ~n8023;
  assign n8036 = ~Ng1319 & n8023;
  assign n3717_1 = n8035 | n8036;
  assign n8038 = Ng1389 & ~n8027;
  assign n8039 = ~Ng1319 & n8027;
  assign n3722_1 = n8038 | n8039;
  assign n8041 = Ng1387 & ~n8031;
  assign n8042 = ~Ng1319 & n8031;
  assign n3727_1 = n8041 | n8042;
  assign n8044 = Ng1391 & ~n8023;
  assign n8045 = ~Ng1339 & n8023;
  assign n3732_1 = n8044 | n8045;
  assign n8047 = Ng1392 & ~n8027;
  assign n8048 = ~Ng1339 & n8027;
  assign n3737_1 = n8047 | n8048;
  assign n8050 = Ng1390 & ~n8031;
  assign n8051 = ~Ng1339 & n8031;
  assign n3742_1 = n8050 | n8051;
  assign n8053 = Ng1394 & ~n8023;
  assign n8054 = ~Ng1332 & n8023;
  assign n3747 = n8053 | n8054;
  assign n8056 = Ng1395 & ~n8027;
  assign n8057 = ~Ng1332 & n8027;
  assign n3752_1 = n8056 | n8057;
  assign n8059 = Ng1393 & ~n8031;
  assign n8060 = ~Ng1332 & n8031;
  assign n3757 = n8059 | n8060;
  assign n8062 = Ng1397 & ~n8023;
  assign n8063 = ~Ng1346 & n8023;
  assign n3762_1 = n8062 | n8063;
  assign n8065 = Ng1398 & ~n8027;
  assign n8066 = ~Ng1346 & n8027;
  assign n3767 = n8065 | n8066;
  assign n8068 = Ng1396 & ~n8031;
  assign n8069 = ~Ng1346 & n8031;
  assign n3772_1 = n8068 | n8069;
  assign n8071 = Ng1400 & ~n8023;
  assign n8072 = ~Ng1358 & n8023;
  assign n3777 = n8071 | n8072;
  assign n8074 = Ng1401 & ~n8027;
  assign n8075 = ~Ng1358 & n8027;
  assign n3782 = n8074 | n8075;
  assign n8077 = Ng1399 & ~n8031;
  assign n8078 = ~Ng1358 & n8031;
  assign n3787_1 = n8077 | n8078;
  assign n8080 = Ng1403 & ~n8023;
  assign n8081 = ~Ng1352 & n8023;
  assign n3792_1 = n8080 | n8081;
  assign n8083 = Ng1404 & ~n8027;
  assign n8084 = ~Ng1352 & n8027;
  assign n3797 = n8083 | n8084;
  assign n8086 = Ng1402 & ~n8031;
  assign n8087 = ~Ng1352 & n8031;
  assign n3802_1 = n8086 | n8087;
  assign n8089 = Ng1406 & ~n8023;
  assign n8090 = ~Ng1365 & n8023;
  assign n3807_1 = n8089 | n8090;
  assign n8092 = Ng1407 & ~n8027;
  assign n8093 = ~Ng1365 & n8027;
  assign n3812 = n8092 | n8093;
  assign n8095 = Ng1405 & ~n8031;
  assign n8096 = ~Ng1365 & n8031;
  assign n3817 = n8095 | n8096;
  assign n8098 = Ng1409 & ~n8023;
  assign n8099 = ~Ng1372 & n8023;
  assign n3822_1 = n8098 | n8099;
  assign n8101 = Ng1410 & ~n8027;
  assign n8102 = ~Ng1372 & n8027;
  assign n3827 = n8101 | n8102;
  assign n8104 = Ng1408 & ~n8031;
  assign n8105 = ~Ng1372 & n8031;
  assign n3832_1 = n8104 | n8105;
  assign n8107 = Ng1412 & ~n8023;
  assign n8108 = ~Ng1378 & n8023;
  assign n3837 = n8107 | n8108;
  assign n8110 = Ng1413 & ~n8027;
  assign n8111 = ~Ng1378 & n8027;
  assign n3842_1 = n8110 | n8111;
  assign n8113 = Ng1411 & ~n8031;
  assign n8114 = ~Ng1378 & n8031;
  assign n3847_1 = n8113 | n8114;
  assign n8116 = \[1605]  & Ng1316;
  assign n8117 = ~n7722 & n8116;
  assign n8118 = ~Ng1415 & ~n8116;
  assign n3852_1 = ~n8117 & ~n8118;
  assign n8120 = ~n7722 & n7979;
  assign n8121 = ~Ng1416 & ~n7979;
  assign n3857_1 = ~n8120 & ~n8121;
  assign n8123 = Ng1315 & Ng1316;
  assign n8124 = ~Ng1414 & ~n8123;
  assign n8125 = ~n7722 & n8123;
  assign n3862_1 = ~n8124 & ~n8125;
  assign n8127 = ~n7734 & n8116;
  assign n8128 = ~Ng1418 & ~n8116;
  assign n3867 = ~n8127 & ~n8128;
  assign n8130 = ~n7734 & n7979;
  assign n8131 = ~Ng1419 & ~n7979;
  assign n3872_1 = ~n8130 & ~n8131;
  assign n8133 = ~Ng1417 & ~n8123;
  assign n8134 = ~n7734 & n8123;
  assign n3877_1 = ~n8133 & ~n8134;
  assign n8136 = Ng1315 & ~Ng1387;
  assign n8137 = \[1605]  & ~Ng1388;
  assign n8138 = \[1603]  & ~Ng1389;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ~n8136 & n8139;
  assign n8141 = ~Ng1319 & ~n8140;
  assign n8142 = Ng1315 & ~Ng1402;
  assign n8143 = \[1605]  & ~Ng1403;
  assign n8144 = \[1603]  & ~Ng1404;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = ~n8142 & n8145;
  assign n8147 = Ng1352 & n8146;
  assign n8148 = ~n8141 & ~n8147;
  assign n8149 = Ng1315 & ~Ng1384;
  assign n8150 = \[1605]  & ~Ng1385;
  assign n8151 = \[1603]  & ~Ng1386;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = ~n8149 & n8152;
  assign n8154 = Ng1326 & n8153;
  assign n8155 = ~Ng1326 & ~n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = n8148 & n8156;
  assign n8158 = Ng1315 & ~Ng1393;
  assign n8159 = \[1605]  & ~Ng1394;
  assign n8160 = \[1603]  & ~Ng1395;
  assign n8161 = ~n8159 & ~n8160;
  assign n8162 = ~n8158 & n8161;
  assign n8163 = Ng1332 & n8162;
  assign n8164 = Ng1315 & ~Ng1396;
  assign n8165 = \[1605]  & ~Ng1397;
  assign n8166 = \[1603]  & ~Ng1398;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n8164 & n8167;
  assign n8169 = Ng1346 & n8168;
  assign n8170 = Ng1315 & ~Ng1390;
  assign n8171 = \[1605]  & ~Ng1391;
  assign n8172 = \[1603]  & ~Ng1392;
  assign n8173 = ~n8171 & ~n8172;
  assign n8174 = ~n8170 & n8173;
  assign n8175 = Ng1339 & n8174;
  assign n8176 = ~n8169 & ~n8175;
  assign n8177 = ~n8163 & n8176;
  assign n8178 = n8157 & n8177;
  assign n8179 = Ng1315 & ~Ng1399;
  assign n8180 = \[1605]  & ~Ng1400;
  assign n8181 = \[1603]  & ~Ng1401;
  assign n8182 = ~n8180 & ~n8181;
  assign n8183 = ~n8179 & n8182;
  assign n8184 = Ng1358 & ~n8183;
  assign n8185 = ~Ng1358 & n8183;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = n8178 & ~n8186;
  assign n8188 = ~Ng1339 & ~n8174;
  assign n8189 = Ng1319 & n8140;
  assign n8190 = ~Ng1352 & ~n8146;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = ~n8188 & n8191;
  assign n8193 = Ng1315 & ~Ng1405;
  assign n8194 = \[1605]  & ~Ng1406;
  assign n8195 = \[1603]  & ~Ng1407;
  assign n8196 = ~n8194 & ~n8195;
  assign n8197 = ~n8193 & n8196;
  assign n8198 = ~Ng1365 & n8197;
  assign n8199 = Ng1365 & ~n8197;
  assign n8200 = ~n8198 & ~n8199;
  assign n8201 = n8192 & ~n8200;
  assign n8202 = ~Ng1346 & ~n8168;
  assign n8203 = Ng1315 & ~Ng1411;
  assign n8204 = \[1605]  & ~Ng1412;
  assign n8205 = \[1603]  & ~Ng1413;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = ~n8203 & n8206;
  assign n8208 = ~Ng1378 & ~n8207;
  assign n8209 = ~Ng1332 & ~n8162;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8202 & n8210;
  assign n8212 = Ng1378 & n8207;
  assign n8213 = Ng1315 & ~Ng1408;
  assign n8214 = \[1605]  & ~Ng1409;
  assign n8215 = \[1603]  & ~Ng1410;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = ~n8213 & n8216;
  assign n8218 = ~Ng1372 & n8217;
  assign n8219 = Ng1372 & ~n8217;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = ~n8212 & ~n8220;
  assign n8222 = n8211 & n8221;
  assign n8223 = n8201 & n8222;
  assign n8224 = n8187 & n8223;
  assign n8225 = Ng1315 & ~Ng1414;
  assign n8226 = Ng1315 & ~Ng1417;
  assign n8227 = \[1605]  & ~Ng1418;
  assign n8228 = \[1603]  & ~Ng1419;
  assign n8229 = ~n8227 & ~n8228;
  assign n8230 = ~n8226 & n8229;
  assign n8231 = \[1605]  & ~Ng1415;
  assign n8232 = \[1603]  & ~Ng1416;
  assign n8233 = ~n8231 & ~n8232;
  assign n8234 = n8230 & n8233;
  assign n8235 = ~n8225 & n8234;
  assign n8236 = ~n8224 & n8235;
  assign n8237 = n8023 & n8236;
  assign n8238 = Ng1421 & ~n8023;
  assign n3882 = n8237 | n8238;
  assign n8240 = n8027 & n8236;
  assign n8241 = Ng1422 & ~n8027;
  assign n3887 = n8240 | n8241;
  assign n8243 = n8031 & n8236;
  assign n8244 = Ng1420 & ~n8031;
  assign n3892_1 = n8243 | n8244;
  assign n8246 = ~Ng1424 & ~n8023;
  assign n3897_1 = ~n8116 & ~n8246;
  assign n8248 = ~Ng1425 & ~n8027;
  assign n3902 = ~n7979 & ~n8248;
  assign n8250 = ~Ng1423 & ~n8031;
  assign n3907_1 = ~n8123 & ~n8250;
  assign n8252 = Ng1512 & ~n5019_1;
  assign n8253 = ~Ng1471 & n5019_1;
  assign n3912_1 = n8252 | n8253;
  assign n8255 = Ng1513 & ~n5023;
  assign n8256 = ~Ng1471 & n5023;
  assign n3917 = n8255 | n8256;
  assign n8258 = Ng1511 & ~n5027;
  assign n8259 = ~Ng1471 & n5027;
  assign n3922 = n8258 | n8259;
  assign n8261 = Ng1515 & ~n5019_1;
  assign n8262 = ~Ng1476 & n5019_1;
  assign n3927 = n8261 | n8262;
  assign n8264 = Ng1516 & ~n5023;
  assign n8265 = ~Ng1476 & n5023;
  assign n3932_1 = n8264 | n8265;
  assign n8267 = Ng1514 & ~n5027;
  assign n8268 = ~Ng1476 & n5027;
  assign n3937 = n8267 | n8268;
  assign n8270 = Ng1524 & ~n5019_1;
  assign n8271 = ~Ng1481 & n5019_1;
  assign n3942_1 = n8270 | n8271;
  assign n8273 = Ng1525 & ~n5023;
  assign n8274 = ~Ng1481 & n5023;
  assign n3947 = n8273 | n8274;
  assign n8276 = Ng1523 & ~n5027;
  assign n8277 = ~Ng1481 & n5027;
  assign n3952 = n8276 | n8277;
  assign n8279 = Ng1527 & ~n5019_1;
  assign n8280 = ~Ng1486 & n5019_1;
  assign n3957_1 = n8279 | n8280;
  assign n8282 = Ng1528 & ~n5023;
  assign n8283 = ~Ng1486 & n5023;
  assign n3962 = n8282 | n8283;
  assign n8285 = Ng1526 & ~n5027;
  assign n8286 = ~Ng1486 & n5027;
  assign n3967 = n8285 | n8286;
  assign n8288 = Ng1530 & ~n5019_1;
  assign n8289 = ~Ng1491 & n5019_1;
  assign n3972 = n8288 | n8289;
  assign n8291 = Ng1531 & ~n5023;
  assign n8292 = ~Ng1491 & n5023;
  assign n3977 = n8291 | n8292;
  assign n8294 = Ng1529 & ~n5027;
  assign n8295 = ~Ng1491 & n5027;
  assign n3982 = n8294 | n8295;
  assign n8297 = Ng1533 & ~n5019_1;
  assign n8298 = ~Ng1496 & n5019_1;
  assign n3987 = n8297 | n8298;
  assign n8300 = Ng1534 & ~n5023;
  assign n8301 = ~Ng1496 & n5023;
  assign n3992 = n8300 | n8301;
  assign n8303 = Ng1532 & ~n5027;
  assign n8304 = ~Ng1496 & n5027;
  assign n3997_1 = n8303 | n8304;
  assign n8306 = Ng1536 & ~n5019_1;
  assign n8307 = ~Ng1501 & n5019_1;
  assign n4002_1 = n8306 | n8307;
  assign n8309 = Ng1537 & ~n5023;
  assign n8310 = ~Ng1501 & n5023;
  assign n4007_1 = n8309 | n8310;
  assign n8312 = Ng1535 & ~n5027;
  assign n8313 = ~Ng1501 & n5027;
  assign n4012 = n8312 | n8313;
  assign n8315 = Ng1539 & ~n5019_1;
  assign n8316 = ~Ng1506 & n5019_1;
  assign n4017 = n8315 | n8316;
  assign n8318 = Ng1540 & ~n5023;
  assign n8319 = ~Ng1506 & n5023;
  assign n4022_1 = n8318 | n8319;
  assign n8321 = Ng1538 & ~n5027;
  assign n8322 = ~Ng1506 & n5027;
  assign n4027 = n8321 | n8322;
  assign n8324 = ~Ng1542 & ~n5019_1;
  assign n8325 = Ng853 & ~Ng1556;
  assign n8326 = \[1612]  & ~Ng1557;
  assign n8327 = \[1594]  & ~Ng1558;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = ~n8325 & n8328;
  assign n8330 = n5019_1 & ~n8329;
  assign n4032_1 = ~n8324 & ~n8330;
  assign n8332 = n5023 & n8329;
  assign n8333 = Ng1543 & ~n5023;
  assign n4037_1 = n8332 | n8333;
  assign n8335 = ~Ng1541 & ~n5027;
  assign n8336 = n5027 & ~n8329;
  assign n4042 = ~n8335 & ~n8336;
  assign n8338 = ~Ng1545 & ~n5019_1;
  assign n8339 = Ng853 & ~Ng1553;
  assign n8340 = \[1612]  & ~Ng1554;
  assign n8341 = \[1594]  & ~Ng1555;
  assign n8342 = ~n8340 & ~n8341;
  assign n8343 = ~n8339 & n8342;
  assign n8344 = n5019_1 & ~n8343;
  assign n4047 = ~n8338 & ~n8344;
  assign n8346 = n5023 & n8343;
  assign n8347 = Ng1546 & ~n5023;
  assign n4052 = n8346 | n8347;
  assign n8349 = ~Ng1544 & ~n5027;
  assign n8350 = n5027 & ~n8343;
  assign n4057_1 = ~n8349 & ~n8350;
  assign n8352 = Ng1506 & Ng1491;
  assign n8353 = ~Ng1496 & n8352;
  assign n8354 = ~Ng1501 & n8353;
  assign n8355 = n5131_1 & n8354;
  assign n8356 = Ng1551 & ~n5131_1;
  assign n4062_1 = n8355 | n8356;
  assign n8358 = n5138 & n8354;
  assign n8359 = Ng1552 & ~n5138;
  assign n4067 = n8358 | n8359;
  assign n8361 = n5142 & n8354;
  assign n8362 = Ng1550 & ~n5142;
  assign n4072_1 = n8361 | n8362;
  assign n8364 = Ng1554 & ~n5131_1;
  assign n8365 = ~Ng1476 & n5131_1;
  assign n4077 = n8364 | n8365;
  assign n8367 = Ng1555 & ~n5138;
  assign n8368 = ~Ng1476 & n5138;
  assign n4082 = n8367 | n8368;
  assign n8370 = Ng1553 & ~n5142;
  assign n8371 = ~Ng1476 & n5142;
  assign n4087 = n8370 | n8371;
  assign n8373 = Ng1557 & ~n5131_1;
  assign n8374 = ~Ng1471 & n5131_1;
  assign n4092 = n8373 | n8374;
  assign n8376 = Ng1558 & ~n5138;
  assign n8377 = ~Ng1471 & n5138;
  assign n4097 = n8376 | n8377;
  assign n8379 = Ng1556 & ~n5142;
  assign n8380 = ~Ng1471 & n5142;
  assign n4102_1 = n8379 | n8380;
  assign n8382 = Ng1560 & ~n5131_1;
  assign n8383 = Ng1476 & Ng1471;
  assign n8384 = Ng1486 & Ng1481;
  assign n8385 = n8383 & n8384;
  assign n8386 = Ng1501 & Ng1496;
  assign n8387 = n8352 & n8386;
  assign n8388 = n8385 & n8387;
  assign n8389 = n5131_1 & ~n8388;
  assign n4107_1 = n8382 | n8389;
  assign n8391 = Ng1561 & ~n5138;
  assign n8392 = n5138 & ~n8388;
  assign n4112_1 = n8391 | n8392;
  assign n8394 = Ng1559 & ~n5142;
  assign n8395 = n5142 & ~n8388;
  assign n4117 = n8394 | n8395;
  assign n8397 = ~\[1612]  & ~Ng1567;
  assign n8398 = Ng853 & Ng1573;
  assign n8399 = \[1612]  & Ng1567;
  assign n8400 = \[1594]  & Ng1570;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = ~n8398 & n8401;
  assign n8403 = Ng853 & ~Ng1701;
  assign n8404 = \[1612]  & ~Ng1699;
  assign n8405 = \[1594]  & ~Ng1700;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = ~n8403 & n8406;
  assign n8408 = Ng853 & ~Ng1695;
  assign n8409 = \[1612]  & ~Ng1693;
  assign n8410 = \[1594]  & ~Ng1694;
  assign n8411 = ~n8409 & ~n8410;
  assign n8412 = ~n8408 & n8411;
  assign n8413 = n8407 & n8412;
  assign n8414 = n8402 & n8413;
  assign n8415 = Ng853 & Ng1645;
  assign n8416 = \[1612]  & Ng1639;
  assign n8417 = \[1594]  & Ng1642;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = ~n8415 & n8418;
  assign n8420 = Ng853 & Ng1600;
  assign n8421 = \[1612]  & Ng1594;
  assign n8422 = \[1594]  & Ng1597;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n8420 & n8423;
  assign n8425 = n8419 & n8424;
  assign n8426 = Ng853 & Ng1636;
  assign n8427 = \[1612]  & Ng1630;
  assign n8428 = \[1594]  & Ng1633;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~n8426 & n8429;
  assign n8431 = Ng853 & Ng1591;
  assign n8432 = \[1612]  & Ng1585;
  assign n8433 = \[1594]  & Ng1588;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = ~n8431 & n8434;
  assign n8436 = n8430 & n8435;
  assign n8437 = n8425 & n8436;
  assign n8438 = n8414 & n8437;
  assign n8439 = Ng853 & ~Ng1698;
  assign n8440 = \[1612]  & ~Ng1696;
  assign n8441 = \[1594]  & ~Ng1697;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = ~n8439 & n8442;
  assign n8444 = Ng853 & Ng1582;
  assign n8445 = \[1612]  & Ng1576;
  assign n8446 = \[1594]  & Ng1579;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = ~n8444 & n8447;
  assign n8449 = n8443 & n8448;
  assign n8450 = Ng853 & Ng1654;
  assign n8451 = \[1612]  & Ng1648;
  assign n8452 = \[1594]  & Ng1651;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = ~n8450 & n8453;
  assign n8455 = Ng853 & Ng1627;
  assign n8456 = \[1612]  & Ng1621;
  assign n8457 = \[1594]  & Ng1624;
  assign n8458 = ~n8456 & ~n8457;
  assign n8459 = ~n8455 & n8458;
  assign n8460 = n8454 & n8459;
  assign n8461 = n8449 & n8460;
  assign n8462 = Ng853 & Ng1618;
  assign n8463 = \[1612]  & Ng1612;
  assign n8464 = \[1594]  & Ng1615;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = ~n8462 & n8465;
  assign n8467 = Ng853 & Ng1609;
  assign n8468 = \[1612]  & Ng1603;
  assign n8469 = \[1594]  & Ng1606;
  assign n8470 = ~n8468 & ~n8469;
  assign n8471 = ~n8467 & n8470;
  assign n8472 = n8466 & n8471;
  assign n8473 = n8461 & n8472;
  assign n8474 = n8438 & n8473;
  assign n8475 = ~n8412 & n8443;
  assign n8476 = ~n8407 & n8475;
  assign n8477 = n8407 & ~n8412;
  assign n8478 = Ng853 & ~Ng1550;
  assign n8479 = \[1612]  & ~Ng1551;
  assign n8480 = \[1594]  & ~Ng1552;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n8478 & n8481;
  assign n8483 = Ng2257 & ~n8482;
  assign n8484 = ~Ng1506 & ~n8419;
  assign n8485 = Ng1506 & n8419;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = ~Ng1476 & ~n8466;
  assign n8488 = Ng1476 & n8466;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = n8486 & n8489;
  assign n8491 = ~Ng1486 & ~n8459;
  assign n8492 = Ng1486 & n8459;
  assign n8493 = ~n8491 & ~n8492;
  assign n8494 = ~n8343 & ~n8454;
  assign n8495 = n8343 & n8454;
  assign n8496 = ~n8494 & ~n8495;
  assign n8497 = n8493 & ~n8496;
  assign n8498 = ~Ng1496 & ~n8430;
  assign n8499 = Ng1496 & n8430;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~n8497 & ~n8500;
  assign n8502 = n8486 & ~n8496;
  assign n8503 = ~n8489 & ~n8502;
  assign n8504 = ~n8501 & ~n8503;
  assign n8505 = n8493 & n8500;
  assign n8506 = ~n8504 & ~n8505;
  assign n8507 = ~n8490 & n8506;
  assign n8508 = n8486 & n8500;
  assign n8509 = n8489 & n8493;
  assign n8510 = n8496 & ~n8509;
  assign n8511 = ~n8508 & n8510;
  assign n8512 = ~n8507 & ~n8511;
  assign n8513 = n8483 & ~n8512;
  assign n8514 = ~Ng1471 & ~n8402;
  assign n8515 = Ng1471 & n8402;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = ~Ng1481 & ~n8448;
  assign n8518 = Ng1481 & n8448;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = n8516 & n8519;
  assign n8521 = ~Ng1491 & ~n8435;
  assign n8522 = Ng1491 & n8435;
  assign n8523 = ~n8521 & ~n8522;
  assign n8524 = ~Ng1501 & ~n8424;
  assign n8525 = Ng1501 & n8424;
  assign n8526 = ~n8524 & ~n8525;
  assign n8527 = n8523 & n8526;
  assign n8528 = ~n8520 & ~n8527;
  assign n8529 = ~n8523 & ~n8526;
  assign n8530 = ~n8516 & ~n8519;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = n8329 & ~n8471;
  assign n8533 = ~n8329 & n8471;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = ~n8531 & ~n8534;
  assign n8536 = ~n8528 & ~n8535;
  assign n8537 = n8531 & n8534;
  assign n8538 = n8483 & ~n8537;
  assign n8539 = ~n8536 & n8538;
  assign n8540 = ~n8513 & ~n8539;
  assign n8541 = n8477 & n8540;
  assign n8542 = ~n8476 & ~n8541;
  assign n8543 = Ng853 & ~Ng1514;
  assign n8544 = \[1612]  & ~Ng1515;
  assign n8545 = \[1594]  & ~Ng1516;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = ~n8543 & n8546;
  assign n8548 = Ng1476 & n8547;
  assign n8549 = n8483 & ~n8548;
  assign n8550 = Ng853 & ~Ng1538;
  assign n8551 = \[1612]  & ~Ng1539;
  assign n8552 = \[1594]  & ~Ng1540;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 = ~n8550 & n8553;
  assign n8555 = Ng1506 & n8554;
  assign n8556 = ~Ng1506 & ~n8554;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = n8549 & n8557;
  assign n8559 = Ng853 & ~Ng1511;
  assign n8560 = \[1612]  & ~Ng1512;
  assign n8561 = \[1594]  & ~Ng1513;
  assign n8562 = ~n8560 & ~n8561;
  assign n8563 = ~n8559 & n8562;
  assign n8564 = Ng1471 & n8563;
  assign n8565 = Ng853 & ~Ng1544;
  assign n8566 = \[1612]  & ~Ng1545;
  assign n8567 = \[1594]  & ~Ng1546;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = ~n8565 & n8568;
  assign n8570 = ~n8343 & n8569;
  assign n8571 = ~n8564 & ~n8570;
  assign n8572 = Ng853 & ~Ng1526;
  assign n8573 = \[1594]  & ~Ng1528;
  assign n8574 = \[1612]  & ~Ng1527;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = ~n8572 & n8575;
  assign n8577 = ~Ng1486 & n8576;
  assign n8578 = Ng1486 & ~n8576;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = n8571 & ~n8579;
  assign n8581 = n8558 & n8580;
  assign n8582 = n8343 & ~n8569;
  assign n8583 = ~Ng1471 & ~n8563;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8581 & n8584;
  assign n8586 = Ng853 & ~Ng1541;
  assign n8587 = \[1612]  & ~Ng1542;
  assign n8588 = \[1594]  & ~Ng1543;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = ~n8586 & n8589;
  assign n8591 = ~n8329 & n8590;
  assign n8592 = Ng853 & ~Ng1535;
  assign n8593 = \[1612]  & ~Ng1536;
  assign n8594 = \[1594]  & ~Ng1537;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = ~n8592 & n8595;
  assign n8597 = ~Ng1501 & n8596;
  assign n8598 = Ng1501 & ~n8596;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8591 & ~n8599;
  assign n8601 = Ng853 & ~Ng1523;
  assign n8602 = \[1594]  & ~Ng1525;
  assign n8603 = \[1612]  & ~Ng1524;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8601 & n8604;
  assign n8606 = Ng1481 & n8605;
  assign n8607 = n8600 & ~n8606;
  assign n8608 = Ng853 & ~Ng1532;
  assign n8609 = \[1612]  & ~Ng1533;
  assign n8610 = \[1594]  & ~Ng1534;
  assign n8611 = ~n8609 & ~n8610;
  assign n8612 = ~n8608 & n8611;
  assign n8613 = ~Ng1496 & n8612;
  assign n8614 = Ng1496 & ~n8612;
  assign n8615 = ~n8613 & ~n8614;
  assign n8616 = Ng853 & ~Ng1529;
  assign n8617 = \[1612]  & ~Ng1530;
  assign n8618 = \[1594]  & ~Ng1531;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = ~n8616 & n8619;
  assign n8621 = ~Ng1491 & ~n8620;
  assign n8622 = ~Ng1481 & ~n8605;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8615 & n8623;
  assign n8625 = Ng1491 & n8620;
  assign n8626 = ~Ng1476 & ~n8547;
  assign n8627 = n8329 & ~n8590;
  assign n8628 = ~n8626 & ~n8627;
  assign n8629 = ~n8625 & n8628;
  assign n8630 = n8624 & n8629;
  assign n8631 = n8607 & n8630;
  assign n8632 = n8585 & n8631;
  assign n8633 = \[1594]  & ~Ng1704;
  assign n8634 = Ng853 & ~Ng1702;
  assign n8635 = \[1612]  & ~Ng1703;
  assign n8636 = ~n8634 & ~n8635;
  assign n8637 = ~n8633 & n8636;
  assign n8638 = n8632 & ~n8637;
  assign n8639 = n8443 & n8638;
  assign n8640 = ~n8542 & n8639;
  assign n8641 = Ng2257 & n8482;
  assign n8642 = ~n8412 & n8641;
  assign n8643 = Ng853 & ~Ng1783;
  assign n8644 = \[1612]  & ~Ng1784;
  assign n8645 = \[1594]  & ~Ng1785;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n8643 & n8646;
  assign n8648 = n8632 & ~n8647;
  assign n8649 = ~n8642 & ~n8648;
  assign n8650 = ~n8640 & n8649;
  assign n8651 = ~n8454 & ~n8466;
  assign n8652 = ~n8448 & n8651;
  assign n8653 = n8413 & ~n8443;
  assign n8654 = ~n8471 & n8653;
  assign n8655 = n8402 & n8437;
  assign n8656 = n8654 & n8655;
  assign n8657 = n8652 & n8656;
  assign n8658 = ~n8459 & n8657;
  assign n8659 = n8650 & ~n8658;
  assign n8660 = ~n8474 & n8659;
  assign n8661 = Ng1471 & ~n8650;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = ~n8402 & ~n8413;
  assign n8664 = ~n8414 & ~n8663;
  assign n8665 = n8659 & n8664;
  assign n8666 = ~n8662 & ~n8665;
  assign n8667 = \[1612]  & ~n8666;
  assign n4122_1 = ~n8397 & ~n8667;
  assign n8669 = ~\[1594]  & ~Ng1570;
  assign n8670 = \[1594]  & ~n8666;
  assign n4127_1 = ~n8669 & ~n8670;
  assign n8672 = ~Ng853 & ~Ng1573;
  assign n8673 = Ng853 & ~n8666;
  assign n4132_1 = ~n8672 & ~n8673;
  assign n8675 = ~\[1612]  & ~Ng1612;
  assign n8676 = Ng1476 & ~n8650;
  assign n8677 = ~n8659 & ~n8676;
  assign n8678 = n8402 & n8443;
  assign n8679 = ~n8402 & ~n8443;
  assign n8680 = ~n8678 & ~n8679;
  assign n8681 = n8413 & ~n8680;
  assign n8682 = ~n8466 & n8681;
  assign n8683 = n8466 & ~n8681;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = n8660 & ~n8684;
  assign n8686 = ~n8677 & ~n8685;
  assign n8687 = \[1612]  & ~n8686;
  assign n4137_1 = ~n8675 & ~n8687;
  assign n8689 = ~\[1594]  & ~Ng1615;
  assign n8690 = \[1594]  & ~n8686;
  assign n4142_1 = ~n8689 & ~n8690;
  assign n8692 = ~Ng853 & ~Ng1618;
  assign n8693 = Ng853 & ~n8686;
  assign n4147_1 = ~n8692 & ~n8693;
  assign n8695 = ~\[1612]  & ~Ng1576;
  assign n8696 = Ng1481 & ~n8650;
  assign n8697 = ~n8659 & ~n8696;
  assign n8698 = ~n8466 & n8679;
  assign n8699 = n8466 & n8678;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = n8413 & ~n8700;
  assign n8702 = n8448 & n8701;
  assign n8703 = ~n8448 & ~n8701;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8660 & n8704;
  assign n8706 = ~n8697 & ~n8705;
  assign n8707 = \[1612]  & ~n8706;
  assign n4152 = ~n8695 & ~n8707;
  assign n8709 = ~\[1594]  & ~Ng1579;
  assign n8710 = \[1594]  & ~n8706;
  assign n4157 = ~n8709 & ~n8710;
  assign n8712 = ~Ng853 & ~Ng1582;
  assign n8713 = Ng853 & ~n8706;
  assign n4162 = ~n8712 & ~n8713;
  assign n8715 = ~\[1612]  & ~Ng1621;
  assign n8716 = Ng1486 & ~n8650;
  assign n8717 = ~n8659 & ~n8716;
  assign n8718 = ~n8443 & ~n8448;
  assign n8719 = ~n8449 & ~n8718;
  assign n8720 = n8701 & ~n8719;
  assign n8721 = ~n8459 & n8720;
  assign n8722 = n8459 & ~n8720;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = n8660 & ~n8723;
  assign n8725 = ~n8717 & ~n8724;
  assign n8726 = \[1612]  & ~n8725;
  assign n4167_1 = ~n8715 & ~n8726;
  assign n8728 = ~\[1594]  & ~Ng1624;
  assign n8729 = \[1594]  & ~n8725;
  assign n4172 = ~n8728 & ~n8729;
  assign n8731 = ~Ng853 & ~Ng1627;
  assign n8732 = Ng853 & ~n8725;
  assign n4177 = ~n8731 & ~n8732;
  assign n8734 = Ng1491 & ~n8650;
  assign n8735 = ~n8459 & ~n8653;
  assign n8736 = n8459 & n8653;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = n8720 & n8737;
  assign n8739 = ~n8435 & n8738;
  assign n8740 = n8435 & ~n8738;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = n8660 & n8741;
  assign n8743 = ~n8734 & ~n8742;
  assign n8744 = \[1612]  & n8743;
  assign n8745 = ~\[1612]  & ~Ng1585;
  assign n4182 = ~n8744 & ~n8745;
  assign n8747 = \[1594]  & n8743;
  assign n8748 = ~\[1594]  & ~Ng1588;
  assign n4187_1 = ~n8747 & ~n8748;
  assign n8750 = Ng853 & n8743;
  assign n8751 = ~Ng853 & ~Ng1591;
  assign n4192 = ~n8750 & ~n8751;
  assign n8753 = ~\[1612]  & Ng1630;
  assign n8754 = Ng1496 & ~n8650;
  assign n8755 = ~n8435 & n8653;
  assign n8756 = n8435 & ~n8653;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = n8738 & ~n8757;
  assign n8759 = n8430 & n8758;
  assign n8760 = ~n8430 & ~n8758;
  assign n8761 = ~n8759 & ~n8760;
  assign n8762 = n8660 & ~n8761;
  assign n8763 = ~n8754 & ~n8762;
  assign n8764 = \[1612]  & ~n8763;
  assign n4197_1 = n8753 | n8764;
  assign n8766 = ~\[1594]  & Ng1633;
  assign n8767 = \[1594]  & ~n8763;
  assign n4202 = n8766 | n8767;
  assign n8769 = ~Ng853 & Ng1636;
  assign n8770 = Ng853 & ~n8763;
  assign n4207 = n8769 | n8770;
  assign n8772 = Ng1501 & ~n8650;
  assign n8773 = n8430 & n8653;
  assign n8774 = n8721 & n8755;
  assign n8775 = ~n8759 & ~n8774;
  assign n8776 = ~n8773 & ~n8775;
  assign n8777 = n8424 & n8776;
  assign n8778 = ~n8424 & ~n8776;
  assign n8779 = ~n8777 & ~n8778;
  assign n8780 = n8660 & ~n8779;
  assign n8781 = ~n8772 & ~n8780;
  assign n8782 = \[1612]  & n8781;
  assign n8783 = ~\[1612]  & ~Ng1594;
  assign n4212_1 = ~n8782 & ~n8783;
  assign n8785 = \[1594]  & n8781;
  assign n8786 = ~\[1594]  & ~Ng1597;
  assign n4217_1 = ~n8785 & ~n8786;
  assign n8788 = Ng853 & n8781;
  assign n8789 = ~Ng853 & ~Ng1600;
  assign n4222 = ~n8788 & ~n8789;
  assign n8791 = Ng1506 & ~n8650;
  assign n8792 = ~n8424 & n8653;
  assign n8793 = n8424 & ~n8653;
  assign n8794 = ~n8792 & ~n8793;
  assign n8795 = n8776 & ~n8794;
  assign n8796 = n8419 & n8795;
  assign n8797 = ~n8419 & ~n8795;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = n8660 & ~n8798;
  assign n8800 = ~n8791 & ~n8799;
  assign n8801 = \[1612]  & n8800;
  assign n8802 = ~\[1612]  & ~Ng1639;
  assign n4227 = ~n8801 & ~n8802;
  assign n8804 = \[1594]  & n8800;
  assign n8805 = ~\[1594]  & ~Ng1642;
  assign n4232 = ~n8804 & ~n8805;
  assign n8807 = Ng853 & n8800;
  assign n8808 = ~Ng853 & ~Ng1645;
  assign n4237 = ~n8807 & ~n8808;
  assign n8810 = ~\[1612]  & ~Ng1603;
  assign n8811 = ~n8329 & ~n8650;
  assign n8812 = ~n8659 & ~n8811;
  assign n8813 = ~n8419 & ~n8430;
  assign n8814 = ~n8425 & ~n8813;
  assign n8815 = ~n8794 & ~n8814;
  assign n8816 = ~n8775 & n8815;
  assign n8817 = ~n8471 & n8816;
  assign n8818 = n8471 & ~n8816;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = n8660 & ~n8819;
  assign n8821 = ~n8812 & ~n8820;
  assign n8822 = \[1612]  & ~n8821;
  assign n4242 = ~n8810 & ~n8822;
  assign n8824 = ~\[1594]  & ~Ng1606;
  assign n8825 = \[1594]  & ~n8821;
  assign n4247 = ~n8824 & ~n8825;
  assign n8827 = ~Ng853 & ~Ng1609;
  assign n8828 = Ng853 & ~n8821;
  assign n4252_1 = ~n8827 & ~n8828;
  assign n8830 = ~\[1612]  & ~Ng1648;
  assign n8831 = ~n8343 & ~n8650;
  assign n8832 = ~n8659 & ~n8831;
  assign n8833 = n8471 & ~n8653;
  assign n8834 = ~n8654 & ~n8833;
  assign n8835 = n8816 & ~n8834;
  assign n8836 = ~n8454 & n8835;
  assign n8837 = n8454 & ~n8835;
  assign n8838 = ~n8836 & ~n8837;
  assign n8839 = n8660 & ~n8838;
  assign n8840 = ~n8832 & ~n8839;
  assign n8841 = \[1612]  & ~n8840;
  assign n4257_1 = ~n8830 & ~n8841;
  assign n8843 = ~\[1594]  & ~Ng1651;
  assign n8844 = \[1594]  & ~n8840;
  assign n4262 = ~n8843 & ~n8844;
  assign n8846 = ~Ng853 & ~Ng1654;
  assign n8847 = Ng853 & ~n8840;
  assign n4267 = ~n8846 & ~n8847;
  assign n8849 = Ng1466 & n5635;
  assign n8850 = Ng1466 & ~n5027;
  assign n8851 = ~n5635 & ~n8850;
  assign n4272 = ~n8849 & ~n8851;
  assign n8853 = Ng1462 & n8849;
  assign n8854 = ~Ng1462 & ~n8849;
  assign n8855 = ~n5642 & ~n8854;
  assign n4277 = ~n8853 & n8855;
  assign n8857 = Ng1457 & n8853;
  assign n8858 = ~Ng1457 & ~n8853;
  assign n8859 = ~n5642 & ~n8858;
  assign n4282 = ~n8857 & n8859;
  assign n8861 = Ng1453 & n8857;
  assign n8862 = ~Ng1453 & ~n8857;
  assign n8863 = ~n5642 & ~n8862;
  assign n4287 = ~n8861 & n8863;
  assign n8865 = Ng1448 & n8861;
  assign n8866 = ~Ng1448 & ~n8861;
  assign n8867 = ~n5642 & ~n8866;
  assign n4292 = ~n8865 & n8867;
  assign n8869 = Ng1444 & n8865;
  assign n8870 = ~Ng1444 & ~n8865;
  assign n8871 = ~n5642 & ~n8870;
  assign n4297 = ~n8869 & n8871;
  assign n8873 = Ng1439 & n8869;
  assign n8874 = ~Ng1439 & ~n8869;
  assign n8875 = ~n5642 & ~n8874;
  assign n4302 = ~n8873 & n8875;
  assign n8877 = Ng1435 & n8873;
  assign n8878 = ~Ng1435 & ~n8873;
  assign n8879 = ~n5642 & ~n8878;
  assign n4307 = ~n8877 & n8879;
  assign n8881 = Ng1430 & n8877;
  assign n8882 = ~Ng1430 & ~n8877;
  assign n8883 = ~n5642 & ~n8882;
  assign n4312 = ~n8881 & n8883;
  assign n8885 = Ng1426 & n8881;
  assign n8886 = ~Ng1426 & ~n8881;
  assign n8887 = ~n8885 & ~n8886;
  assign n4317 = ~n5642 & n8887;
  assign n8889 = n8413 & n8443;
  assign n8890 = n8412 & ~n8443;
  assign n8891 = ~n8407 & n8890;
  assign n8892 = ~n5124 & ~n8891;
  assign n8893 = ~n8889 & ~n8892;
  assign n8894 = \[1612]  & ~n8893;
  assign n8895 = Ng853 & ~Ng11553;
  assign n8896 = \[1612]  & ~Ng11551;
  assign n8897 = \[1594]  & ~Ng11552;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = ~n8895 & n8898;
  assign n8900 = Ng853 & ~Ng11559;
  assign n8901 = \[1612]  & ~Ng11557;
  assign n8902 = \[1594]  & ~Ng11558;
  assign n8903 = ~n8901 & ~n8902;
  assign n8904 = ~n8900 & n8903;
  assign n8905 = Ng853 & ~Ng11556;
  assign n8906 = \[1612]  & ~Ng11554;
  assign n8907 = \[1594]  & ~Ng11555;
  assign n8908 = ~n8906 & ~n8907;
  assign n8909 = ~n8905 & n8908;
  assign n8910 = n8904 & ~n8909;
  assign n8911 = Ng853 & ~Ng11562;
  assign n8912 = \[1612]  & ~Ng11560;
  assign n8913 = \[1594]  & ~Ng11561;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = ~n8911 & n8914;
  assign n8916 = ~n8910 & n8915;
  assign n8917 = ~n8899 & n8916;
  assign n8918 = ~Pg3229 & n8910;
  assign n8919 = Pg3229 & ~n8915;
  assign n8920 = ~n8918 & ~n8919;
  assign n8921 = ~n8917 & n8920;
  assign n8922 = n8894 & ~n8921;
  assign n8923 = ~Ng11551 & ~n8894;
  assign n4322_1 = ~n8922 & ~n8923;
  assign n8925 = \[1594]  & ~n8893;
  assign n8926 = ~n8921 & n8925;
  assign n8927 = ~Ng11552 & ~n8925;
  assign n4327 = ~n8926 & ~n8927;
  assign n8929 = Ng853 & ~n8893;
  assign n8930 = ~n8921 & n8929;
  assign n8931 = ~Ng11553 & ~n8929;
  assign n4332_1 = ~n8930 & ~n8931;
  assign n8933 = ~Pg3229 & ~n8899;
  assign n8934 = Pg3229 & n8899;
  assign n8935 = ~n8933 & ~n8934;
  assign n8936 = ~n8904 & n8935;
  assign n8937 = ~n8910 & ~n8936;
  assign n8938 = n8894 & n8937;
  assign n8939 = Ng11554 & ~n8894;
  assign n4337_1 = n8938 | n8939;
  assign n8941 = n8925 & n8937;
  assign n8942 = Ng11555 & ~n8925;
  assign n4342 = n8941 | n8942;
  assign n8944 = n8929 & n8937;
  assign n8945 = Ng11556 & ~n8929;
  assign n4347_1 = n8944 | n8945;
  assign n8947 = n8909 & ~n8935;
  assign n8948 = n8909 & n8915;
  assign n8949 = n8935 & ~n8948;
  assign n8950 = ~n8947 & ~n8949;
  assign n8951 = n8894 & n8950;
  assign n8952 = ~Ng11557 & ~n8894;
  assign n4352_1 = ~n8951 & ~n8952;
  assign n8954 = n8925 & ~n8950;
  assign n8955 = Ng11558 & ~n8925;
  assign n4357_1 = n8954 | n8955;
  assign n8957 = n8929 & n8950;
  assign n8958 = ~Ng11559 & ~n8929;
  assign n4362_1 = ~n8957 & ~n8958;
  assign n8960 = n8904 & n8947;
  assign n8961 = n8894 & ~n8960;
  assign n8962 = Ng11560 & ~n8894;
  assign n4367 = n8961 | n8962;
  assign n8964 = n8925 & ~n8960;
  assign n8965 = Ng11561 & ~n8925;
  assign n4372 = n8964 | n8965;
  assign n8967 = n8929 & ~n8960;
  assign n8968 = Ng11562 & ~n8929;
  assign n4377 = n8967 | n8968;
  assign n8970 = ~n8343 & n8388;
  assign n8971 = ~n8329 & n8970;
  assign n8972 = Ng853 & Ng1804;
  assign n8973 = \[1612]  & Ng1798;
  assign n8974 = \[1594]  & Ng1801;
  assign n8975 = ~n8973 & ~n8974;
  assign n4627 = n8972 | ~n8975;
  assign n8977 = ~n8641 & ~n4627;
  assign n8978 = n8971 & n8977;
  assign n8979 = ~n8971 & n4627;
  assign n8980 = ~n8978 & ~n8979;
  assign n8981 = Ng853 & Ng1795;
  assign n8982 = \[1612]  & Ng1789;
  assign n8983 = \[1594]  & Ng1792;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = ~n8981 & n8984;
  assign n8986 = Ng2257 & n8985;
  assign n8987 = ~n8980 & n8986;
  assign n8988 = Ng853 & ~Ng1807;
  assign n8989 = \[1612]  & ~Ng1808;
  assign n8990 = \[1594]  & ~Ng1809;
  assign n8991 = ~n8989 & ~n8990;
  assign n8992 = ~n8988 & n8991;
  assign n8993 = ~n8980 & n8992;
  assign n8994 = Ng2257 & ~n8993;
  assign n8995 = ~n8985 & ~n8994;
  assign n8996 = ~n8987 & ~n8995;
  assign n8997 = \[1612]  & n8996;
  assign n8998 = ~\[1612]  & ~Ng1789;
  assign n4382 = ~n8997 & ~n8998;
  assign n9000 = \[1594]  & n8996;
  assign n9001 = ~\[1594]  & ~Ng1792;
  assign n4387 = ~n9000 & ~n9001;
  assign n9003 = Ng853 & n8996;
  assign n9004 = ~Ng853 & ~Ng1795;
  assign n4392 = ~n9003 & ~n9004;
  assign n9006 = ~\[1612]  & Ng1798;
  assign n9007 = Ng2257 & ~n8985;
  assign n9008 = ~n8992 & n9007;
  assign n9009 = n4627 & ~n9008;
  assign n9010 = ~n8641 & ~n9008;
  assign n9011 = n8971 & ~n9010;
  assign n9012 = ~n9009 & ~n9011;
  assign n9013 = \[1612]  & ~n9012;
  assign n4397 = n9006 | n9013;
  assign n9015 = ~\[1594]  & Ng1801;
  assign n9016 = \[1594]  & ~n9012;
  assign n4402 = n9015 | n9016;
  assign n9018 = ~Ng853 & Ng1804;
  assign n9019 = Ng853 & ~n9012;
  assign n4407 = n9018 | n9019;
  assign n9021 = n8993 & n9007;
  assign n9022 = \[1612]  & n9021;
  assign n9023 = \[1612]  & n8987;
  assign n9024 = ~Ng1808 & ~n9023;
  assign n4412 = ~n9022 & ~n9024;
  assign n9026 = \[1594]  & n9021;
  assign n9027 = \[1594]  & n8987;
  assign n9028 = ~Ng1809 & ~n9027;
  assign n4417 = ~n9026 & ~n9028;
  assign n9030 = Ng853 & n9021;
  assign n9031 = Ng853 & n8987;
  assign n9032 = ~Ng1807 & ~n9031;
  assign n4422 = ~n9030 & ~n9032;
  assign n9034 = ~\[1612]  & Ng1810;
  assign n9035 = Ng853 & ~Ng1559;
  assign n9036 = \[1612]  & ~Ng1560;
  assign n9037 = \[1594]  & ~Ng1561;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~n9035 & n9038;
  assign n9040 = n8388 & ~n9039;
  assign n9041 = Ng2257 & n9040;
  assign n9042 = Ng853 & Ng1816;
  assign n9043 = \[1612]  & Ng1810;
  assign n9044 = \[1594]  & Ng1813;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = ~n9042 & n9045;
  assign n9047 = ~Ng2257 & ~n9046;
  assign n9048 = ~n9041 & ~n9047;
  assign n9049 = \[1612]  & ~n9048;
  assign n4427 = n9034 | n9049;
  assign n9051 = ~\[1594]  & Ng1813;
  assign n9052 = \[1594]  & ~n9048;
  assign n4432 = n9051 | n9052;
  assign n9054 = ~Ng853 & Ng1816;
  assign n9055 = Ng853 & ~n9048;
  assign n4437 = n9054 | n9055;
  assign n9057 = ~\[1612]  & ~Ng1819;
  assign n9058 = Ng853 & Ng1825;
  assign n9059 = \[1612]  & Ng1819;
  assign n9060 = \[1594]  & Ng1822;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = ~n9058 & n9061;
  assign n9063 = Ng853 & ~Ng1828;
  assign n9064 = \[1612]  & ~Ng1829;
  assign n9065 = \[1594]  & ~Ng1830;
  assign n9066 = ~n9064 & ~n9065;
  assign n9067 = ~n9063 & n9066;
  assign n9068 = n9040 & n9062;
  assign n9069 = ~n9046 & ~n9068;
  assign n9070 = ~n9040 & ~n9062;
  assign n9071 = n9046 & ~n9070;
  assign n9072 = Ng2257 & ~n9071;
  assign n9073 = ~n9069 & n9072;
  assign n9074 = ~n9067 & n9073;
  assign n9075 = n9062 & n9074;
  assign n9076 = ~n9062 & ~n9074;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = \[1612]  & n9077;
  assign n4442_1 = ~n9057 & ~n9078;
  assign n9080 = ~\[1594]  & ~Ng1822;
  assign n9081 = \[1594]  & n9077;
  assign n4447_1 = ~n9080 & ~n9081;
  assign n9083 = ~Ng853 & ~Ng1825;
  assign n9084 = Ng853 & n9077;
  assign n4452_1 = ~n9083 & ~n9084;
  assign n9086 = n9067 & n9073;
  assign n9087 = \[1612]  & n9086;
  assign n9088 = n9046 & ~n9068;
  assign n9089 = ~n9046 & ~n9070;
  assign n9090 = Ng2257 & ~n9089;
  assign n9091 = ~n9088 & n9090;
  assign n9092 = \[1612]  & n9091;
  assign n9093 = ~Ng1829 & ~n9092;
  assign n4457 = ~n9087 & ~n9093;
  assign n9095 = \[1594]  & n9086;
  assign n9096 = \[1594]  & n9091;
  assign n9097 = ~Ng1830 & ~n9096;
  assign n4462 = ~n9095 & ~n9097;
  assign n9099 = Ng853 & n9086;
  assign n9100 = Ng853 & n9091;
  assign n9101 = ~Ng1828 & ~n9100;
  assign n4467 = ~n9099 & ~n9101;
  assign n9103 = ~\[1612]  & ~Ng1693;
  assign n9104 = ~n8412 & ~n8443;
  assign n9105 = ~n8477 & ~n9104;
  assign n9106 = ~n8540 & ~n9105;
  assign n9107 = ~n8653 & ~n9106;
  assign n9108 = ~n8648 & ~n9107;
  assign n9109 = \[1612]  & ~n9108;
  assign n4472 = ~n9103 & ~n9109;
  assign n9111 = ~\[1594]  & ~Ng1694;
  assign n9112 = \[1594]  & ~n9108;
  assign n4477 = ~n9111 & ~n9112;
  assign n9114 = ~Ng853 & ~Ng1695;
  assign n9115 = Ng853 & ~n9108;
  assign n4482 = ~n9114 & ~n9115;
  assign n9117 = ~\[1612]  & ~Ng1696;
  assign n9118 = n8540 & n8638;
  assign n9119 = ~n8496 & n8534;
  assign n9120 = n8508 & n9119;
  assign n9121 = n8509 & n8527;
  assign n9122 = n9120 & n9121;
  assign n9123 = n8520 & n9122;
  assign n9124 = ~n8482 & ~n9123;
  assign n9125 = Ng2257 & ~n9124;
  assign n9126 = n8407 & ~n8513;
  assign n9127 = ~n9125 & n9126;
  assign n9128 = ~n8638 & ~n8641;
  assign n9129 = ~n8407 & n9128;
  assign n9130 = ~n9127 & ~n9129;
  assign n9131 = ~n9118 & ~n9130;
  assign n9132 = n8475 & ~n9131;
  assign n9133 = n8483 & ~n9123;
  assign n9134 = n9126 & n9133;
  assign n9135 = ~n8443 & ~n8539;
  assign n9136 = ~n9134 & n9135;
  assign n9137 = ~n8413 & ~n8648;
  assign n9138 = ~n9136 & n9137;
  assign n9139 = ~n9132 & n9138;
  assign n9140 = ~n8890 & n9139;
  assign n9141 = \[1612]  & ~n9140;
  assign n4487 = ~n9117 & ~n9141;
  assign n9143 = ~\[1594]  & ~Ng1697;
  assign n9144 = \[1594]  & ~n9140;
  assign n4492 = ~n9143 & ~n9144;
  assign n9146 = ~Ng853 & ~Ng1698;
  assign n9147 = Ng853 & ~n9140;
  assign n4497 = ~n9146 & ~n9147;
  assign n9149 = ~\[1612]  & ~Ng1699;
  assign n9150 = ~n8443 & n9125;
  assign n9151 = Ng2257 & n8443;
  assign n9152 = n8540 & n9151;
  assign n9153 = n8477 & ~n9152;
  assign n9154 = ~n9150 & n9153;
  assign n9155 = ~n8407 & n9133;
  assign n9156 = n9104 & n9155;
  assign n9157 = ~n9154 & ~n9156;
  assign n9158 = ~n8648 & ~n9157;
  assign n9159 = \[1612]  & ~n9158;
  assign n4502 = ~n9149 & ~n9159;
  assign n9161 = ~\[1594]  & ~Ng1700;
  assign n9162 = \[1594]  & ~n9158;
  assign n4507 = ~n9161 & ~n9162;
  assign n9164 = ~Ng853 & ~Ng1701;
  assign n9165 = Ng853 & ~n9158;
  assign n4512 = ~n9164 & ~n9165;
  assign n9167 = ~n8476 & ~n9124;
  assign n9168 = n5019_1 & ~n9167;
  assign n9169 = ~n8542 & n8632;
  assign n9170 = n9168 & ~n9169;
  assign n9171 = Ng1703 & ~n9168;
  assign n4517 = n9170 | n9171;
  assign n9173 = n5023 & ~n9167;
  assign n9174 = n9169 & n9173;
  assign n9175 = ~Ng1704 & ~n9173;
  assign n4522 = ~n9174 & ~n9175;
  assign n9177 = n5027 & ~n9167;
  assign n9178 = Ng1702 & ~n9177;
  assign n9179 = ~n9169 & n9177;
  assign n4527 = n9178 | n9179;
  assign n9181 = n8632 & n8647;
  assign n9182 = n5019_1 & ~n9181;
  assign n9183 = Ng1784 & ~n5019_1;
  assign n4532 = n9182 | n9183;
  assign n9185 = n5023 & ~n9181;
  assign n9186 = Ng1785 & ~n5023;
  assign n4537 = n9185 | n9186;
  assign n9188 = n5027 & ~n9181;
  assign n9189 = Ng1783 & ~n5027;
  assign n4542 = n9188 | n9189;
  assign n9191 = \[1594]  & ~n3125_1;
  assign n9192 = ~\[1594]  & ~Ng1686;
  assign n9193 = Ng1680 & ~n9192;
  assign n9194 = ~n9191 & n9193;
  assign n9195 = ~Ng1680 & ~Ng1679;
  assign n4632 = n9194 | n9195;
  assign n9197 = Ng1453 & n8459;
  assign n9198 = ~Ng1448 & ~n8435;
  assign n9199 = ~Ng1453 & ~n8459;
  assign n9200 = ~n9198 & ~n9199;
  assign n9201 = Ng1426 & n8454;
  assign n9202 = ~Ng1426 & ~n8454;
  assign n9203 = ~n9201 & ~n9202;
  assign n9204 = n9200 & n9203;
  assign n9205 = Ng1444 & n8430;
  assign n9206 = ~Ng1444 & ~n8430;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = n9204 & n9207;
  assign n9209 = ~n9197 & n9208;
  assign n9210 = ~Ng1435 & ~n8419;
  assign n9211 = Ng1439 & n8424;
  assign n9212 = ~Ng1439 & ~n8424;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9210 & n9213;
  assign n9215 = Ng1430 & ~n8471;
  assign n9216 = ~Ng1430 & n8471;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = Ng1462 & n8466;
  assign n9219 = ~Ng1462 & ~n8466;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = ~n9217 & n9220;
  assign n9222 = Ng1435 & n8419;
  assign n9223 = Ng1457 & ~n8448;
  assign n9224 = ~Ng1457 & n8448;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n9222 & ~n9225;
  assign n9227 = n9221 & n9226;
  assign n9228 = n9214 & n9227;
  assign n9229 = Ng1448 & n8435;
  assign n9230 = n8892 & ~n9229;
  assign n9231 = ~Ng1466 & n8402;
  assign n9232 = Ng1466 & ~n8402;
  assign n9233 = ~n9231 & ~n9232;
  assign n9234 = n9230 & ~n9233;
  assign n9235 = n9228 & n9234;
  assign n9236 = n9209 & n9235;
  assign n4637 = ~n8474 & ~n9236;
  assign n9238 = ~Ng1315 & Ng1934;
  assign n4738 = n6033 | n9238;
  assign n9240 = Ng1315 & Ng1934;
  assign n9241 = ~Ng1315 & ~Ng1937;
  assign n4743 = ~n9240 & ~n9241;
  assign n9243 = Ng1315 & Ng1937;
  assign n9244 = ~Ng1315 & Ng1890;
  assign n4748 = n9243 | n9244;
  assign n9246 = Ng1315 & Ng1953;
  assign n9247 = \[1605]  & Ng1949;
  assign n9248 = \[1603]  & Ng1951;
  assign n9249 = ~n9247 & ~n9248;
  assign n4753 = ~n9246 & n9249;
  assign n9251 = ~\[1612]  & Ng1867;
  assign n9252 = \[1612]  & ~n9062;
  assign n4820 = n9251 | n9252;
  assign n9254 = ~\[1594]  & Ng1868;
  assign n9255 = \[1594]  & ~n9062;
  assign n4825 = n9254 | n9255;
  assign n9257 = ~Ng853 & Ng1869;
  assign n9258 = Ng853 & ~n9062;
  assign n4830 = n9257 | n9258;
  assign n9260 = ~\[1612]  & ~Ng11566;
  assign n9261 = \[1612]  & ~n8891;
  assign n4835 = ~n9260 & ~n9261;
  assign n9263 = ~\[1594]  & ~Ng11569;
  assign n9264 = \[1594]  & ~n8891;
  assign n4839 = ~n9263 & ~n9264;
  assign n9266 = ~Ng853 & ~Ng11570;
  assign n9267 = Ng853 & ~n8891;
  assign n4843 = ~n9266 & ~n9267;
  assign n9269 = ~\[1612]  & ~Ng1858;
  assign n9270 = \[1612]  & ~n8476;
  assign n4847 = ~n9269 & ~n9270;
  assign n9272 = ~\[1594]  & ~Ng1859;
  assign n9273 = \[1594]  & ~n8476;
  assign n4852 = ~n9272 & ~n9273;
  assign n9275 = ~Ng853 & ~Ng1860;
  assign n9276 = Ng853 & ~n8476;
  assign n4857 = ~n9275 & ~n9276;
  assign n9278 = ~\[1612]  & ~Ng1861;
  assign n9279 = \[1612]  & n4627;
  assign n4862 = ~n9278 & ~n9279;
  assign n9281 = ~\[1594]  & ~Ng1865;
  assign n9282 = \[1594]  & n4627;
  assign n4867 = ~n9281 & ~n9282;
  assign n9284 = ~Ng853 & ~Ng1845;
  assign n9285 = Ng853 & n4627;
  assign n4872_1 = ~n9284 & ~n9285;
  assign n9287 = ~\[1612]  & ~Ng11571;
  assign n9288 = \[1612]  & ~n8889;
  assign n4877 = ~n9287 & ~n9288;
  assign n9290 = ~\[1594]  & ~Ng11567;
  assign n9291 = \[1594]  & ~n8889;
  assign n4881 = ~n9290 & ~n9291;
  assign n9293 = ~Ng853 & ~Ng11568;
  assign n9294 = Ng853 & ~n8889;
  assign n4885 = ~n9293 & ~n9294;
  assign n9296 = Ng1315 & Ng1870;
  assign n9297 = \[1605]  & Ng1945;
  assign n9298 = \[1603]  & Ng1947;
  assign n9299 = ~n9297 & ~n9298;
  assign n4889 = ~n9296 & n9299;
  assign n9301 = \[1605]  & ~Ng1860;
  assign n9302 = \[1603]  & ~Ng1858;
  assign n9303 = Ng1315 & ~Ng1859;
  assign n9304 = ~n9302 & ~n9303;
  assign n4902 = ~n9301 & n9304;
  assign n9306 = \[1605]  & ~Ng1845;
  assign n9307 = \[1603]  & ~Ng1861;
  assign n9308 = Ng1315 & ~Ng1865;
  assign n9309 = ~n9307 & ~n9308;
  assign n4916 = ~n9306 & n9309;
  assign n9311 = \[1605]  & ~Ng1869;
  assign n9312 = \[1603]  & ~Ng1867;
  assign n9313 = Ng1315 & ~Ng1868;
  assign n9314 = ~n9312 & ~n9313;
  assign n4925 = ~n9311 & n9314;
  assign n9316 = Ng1315 & Ng2000;
  assign n9317 = \[1605]  & Ng1994;
  assign n9318 = \[1603]  & Ng1997;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = ~n9316 & n9319;
  assign n9321 = Ng1315 & Ng1877;
  assign n9322 = \[1605]  & Ng1871;
  assign n9323 = \[1603]  & Ng1874;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = ~n9321 & n9324;
  assign n9326 = Ng1890 & n9325;
  assign n9327 = ~n9320 & n9326;
  assign n9328 = Ng1315 & Ng1991;
  assign n9329 = \[1605]  & Ng1985;
  assign n9330 = \[1603]  & Ng1988;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~n9328 & n9331;
  assign n9333 = ~n9325 & ~n9332;
  assign n9334 = ~n6126 & ~n9333;
  assign n5073 = n9327 | n9334;
  assign n9336 = \[1605]  & n5073;
  assign n9337 = ~Ng1956 & ~n9336;
  assign n9338 = Ng1315 & ~Ng1964;
  assign n9339 = \[1605]  & ~Ng1965;
  assign n9340 = \[1603]  & ~Ng1966;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n9338 & n9341;
  assign n9343 = Pg3229 & ~n9342;
  assign n9344 = Ng1315 & ~Ng1961;
  assign n9345 = \[1605]  & ~Ng1962;
  assign n9346 = \[1603]  & ~Ng1963;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = ~n9344 & n9347;
  assign n9349 = Ng1315 & ~Ng1958;
  assign n9350 = \[1605]  & ~Ng1959;
  assign n9351 = \[1603]  & ~Ng1960;
  assign n9352 = ~n9350 & ~n9351;
  assign n9353 = ~n9349 & n9352;
  assign n9354 = n9348 & ~n9353;
  assign n9355 = Ng1315 & ~Ng1955;
  assign n9356 = \[1605]  & ~Ng1956;
  assign n9357 = \[1603]  & ~Ng1957;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = ~n9355 & n9358;
  assign n9360 = n9342 & ~n9359;
  assign n9361 = ~n9354 & n9360;
  assign n9362 = ~Pg3229 & n9354;
  assign n9363 = ~n9361 & ~n9362;
  assign n9364 = ~n9343 & n9363;
  assign n9365 = n9336 & ~n9364;
  assign n4934 = ~n9337 & ~n9365;
  assign n9367 = \[1603]  & n5073;
  assign n9368 = ~n9364 & n9367;
  assign n9369 = ~Ng1957 & ~n9367;
  assign n4939 = ~n9368 & ~n9369;
  assign n9371 = Ng1315 & n5073;
  assign n9372 = ~n9364 & n9371;
  assign n9373 = ~Ng1955 & ~n9371;
  assign n4944 = ~n9372 & ~n9373;
  assign n9375 = ~Pg3229 & ~n9359;
  assign n9376 = Pg3229 & n9359;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = ~n9348 & n9377;
  assign n9379 = ~n9354 & ~n9378;
  assign n9380 = n9336 & n9379;
  assign n9381 = Ng1959 & ~n9336;
  assign n4949 = n9380 | n9381;
  assign n9383 = n9367 & n9379;
  assign n9384 = Ng1960 & ~n9367;
  assign n4954 = n9383 | n9384;
  assign n9386 = n9371 & n9379;
  assign n9387 = Ng1958 & ~n9371;
  assign n4959 = n9386 | n9387;
  assign n9389 = n9342 & n9353;
  assign n9390 = n9377 & ~n9389;
  assign n9391 = n9353 & ~n9377;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = n9336 & ~n9392;
  assign n9394 = Ng1962 & ~n9336;
  assign n4964 = n9393 | n9394;
  assign n9396 = n9367 & ~n9392;
  assign n9397 = Ng1963 & ~n9367;
  assign n4969 = n9396 | n9397;
  assign n9399 = n9371 & ~n9392;
  assign n9400 = Ng1961 & ~n9371;
  assign n4974 = n9399 | n9400;
  assign n9402 = n9348 & n9353;
  assign n9403 = ~n9377 & n9402;
  assign n9404 = n9336 & ~n9403;
  assign n9405 = Ng1965 & ~n9336;
  assign n4979 = n9404 | n9405;
  assign n9407 = n9367 & ~n9403;
  assign n9408 = Ng1966 & ~n9367;
  assign n4984 = n9407 | n9408;
  assign n9410 = n9371 & ~n9403;
  assign n9411 = Ng1964 & ~n9371;
  assign n4989 = n9410 | n9411;
  assign n9413 = ~\[1605]  & ~Ng1967;
  assign n9414 = Ng185 & Ng1904;
  assign n9415 = ~n4753 & n9414;
  assign n9416 = \[1603]  & Ng1970;
  assign n9417 = Ng1315 & Ng1973;
  assign n9418 = \[1605]  & Ng1967;
  assign n9419 = ~n9417 & ~n9418;
  assign n9420 = ~n9416 & n9419;
  assign n9421 = ~n9415 & n9420;
  assign n9422 = ~n6032 & ~n9421;
  assign n9423 = \[1605]  & ~n9422;
  assign n4994 = ~n9413 & ~n9423;
  assign n9425 = ~\[1603]  & ~Ng1970;
  assign n9426 = \[1603]  & ~n9422;
  assign n4999 = ~n9425 & ~n9426;
  assign n9428 = ~Ng1315 & Ng1973;
  assign n9429 = n6033 & ~n9421;
  assign n5004 = n9428 | n9429;
  assign n9431 = ~\[1605]  & ~Ng1976;
  assign n9432 = Ng185 & Ng1922;
  assign n9433 = ~n4889 & n9432;
  assign n9434 = Ng1315 & Ng1982;
  assign n9435 = \[1603]  & Ng1979;
  assign n9436 = \[1605]  & Ng1976;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = ~n9434 & n9437;
  assign n9439 = ~n9433 & n9438;
  assign n9440 = ~n6032 & ~n9439;
  assign n9441 = \[1605]  & ~n9440;
  assign n5009 = ~n9431 & ~n9441;
  assign n9443 = ~\[1603]  & ~Ng1979;
  assign n9444 = \[1603]  & ~n9440;
  assign n5014 = ~n9443 & ~n9444;
  assign n9446 = ~Ng1315 & Ng1982;
  assign n9447 = n6033 & ~n9439;
  assign n5019 = n9446 | n9447;
  assign n9449 = ~\[1605]  & Ng1994;
  assign n9450 = ~n6032 & ~n9320;
  assign n9451 = ~n9421 & ~n9439;
  assign n9452 = n6032 & ~n9451;
  assign n9453 = Ng1315 & Ng1749;
  assign n9454 = \[1605]  & Ng1745;
  assign n9455 = \[1603]  & Ng1747;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = ~n9453 & n9456;
  assign n9458 = Ng1315 & Ng1764;
  assign n9459 = \[1605]  & Ng1760;
  assign n9460 = \[1603]  & Ng1762;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9458 & n9461;
  assign n9463 = n9359 & ~n9462;
  assign n9464 = Ng1315 & Ng1734;
  assign n9465 = \[1605]  & Ng1730;
  assign n9466 = \[1603]  & Ng1732;
  assign n9467 = ~n9465 & ~n9466;
  assign n9468 = ~n9464 & n9467;
  assign n9469 = n9348 & n9468;
  assign n9470 = ~n9463 & ~n9469;
  assign n9471 = n9457 & ~n9470;
  assign n9472 = ~n9353 & n9471;
  assign n9473 = ~n9457 & ~n9462;
  assign n9474 = ~n9342 & n9473;
  assign n9475 = ~n9348 & n9457;
  assign n9476 = n9389 & n9462;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = Ng1315 & Ng1705;
  assign n9479 = \[1605]  & Ng1775;
  assign n9480 = \[1603]  & Ng1777;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = ~n9478 & n9481;
  assign n9483 = ~n9457 & ~n9482;
  assign n9484 = n9348 & n9483;
  assign n9485 = n9353 & n9484;
  assign n9486 = n9477 & ~n9485;
  assign n9487 = n9359 & ~n9486;
  assign n9488 = ~n9474 & ~n9487;
  assign n9489 = ~n9468 & ~n9488;
  assign n9490 = n9402 & n9482;
  assign n9491 = n9389 & n9473;
  assign n9492 = ~n9348 & n9483;
  assign n9493 = ~n9353 & n9462;
  assign n9494 = ~n9492 & ~n9493;
  assign n9495 = ~n9491 & n9494;
  assign n9496 = n9468 & ~n9495;
  assign n9497 = ~n9490 & ~n9496;
  assign n9498 = ~n9359 & ~n9497;
  assign n9499 = ~n9489 & ~n9498;
  assign n9500 = ~n9472 & n9499;
  assign n9501 = n9342 & ~n9468;
  assign n9502 = n9348 & ~n9501;
  assign n9503 = n9482 & ~n9502;
  assign n9504 = n9348 & ~n9468;
  assign n9505 = ~n9353 & n9468;
  assign n9506 = ~n9504 & ~n9505;
  assign n9507 = n9473 & n9506;
  assign n9508 = ~n9503 & ~n9507;
  assign n9509 = n9359 & ~n9508;
  assign n9510 = n9402 & ~n9457;
  assign n9511 = n9342 & ~n9510;
  assign n9512 = ~n9342 & ~n9482;
  assign n9513 = ~n9462 & ~n9512;
  assign n9514 = ~n9463 & ~n9513;
  assign n9515 = n9468 & n9514;
  assign n9516 = ~n9511 & n9515;
  assign n9517 = ~n9509 & ~n9516;
  assign n9518 = n9462 & ~n9475;
  assign n9519 = ~n9484 & ~n9518;
  assign n9520 = ~n9353 & ~n9519;
  assign n9521 = ~n9468 & n9520;
  assign n9522 = ~n9462 & ~n9502;
  assign n9523 = ~n9506 & ~n9522;
  assign n9524 = ~n9359 & n9457;
  assign n9525 = ~n9523 & n9524;
  assign n9526 = ~n9521 & ~n9525;
  assign n9527 = n9517 & n9526;
  assign n9528 = n9439 & n9527;
  assign n9529 = n9500 & ~n9528;
  assign n9530 = n9452 & n9529;
  assign n9531 = ~n9450 & ~n9530;
  assign n9532 = \[1605]  & ~n9531;
  assign n5024 = n9449 | n9532;
  assign n9534 = ~\[1603]  & Ng1997;
  assign n9535 = \[1603]  & ~n9531;
  assign n5029 = n9534 | n9535;
  assign n9537 = ~Ng1315 & Ng2000;
  assign n9538 = Ng1315 & ~n9531;
  assign n5034 = n9537 | n9538;
  assign n9540 = ~\[1605]  & Ng1985;
  assign n9541 = ~n6032 & ~n9332;
  assign n9542 = n9421 & n9500;
  assign n9543 = n9452 & n9527;
  assign n9544 = ~n9542 & n9543;
  assign n9545 = ~n9541 & ~n9544;
  assign n9546 = \[1605]  & ~n9545;
  assign n5039 = n9540 | n9546;
  assign n9548 = ~\[1603]  & Ng1988;
  assign n9549 = \[1603]  & ~n9545;
  assign n5044 = n9548 | n9549;
  assign n9551 = ~Ng1315 & Ng1991;
  assign n9552 = Ng1315 & ~n9545;
  assign n5049 = n9551 | n9552;
  assign n9554 = ~\[1605]  & ~Ng1871;
  assign n9555 = n9320 & n9326;
  assign n9556 = \[1605]  & ~n9555;
  assign n5054 = ~n9554 & ~n9556;
  assign n9558 = ~\[1603]  & ~Ng1874;
  assign n9559 = \[1603]  & ~n9555;
  assign n5059 = ~n9558 & ~n9559;
  assign n9561 = ~Ng1315 & ~Ng1877;
  assign n9562 = Ng1315 & ~n9555;
  assign n5064 = ~n9561 & ~n9562;
  assign n9564 = Ng1886 & ~Ng1887;
  assign n9565 = \[1603]  & n3571_1;
  assign n9566 = ~\[1603]  & Pg16399;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = ~Ng1886 & n9567;
  assign n5078 = ~n9564 & ~n9568;
  assign n9570 = Pg3229 & Ng1672;
  assign n9571 = ~Pg3229 & ~Ng1686;
  assign n5126 = ~n9570 & ~n9571;
  assign n9573 = Ng1315 & Ng1890;
  assign n9574 = ~Ng1315 & Ng2010;
  assign n5136 = n9573 | n9574;
  assign n9576 = ~Ng1315 & ~Ng2039;
  assign n5141 = ~n6374_1 & ~n9576;
  assign n9578 = \[1603]  & Ng2010;
  assign n9579 = Ng1315 & ~Ng2039;
  assign n9580 = Ng2020 & n9579;
  assign n9581 = ~Ng2020 & ~n9579;
  assign n9582 = ~n9580 & ~n9581;
  assign n5146 = ~n9578 & n9582;
  assign n9584 = Ng2013 & n9580;
  assign n9585 = ~Ng2013 & ~n9580;
  assign n9586 = ~n9578 & ~n9585;
  assign n5151 = ~n9584 & n9586;
  assign n9588 = Ng2033 & n9584;
  assign n9589 = ~Ng2033 & ~n9584;
  assign n9590 = ~n9578 & ~n9589;
  assign n5156 = ~n9588 & n9590;
  assign n9592 = Ng2026 & n9588;
  assign n9593 = ~Ng2026 & ~n9588;
  assign n9594 = ~n9578 & ~n9593;
  assign n5161 = ~n9592 & n9594;
  assign n9596 = Ng2040 & n9592;
  assign n9597 = ~Ng2040 & ~n9592;
  assign n9598 = ~n9578 & ~n9597;
  assign n5166 = ~n9596 & n9598;
  assign n9600 = Ng2052 & n9596;
  assign n9601 = ~Ng2052 & ~n9596;
  assign n9602 = ~n9578 & ~n9601;
  assign n5171 = ~n9600 & n9602;
  assign n9604 = Ng2046 & n9600;
  assign n9605 = ~Ng2046 & ~n9600;
  assign n9606 = ~n9578 & ~n9605;
  assign n5176 = ~n9604 & n9606;
  assign n9608 = Ng2059 & n9604;
  assign n9609 = ~Ng2059 & ~n9604;
  assign n9610 = ~n9578 & ~n9609;
  assign n5181 = ~n9608 & n9610;
  assign n9612 = Ng2066 & n9608;
  assign n9613 = ~Ng2066 & ~n9608;
  assign n9614 = ~n9578 & ~n9613;
  assign n5186 = ~n9612 & n9614;
  assign n9616 = Ng2072 & n9612;
  assign n9617 = ~Ng2072 & ~n9612;
  assign n9618 = ~n9616 & ~n9617;
  assign n5191 = ~n9578 & n9618;
  assign n9620 = Ng1905 & ~Ng2039;
  assign n9621 = Ng1918 & n9620;
  assign n9622 = \[1605]  & n9621;
  assign n9623 = Ng2079 & ~n9622;
  assign n9624 = ~Ng2020 & n9622;
  assign n5196 = n9623 | n9624;
  assign n9626 = \[1603]  & n9621;
  assign n9627 = Ng2080 & ~n9626;
  assign n9628 = ~Ng2020 & n9626;
  assign n5201 = n9627 | n9628;
  assign n9630 = Ng1315 & n9621;
  assign n9631 = Ng2078 & ~n9630;
  assign n9632 = ~Ng2020 & n9630;
  assign n5206 = n9631 | n9632;
  assign n9634 = Ng2082 & ~n9622;
  assign n9635 = ~Ng2013 & n9622;
  assign n5211 = n9634 | n9635;
  assign n9637 = Ng2083 & ~n9626;
  assign n9638 = ~Ng2013 & n9626;
  assign n5216 = n9637 | n9638;
  assign n9640 = Ng2081 & ~n9630;
  assign n9641 = ~Ng2013 & n9630;
  assign n5221 = n9640 | n9641;
  assign n9643 = Ng2085 & ~n9622;
  assign n9644 = ~Ng2033 & n9622;
  assign n5226 = n9643 | n9644;
  assign n9646 = Ng2086 & ~n9626;
  assign n9647 = ~Ng2033 & n9626;
  assign n5231 = n9646 | n9647;
  assign n9649 = Ng2084 & ~n9630;
  assign n9650 = ~Ng2033 & n9630;
  assign n5236 = n9649 | n9650;
  assign n9652 = Ng2088 & ~n9622;
  assign n9653 = ~Ng2026 & n9622;
  assign n5241 = n9652 | n9653;
  assign n9655 = Ng2089 & ~n9626;
  assign n9656 = ~Ng2026 & n9626;
  assign n5246 = n9655 | n9656;
  assign n9658 = Ng2087 & ~n9630;
  assign n9659 = ~Ng2026 & n9630;
  assign n5251 = n9658 | n9659;
  assign n9661 = Ng2091 & ~n9622;
  assign n9662 = ~Ng2040 & n9622;
  assign n5256 = n9661 | n9662;
  assign n9664 = Ng2092 & ~n9626;
  assign n9665 = ~Ng2040 & n9626;
  assign n5261 = n9664 | n9665;
  assign n9667 = Ng2090 & ~n9630;
  assign n9668 = ~Ng2040 & n9630;
  assign n5266 = n9667 | n9668;
  assign n9670 = Ng2094 & ~n9622;
  assign n9671 = ~Ng2052 & n9622;
  assign n5271 = n9670 | n9671;
  assign n9673 = Ng2095 & ~n9626;
  assign n9674 = ~Ng2052 & n9626;
  assign n5276 = n9673 | n9674;
  assign n9676 = Ng2093 & ~n9630;
  assign n9677 = ~Ng2052 & n9630;
  assign n5281 = n9676 | n9677;
  assign n9679 = Ng2097 & ~n9622;
  assign n9680 = ~Ng2046 & n9622;
  assign n5286 = n9679 | n9680;
  assign n9682 = Ng2098 & ~n9626;
  assign n9683 = ~Ng2046 & n9626;
  assign n5291 = n9682 | n9683;
  assign n9685 = Ng2096 & ~n9630;
  assign n9686 = ~Ng2046 & n9630;
  assign n5296 = n9685 | n9686;
  assign n9688 = Ng2100 & ~n9622;
  assign n9689 = ~Ng2059 & n9622;
  assign n5301 = n9688 | n9689;
  assign n9691 = Ng2101 & ~n9626;
  assign n9692 = ~Ng2059 & n9626;
  assign n5306 = n9691 | n9692;
  assign n9694 = Ng2099 & ~n9630;
  assign n9695 = ~Ng2059 & n9630;
  assign n5311 = n9694 | n9695;
  assign n9697 = Ng2103 & ~n9622;
  assign n9698 = ~Ng2066 & n9622;
  assign n5316 = n9697 | n9698;
  assign n9700 = Ng2104 & ~n9626;
  assign n9701 = ~Ng2066 & n9626;
  assign n5321 = n9700 | n9701;
  assign n9703 = Ng2102 & ~n9630;
  assign n9704 = ~Ng2066 & n9630;
  assign n5326 = n9703 | n9704;
  assign n9706 = Ng2106 & ~n9622;
  assign n9707 = ~Ng2072 & n9622;
  assign n5331 = n9706 | n9707;
  assign n9709 = Ng2107 & ~n9626;
  assign n9710 = ~Ng2072 & n9626;
  assign n5336 = n9709 | n9710;
  assign n9712 = Ng2105 & ~n9630;
  assign n9713 = ~Ng2072 & n9630;
  assign n5341 = n9712 | n9713;
  assign n9715 = \[1605]  & Ng2010;
  assign n9716 = ~Ng2109 & ~n9715;
  assign n9717 = ~n9320 & n9715;
  assign n5346 = ~n9716 & ~n9717;
  assign n9719 = ~Ng2110 & ~n9578;
  assign n9720 = ~n9320 & n9578;
  assign n5351 = ~n9719 & ~n9720;
  assign n9722 = Ng1315 & Ng2010;
  assign n9723 = ~Ng2108 & ~n9722;
  assign n9724 = ~n9320 & n9722;
  assign n5356 = ~n9723 & ~n9724;
  assign n9726 = ~Ng2112 & ~n9715;
  assign n9727 = ~n9332 & n9715;
  assign n5361 = ~n9726 & ~n9727;
  assign n9729 = n9332 & n9578;
  assign n9730 = Ng2113 & ~n9578;
  assign n5366 = n9729 | n9730;
  assign n9732 = ~n9332 & n9722;
  assign n9733 = ~Ng2111 & ~n9722;
  assign n5371 = ~n9732 & ~n9733;
  assign n9735 = Ng1315 & ~Ng2105;
  assign n9736 = \[1605]  & ~Ng2106;
  assign n9737 = \[1603]  & ~Ng2107;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = ~n9735 & n9738;
  assign n9740 = ~Ng2072 & ~n9739;
  assign n9741 = Ng1315 & ~Ng2093;
  assign n9742 = \[1605]  & ~Ng2094;
  assign n9743 = \[1603]  & ~Ng2095;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = ~n9741 & n9744;
  assign n9746 = Ng2052 & n9745;
  assign n9747 = ~Ng2052 & ~n9745;
  assign n9748 = ~n9746 & ~n9747;
  assign n9749 = ~n9740 & n9748;
  assign n9750 = Ng1315 & ~Ng2078;
  assign n9751 = \[1605]  & ~Ng2079;
  assign n9752 = \[1603]  & ~Ng2080;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~n9750 & n9753;
  assign n9755 = ~Ng2020 & ~n9754;
  assign n9756 = Ng1315 & ~Ng2087;
  assign n9757 = \[1605]  & ~Ng2088;
  assign n9758 = \[1603]  & ~Ng2089;
  assign n9759 = ~n9757 & ~n9758;
  assign n9760 = ~n9756 & n9759;
  assign n9761 = ~Ng2026 & ~n9760;
  assign n9762 = ~n9755 & ~n9761;
  assign n9763 = Ng1315 & ~Ng2096;
  assign n9764 = \[1605]  & ~Ng2097;
  assign n9765 = \[1603]  & ~Ng2098;
  assign n9766 = ~n9764 & ~n9765;
  assign n9767 = ~n9763 & n9766;
  assign n9768 = Ng2046 & n9767;
  assign n9769 = n9762 & ~n9768;
  assign n9770 = n9749 & n9769;
  assign n9771 = Ng2026 & n9760;
  assign n9772 = Ng1315 & ~Ng2099;
  assign n9773 = \[1605]  & ~Ng2100;
  assign n9774 = \[1603]  & ~Ng2101;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = ~n9772 & n9775;
  assign n9777 = ~Ng2059 & ~n9776;
  assign n9778 = ~n9771 & ~n9777;
  assign n9779 = Ng1315 & ~Ng2081;
  assign n9780 = \[1605]  & ~Ng2082;
  assign n9781 = \[1603]  & ~Ng2083;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = ~n9779 & n9782;
  assign n9784 = Ng2013 & n9783;
  assign n9785 = ~Ng2013 & ~n9783;
  assign n9786 = ~n9784 & ~n9785;
  assign n9787 = n9778 & n9786;
  assign n9788 = Ng2059 & n9776;
  assign n9789 = Ng1315 & ~Ng2090;
  assign n9790 = \[1605]  & ~Ng2091;
  assign n9791 = \[1603]  & ~Ng2092;
  assign n9792 = ~n9790 & ~n9791;
  assign n9793 = ~n9789 & n9792;
  assign n9794 = Ng2040 & n9793;
  assign n9795 = ~Ng2040 & ~n9793;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = ~n9788 & n9796;
  assign n9798 = n9787 & n9797;
  assign n9799 = n9770 & n9798;
  assign n9800 = Ng1315 & ~Ng2102;
  assign n9801 = \[1605]  & ~Ng2103;
  assign n9802 = \[1603]  & ~Ng2104;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = ~n9800 & n9803;
  assign n9805 = Ng2066 & n9804;
  assign n9806 = ~Ng2066 & ~n9804;
  assign n9807 = ~n9805 & ~n9806;
  assign n9808 = Ng2020 & n9754;
  assign n9809 = Ng2072 & n9739;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = ~Ng2046 & ~n9767;
  assign n9812 = n9810 & ~n9811;
  assign n9813 = Ng1315 & ~Ng2084;
  assign n9814 = \[1605]  & ~Ng2085;
  assign n9815 = \[1603]  & ~Ng2086;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9813 & n9816;
  assign n9818 = Ng2033 & ~n9817;
  assign n9819 = ~Ng2033 & n9817;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = n9812 & ~n9820;
  assign n9822 = n9807 & n9821;
  assign n9823 = n9799 & n9822;
  assign n9824 = Ng1315 & ~Ng2108;
  assign n9825 = Ng1315 & ~Ng2111;
  assign n9826 = \[1605]  & ~Ng2112;
  assign n9827 = \[1603]  & ~Ng2113;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = ~n9825 & n9828;
  assign n9830 = \[1605]  & ~Ng2109;
  assign n9831 = \[1603]  & ~Ng2110;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = n9829 & n9832;
  assign n9834 = ~n9824 & n9833;
  assign n9835 = ~n9823 & n9834;
  assign n9836 = n9622 & n9835;
  assign n9837 = Ng2115 & ~n9622;
  assign n5376 = n9836 | n9837;
  assign n9839 = n9626 & n9835;
  assign n9840 = Ng2116 & ~n9626;
  assign n5381 = n9839 | n9840;
  assign n9842 = n9630 & n9835;
  assign n9843 = Ng2114 & ~n9630;
  assign n5386 = n9842 | n9843;
  assign n9845 = ~Ng2118 & ~n9622;
  assign n5391 = ~n9715 & ~n9845;
  assign n9847 = ~Ng2119 & ~n9626;
  assign n5396 = ~n9578 & ~n9847;
  assign n9849 = ~Ng2117 & ~n9630;
  assign n5401 = ~n9722 & ~n9849;
  assign n9851 = Ng2206 & ~n5019_1;
  assign n9852 = ~Ng2165 & n5019_1;
  assign n5406 = n9851 | n9852;
  assign n9854 = Ng2207 & ~n5023;
  assign n9855 = ~Ng2165 & n5023;
  assign n5411 = n9854 | n9855;
  assign n9857 = Ng2205 & ~n5027;
  assign n9858 = ~Ng2165 & n5027;
  assign n5416 = n9857 | n9858;
  assign n9860 = Ng2209 & ~n5019_1;
  assign n9861 = ~Ng2170 & n5019_1;
  assign n5421 = n9860 | n9861;
  assign n9863 = Ng2210 & ~n5023;
  assign n9864 = ~Ng2170 & n5023;
  assign n5426 = n9863 | n9864;
  assign n9866 = Ng2208 & ~n5027;
  assign n9867 = ~Ng2170 & n5027;
  assign n5431 = n9866 | n9867;
  assign n9869 = Ng2218 & ~n5019_1;
  assign n9870 = ~Ng2175 & n5019_1;
  assign n5436 = n9869 | n9870;
  assign n9872 = Ng2219 & ~n5023;
  assign n9873 = ~Ng2175 & n5023;
  assign n5441 = n9872 | n9873;
  assign n9875 = Ng2217 & ~n5027;
  assign n9876 = ~Ng2175 & n5027;
  assign n5446 = n9875 | n9876;
  assign n9878 = Ng2221 & ~n5019_1;
  assign n9879 = ~Ng2180 & n5019_1;
  assign n5451 = n9878 | n9879;
  assign n9881 = Ng2222 & ~n5023;
  assign n9882 = ~Ng2180 & n5023;
  assign n5456 = n9881 | n9882;
  assign n9884 = Ng2220 & ~n5027;
  assign n9885 = ~Ng2180 & n5027;
  assign n5461 = n9884 | n9885;
  assign n9887 = Ng2224 & ~n5019_1;
  assign n9888 = ~Ng2185 & n5019_1;
  assign n5466 = n9887 | n9888;
  assign n9890 = Ng2225 & ~n5023;
  assign n9891 = ~Ng2185 & n5023;
  assign n5471 = n9890 | n9891;
  assign n9893 = Ng2223 & ~n5027;
  assign n9894 = ~Ng2185 & n5027;
  assign n5476 = n9893 | n9894;
  assign n9896 = Ng2227 & ~n5019_1;
  assign n9897 = ~Ng2190 & n5019_1;
  assign n5481 = n9896 | n9897;
  assign n9899 = Ng2228 & ~n5023;
  assign n9900 = ~Ng2190 & n5023;
  assign n5486 = n9899 | n9900;
  assign n9902 = Ng2226 & ~n5027;
  assign n9903 = ~Ng2190 & n5027;
  assign n5491 = n9902 | n9903;
  assign n9905 = Ng2230 & ~n5019_1;
  assign n9906 = ~Ng2195 & n5019_1;
  assign n5496 = n9905 | n9906;
  assign n9908 = Ng2231 & ~n5023;
  assign n9909 = ~Ng2195 & n5023;
  assign n5501 = n9908 | n9909;
  assign n9911 = Ng2229 & ~n5027;
  assign n9912 = ~Ng2195 & n5027;
  assign n5506 = n9911 | n9912;
  assign n9914 = Ng2233 & ~n5019_1;
  assign n9915 = ~Ng2200 & n5019_1;
  assign n5511 = n9914 | n9915;
  assign n9917 = Ng2234 & ~n5023;
  assign n9918 = ~Ng2200 & n5023;
  assign n5516 = n9917 | n9918;
  assign n9920 = Ng2232 & ~n5027;
  assign n9921 = ~Ng2200 & n5027;
  assign n5521 = n9920 | n9921;
  assign n9923 = ~Ng2236 & ~n5019_1;
  assign n9924 = Ng853 & ~Ng2250;
  assign n9925 = \[1612]  & ~Ng2251;
  assign n9926 = \[1594]  & ~Ng2252;
  assign n9927 = ~n9925 & ~n9926;
  assign n9928 = ~n9924 & n9927;
  assign n9929 = n5019_1 & ~n9928;
  assign n5526 = ~n9923 & ~n9929;
  assign n9931 = n5023 & n9928;
  assign n9932 = Ng2237 & ~n5023;
  assign n5531 = n9931 | n9932;
  assign n9934 = ~Ng2235 & ~n5027;
  assign n9935 = n5027 & ~n9928;
  assign n5536 = ~n9934 & ~n9935;
  assign n9937 = ~Ng2239 & ~n5019_1;
  assign n9938 = Ng853 & ~Ng2247;
  assign n9939 = \[1612]  & ~Ng2248;
  assign n9940 = \[1594]  & ~Ng2249;
  assign n9941 = ~n9939 & ~n9940;
  assign n9942 = ~n9938 & n9941;
  assign n9943 = n5019_1 & ~n9942;
  assign n5541 = ~n9937 & ~n9943;
  assign n9945 = n5023 & n9942;
  assign n9946 = Ng2240 & ~n5023;
  assign n5546 = n9945 | n9946;
  assign n9948 = ~Ng2238 & ~n5027;
  assign n9949 = n5027 & ~n9942;
  assign n5551 = ~n9948 & ~n9949;
  assign n9951 = Ng2200 & Ng2185;
  assign n9952 = ~Ng2190 & n9951;
  assign n9953 = ~Ng2195 & n9952;
  assign n9954 = n5131_1 & n9953;
  assign n9955 = Ng2245 & ~n5131_1;
  assign n5556 = n9954 | n9955;
  assign n9957 = n5138 & n9953;
  assign n9958 = Ng2246 & ~n5138;
  assign n5561 = n9957 | n9958;
  assign n9960 = n5142 & n9953;
  assign n9961 = Ng2244 & ~n5142;
  assign n5566 = n9960 | n9961;
  assign n9963 = Ng2248 & ~n5131_1;
  assign n9964 = ~Ng2170 & n5131_1;
  assign n5571 = n9963 | n9964;
  assign n9966 = Ng2249 & ~n5138;
  assign n9967 = ~Ng2170 & n5138;
  assign n5576 = n9966 | n9967;
  assign n9969 = Ng2247 & ~n5142;
  assign n9970 = ~Ng2170 & n5142;
  assign n5581 = n9969 | n9970;
  assign n9972 = Ng2251 & ~n5131_1;
  assign n9973 = ~Ng2165 & n5131_1;
  assign n5586 = n9972 | n9973;
  assign n9975 = Ng2252 & ~n5138;
  assign n9976 = ~Ng2165 & n5138;
  assign n5591 = n9975 | n9976;
  assign n9978 = Ng2250 & ~n5142;
  assign n9979 = ~Ng2165 & n5142;
  assign n5596 = n9978 | n9979;
  assign n9981 = Ng2254 & ~n5131_1;
  assign n9982 = Ng2170 & Ng2165;
  assign n9983 = Ng2180 & Ng2175;
  assign n9984 = n9982 & n9983;
  assign n9985 = Ng2195 & Ng2190;
  assign n9986 = n9951 & n9985;
  assign n9987 = n9984 & n9986;
  assign n9988 = n5131_1 & ~n9987;
  assign n5601 = n9981 | n9988;
  assign n9990 = Ng2255 & ~n5138;
  assign n9991 = n5138 & ~n9987;
  assign n5606 = n9990 | n9991;
  assign n9993 = Ng2253 & ~n5142;
  assign n9994 = n5142 & ~n9987;
  assign n5611 = n9993 | n9994;
  assign n9996 = Ng853 & Ng2339;
  assign n9997 = \[1612]  & Ng2333;
  assign n9998 = \[1594]  & Ng2336;
  assign n9999 = ~n9997 & ~n9998;
  assign n10000 = ~n9996 & n9999;
  assign n10001 = Ng853 & Ng2294;
  assign n10002 = \[1612]  & Ng2288;
  assign n10003 = \[1594]  & Ng2291;
  assign n10004 = ~n10002 & ~n10003;
  assign n10005 = ~n10001 & n10004;
  assign n10006 = n10000 & n10005;
  assign n10007 = Ng853 & Ng2285;
  assign n10008 = \[1612]  & Ng2279;
  assign n10009 = \[1594]  & Ng2282;
  assign n10010 = ~n10008 & ~n10009;
  assign n10011 = ~n10007 & n10010;
  assign n10012 = Ng853 & Ng2330;
  assign n10013 = \[1612]  & Ng2324;
  assign n10014 = \[1594]  & Ng2327;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = ~n10012 & n10015;
  assign n10017 = n10011 & n10016;
  assign n10018 = n10006 & n10017;
  assign n10019 = Ng853 & Ng2267;
  assign n10020 = \[1612]  & Ng2261;
  assign n10021 = \[1594]  & Ng2264;
  assign n10022 = ~n10020 & ~n10021;
  assign n10023 = ~n10019 & n10022;
  assign n10024 = Ng853 & ~Ng2395;
  assign n10025 = \[1612]  & ~Ng2393;
  assign n10026 = \[1594]  & ~Ng2394;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = ~n10024 & n10027;
  assign n10029 = Ng853 & ~Ng2389;
  assign n10030 = \[1612]  & ~Ng2387;
  assign n10031 = \[1594]  & ~Ng2388;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = ~n10029 & n10032;
  assign n10034 = n10028 & n10033;
  assign n10035 = n10023 & n10034;
  assign n10036 = n10018 & n10035;
  assign n10037 = Ng853 & ~Ng2392;
  assign n10038 = \[1612]  & ~Ng2390;
  assign n10039 = \[1594]  & ~Ng2391;
  assign n10040 = ~n10038 & ~n10039;
  assign n10041 = ~n10037 & n10040;
  assign n10042 = Ng853 & Ng2276;
  assign n10043 = \[1612]  & Ng2270;
  assign n10044 = \[1594]  & Ng2273;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = ~n10042 & n10045;
  assign n10047 = n10041 & n10046;
  assign n10048 = Ng853 & Ng2348;
  assign n10049 = \[1612]  & Ng2342;
  assign n10050 = \[1594]  & Ng2345;
  assign n10051 = ~n10049 & ~n10050;
  assign n10052 = ~n10048 & n10051;
  assign n10053 = Ng853 & Ng2303;
  assign n10054 = \[1612]  & Ng2297;
  assign n10055 = \[1594]  & Ng2300;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = ~n10053 & n10056;
  assign n10058 = n10052 & n10057;
  assign n10059 = n10047 & n10058;
  assign n10060 = Ng853 & Ng2321;
  assign n10061 = \[1612]  & Ng2315;
  assign n10062 = \[1594]  & Ng2318;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10060 & n10063;
  assign n10065 = Ng853 & Ng2312;
  assign n10066 = \[1612]  & Ng2306;
  assign n10067 = \[1594]  & Ng2309;
  assign n10068 = ~n10066 & ~n10067;
  assign n10069 = ~n10065 & n10068;
  assign n10070 = n10064 & n10069;
  assign n10071 = n10059 & n10070;
  assign n10072 = n10036 & n10071;
  assign n10073 = ~n10033 & n10041;
  assign n10074 = ~n10028 & n10073;
  assign n10075 = n10028 & ~n10033;
  assign n10076 = ~Ng2180 & ~n10064;
  assign n10077 = Ng2180 & n10064;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = ~Ng2170 & ~n10069;
  assign n10080 = Ng2170 & n10069;
  assign n10081 = ~n10079 & ~n10080;
  assign n10082 = n10078 & n10081;
  assign n10083 = ~Ng2190 & ~n10016;
  assign n10084 = Ng2190 & n10016;
  assign n10085 = ~n10083 & ~n10084;
  assign n10086 = ~Ng2200 & ~n10000;
  assign n10087 = Ng2200 & n10000;
  assign n10088 = ~n10086 & ~n10087;
  assign n10089 = n10085 & n10088;
  assign n10090 = ~n10082 & ~n10089;
  assign n10091 = n10078 & n10088;
  assign n10092 = n10090 & ~n10091;
  assign n10093 = ~n9942 & ~n10052;
  assign n10094 = n9942 & n10052;
  assign n10095 = ~n10093 & ~n10094;
  assign n10096 = ~n10092 & ~n10095;
  assign n10097 = Ng853 & ~Ng2244;
  assign n10098 = \[1612]  & ~Ng2245;
  assign n10099 = \[1594]  & ~Ng2246;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = ~n10097 & n10100;
  assign n10102 = Ng2257 & ~n10101;
  assign n10103 = n10090 & n10095;
  assign n10104 = n10078 & n10085;
  assign n10105 = ~n10085 & ~n10088;
  assign n10106 = n10081 & ~n10105;
  assign n10107 = ~n10104 & ~n10106;
  assign n10108 = ~n10103 & ~n10107;
  assign n10109 = n10102 & ~n10108;
  assign n10110 = ~n10096 & n10109;
  assign n10111 = n9928 & ~n10057;
  assign n10112 = ~n9928 & n10057;
  assign n10113 = ~n10111 & ~n10112;
  assign n10114 = ~Ng2185 & ~n10011;
  assign n10115 = Ng2185 & n10011;
  assign n10116 = ~n10114 & ~n10115;
  assign n10117 = ~Ng2195 & ~n10005;
  assign n10118 = Ng2195 & n10005;
  assign n10119 = ~n10117 & ~n10118;
  assign n10120 = n10116 & n10119;
  assign n10121 = ~Ng2175 & ~n10046;
  assign n10122 = Ng2175 & n10046;
  assign n10123 = ~n10121 & ~n10122;
  assign n10124 = ~Ng2165 & ~n10023;
  assign n10125 = Ng2165 & n10023;
  assign n10126 = ~n10124 & ~n10125;
  assign n10127 = n10123 & n10126;
  assign n10128 = ~n10120 & ~n10127;
  assign n10129 = ~n10113 & n10128;
  assign n10130 = n10119 & n10126;
  assign n10131 = n10113 & n10123;
  assign n10132 = ~n10116 & ~n10131;
  assign n10133 = ~n10130 & n10132;
  assign n10134 = n10116 & n10123;
  assign n10135 = n10113 & n10119;
  assign n10136 = ~n10126 & ~n10135;
  assign n10137 = ~n10134 & n10136;
  assign n10138 = ~n10133 & ~n10137;
  assign n10139 = ~n10129 & n10138;
  assign n10140 = n10102 & ~n10139;
  assign n10141 = ~n10110 & ~n10140;
  assign n10142 = n10075 & n10141;
  assign n10143 = ~n10074 & ~n10142;
  assign n10144 = Ng853 & ~Ng2226;
  assign n10145 = \[1612]  & ~Ng2227;
  assign n10146 = \[1594]  & ~Ng2228;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = ~n10144 & n10147;
  assign n10149 = ~Ng2190 & n10148;
  assign n10150 = Ng2190 & ~n10148;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = Ng853 & ~Ng2217;
  assign n10153 = \[1594]  & ~Ng2219;
  assign n10154 = \[1612]  & ~Ng2218;
  assign n10155 = ~n10153 & ~n10154;
  assign n10156 = ~n10152 & n10155;
  assign n10157 = Ng2175 & n10156;
  assign n10158 = n10102 & ~n10157;
  assign n10159 = ~n10151 & n10158;
  assign n10160 = Ng853 & ~Ng2238;
  assign n10161 = \[1612]  & ~Ng2239;
  assign n10162 = \[1594]  & ~Ng2240;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = ~n10160 & n10163;
  assign n10165 = ~n9942 & n10164;
  assign n10166 = n10159 & ~n10165;
  assign n10167 = Ng853 & ~Ng2205;
  assign n10168 = \[1612]  & ~Ng2206;
  assign n10169 = \[1594]  & ~Ng2207;
  assign n10170 = ~n10168 & ~n10169;
  assign n10171 = ~n10167 & n10170;
  assign n10172 = ~Ng2165 & ~n10171;
  assign n10173 = ~Ng2175 & ~n10156;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = Ng853 & ~Ng2223;
  assign n10176 = \[1612]  & ~Ng2224;
  assign n10177 = \[1594]  & ~Ng2225;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10175 & n10178;
  assign n10180 = Ng2185 & n10179;
  assign n10181 = ~Ng2185 & ~n10179;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = n10174 & n10182;
  assign n10184 = Ng853 & ~Ng2208;
  assign n10185 = \[1612]  & ~Ng2209;
  assign n10186 = \[1594]  & ~Ng2210;
  assign n10187 = ~n10185 & ~n10186;
  assign n10188 = ~n10184 & n10187;
  assign n10189 = ~Ng2170 & ~n10188;
  assign n10190 = Ng853 & ~Ng2232;
  assign n10191 = \[1612]  & ~Ng2233;
  assign n10192 = \[1594]  & ~Ng2234;
  assign n10193 = ~n10191 & ~n10192;
  assign n10194 = ~n10190 & n10193;
  assign n10195 = ~Ng2200 & n10194;
  assign n10196 = Ng2200 & ~n10194;
  assign n10197 = ~n10195 & ~n10196;
  assign n10198 = ~n10189 & ~n10197;
  assign n10199 = n10183 & n10198;
  assign n10200 = n10166 & n10199;
  assign n10201 = Ng853 & ~Ng2229;
  assign n10202 = \[1612]  & ~Ng2230;
  assign n10203 = \[1594]  & ~Ng2231;
  assign n10204 = ~n10202 & ~n10203;
  assign n10205 = ~n10201 & n10204;
  assign n10206 = Ng2195 & ~n10205;
  assign n10207 = ~Ng2195 & n10205;
  assign n10208 = ~n10206 & ~n10207;
  assign n10209 = n9942 & ~n10164;
  assign n10210 = Ng853 & ~Ng2235;
  assign n10211 = \[1612]  & ~Ng2236;
  assign n10212 = \[1594]  & ~Ng2237;
  assign n10213 = ~n10211 & ~n10212;
  assign n10214 = ~n10210 & n10213;
  assign n10215 = n9928 & ~n10214;
  assign n10216 = ~n9928 & n10214;
  assign n10217 = ~n10215 & ~n10216;
  assign n10218 = ~n10209 & n10217;
  assign n10219 = ~n10208 & n10218;
  assign n10220 = Ng2165 & n10171;
  assign n10221 = Ng2170 & n10188;
  assign n10222 = ~n10220 & ~n10221;
  assign n10223 = Ng853 & ~Ng2220;
  assign n10224 = \[1612]  & ~Ng2221;
  assign n10225 = \[1594]  & ~Ng2222;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = ~n10223 & n10226;
  assign n10228 = ~Ng2180 & n10227;
  assign n10229 = Ng2180 & ~n10227;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = n10222 & ~n10230;
  assign n10232 = n10219 & n10231;
  assign n10233 = n10200 & n10232;
  assign n10234 = \[1594]  & ~Ng2398;
  assign n10235 = Ng853 & ~Ng2396;
  assign n10236 = \[1612]  & ~Ng2397;
  assign n10237 = ~n10235 & ~n10236;
  assign n10238 = ~n10234 & n10237;
  assign n10239 = n10233 & ~n10238;
  assign n10240 = n10041 & n10239;
  assign n10241 = ~n10143 & n10240;
  assign n10242 = Ng853 & ~Ng2477;
  assign n10243 = \[1612]  & ~Ng2478;
  assign n10244 = \[1594]  & ~Ng2479;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~n10242 & n10245;
  assign n10247 = n10233 & ~n10246;
  assign n10248 = Ng2257 & n10101;
  assign n10249 = ~n10033 & n10248;
  assign n10250 = ~n10247 & ~n10249;
  assign n10251 = ~n10241 & n10250;
  assign n10252 = n10034 & ~n10041;
  assign n10253 = ~n10057 & n10252;
  assign n10254 = n10018 & ~n10052;
  assign n10255 = ~n10046 & ~n10069;
  assign n10256 = ~n10064 & n10255;
  assign n10257 = n10254 & n10256;
  assign n10258 = n10253 & n10257;
  assign n10259 = n10023 & n10258;
  assign n10260 = n10251 & ~n10259;
  assign n10261 = ~n10072 & n10260;
  assign n10262 = ~n10023 & ~n10034;
  assign n10263 = ~n10035 & ~n10262;
  assign n10264 = n10261 & ~n10263;
  assign n10265 = Ng2165 & ~n10251;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = \[1612]  & n10266;
  assign n10268 = ~\[1612]  & ~Ng2261;
  assign n5616 = ~n10267 & ~n10268;
  assign n10270 = \[1594]  & n10266;
  assign n10271 = ~\[1594]  & ~Ng2264;
  assign n5621 = ~n10270 & ~n10271;
  assign n10273 = Ng853 & n10266;
  assign n10274 = ~Ng853 & ~Ng2267;
  assign n5626 = ~n10273 & ~n10274;
  assign n10276 = ~\[1612]  & ~Ng2306;
  assign n10277 = Ng2170 & ~n10251;
  assign n10278 = ~n10260 & ~n10277;
  assign n10279 = n10023 & n10041;
  assign n10280 = ~n10023 & ~n10041;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n10034 & ~n10281;
  assign n10283 = ~n10069 & n10282;
  assign n10284 = n10069 & ~n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = n10261 & ~n10285;
  assign n10287 = ~n10278 & ~n10286;
  assign n10288 = \[1612]  & ~n10287;
  assign n5631 = ~n10276 & ~n10288;
  assign n10290 = ~\[1594]  & ~Ng2309;
  assign n10291 = \[1594]  & ~n10287;
  assign n5636 = ~n10290 & ~n10291;
  assign n10293 = ~Ng853 & ~Ng2312;
  assign n10294 = Ng853 & ~n10287;
  assign n5641 = ~n10293 & ~n10294;
  assign n10296 = ~\[1612]  & ~Ng2270;
  assign n10297 = Ng2175 & ~n10251;
  assign n10298 = ~n10260 & ~n10297;
  assign n10299 = ~n10069 & ~n10280;
  assign n10300 = n10069 & ~n10279;
  assign n10301 = n10034 & ~n10300;
  assign n10302 = ~n10299 & n10301;
  assign n10303 = n10046 & n10302;
  assign n10304 = ~n10046 & ~n10302;
  assign n10305 = ~n10303 & ~n10304;
  assign n10306 = n10261 & n10305;
  assign n10307 = ~n10298 & ~n10306;
  assign n10308 = \[1612]  & ~n10307;
  assign n5646 = ~n10296 & ~n10308;
  assign n10310 = ~\[1594]  & ~Ng2273;
  assign n10311 = \[1594]  & ~n10307;
  assign n5651 = ~n10310 & ~n10311;
  assign n10313 = ~Ng853 & ~Ng2276;
  assign n10314 = Ng853 & ~n10307;
  assign n5656 = ~n10313 & ~n10314;
  assign n10316 = ~\[1612]  & ~Ng2315;
  assign n10317 = Ng2180 & ~n10251;
  assign n10318 = ~n10260 & ~n10317;
  assign n10319 = ~n10041 & ~n10046;
  assign n10320 = ~n10047 & ~n10319;
  assign n10321 = n10302 & ~n10320;
  assign n10322 = ~n10064 & n10321;
  assign n10323 = n10064 & ~n10321;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = n10261 & ~n10324;
  assign n10326 = ~n10318 & ~n10325;
  assign n10327 = \[1612]  & ~n10326;
  assign n5661 = ~n10316 & ~n10327;
  assign n10329 = ~\[1594]  & ~Ng2318;
  assign n10330 = \[1594]  & ~n10326;
  assign n5666 = ~n10329 & ~n10330;
  assign n10332 = ~Ng853 & ~Ng2321;
  assign n10333 = Ng853 & ~n10326;
  assign n5671 = ~n10332 & ~n10333;
  assign n10335 = Ng2185 & ~n10251;
  assign n10336 = ~n10064 & ~n10252;
  assign n10337 = n10064 & n10252;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = n10321 & n10338;
  assign n10340 = n10011 & n10339;
  assign n10341 = ~n10011 & ~n10339;
  assign n10342 = ~n10340 & ~n10341;
  assign n10343 = n10261 & ~n10342;
  assign n10344 = ~n10335 & ~n10343;
  assign n10345 = \[1612]  & n10344;
  assign n10346 = ~\[1612]  & ~Ng2279;
  assign n5676 = ~n10345 & ~n10346;
  assign n10348 = \[1594]  & n10344;
  assign n10349 = ~\[1594]  & ~Ng2282;
  assign n5681 = ~n10348 & ~n10349;
  assign n10351 = Ng853 & n10344;
  assign n10352 = ~Ng853 & ~Ng2285;
  assign n5686 = ~n10351 & ~n10352;
  assign n10354 = ~\[1612]  & Ng2324;
  assign n10355 = Ng2190 & ~n10251;
  assign n10356 = ~n10011 & n10252;
  assign n10357 = n10011 & ~n10252;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = n10339 & ~n10358;
  assign n10360 = n10016 & n10359;
  assign n10361 = ~n10016 & ~n10359;
  assign n10362 = ~n10360 & ~n10361;
  assign n10363 = n10261 & ~n10362;
  assign n10364 = ~n10355 & ~n10363;
  assign n10365 = \[1612]  & ~n10364;
  assign n5691 = n10354 | n10365;
  assign n10367 = ~\[1594]  & Ng2327;
  assign n10368 = \[1594]  & ~n10364;
  assign n5696 = n10367 | n10368;
  assign n10370 = ~Ng853 & Ng2330;
  assign n10371 = Ng853 & ~n10364;
  assign n5701 = n10370 | n10371;
  assign n10373 = Ng2195 & ~n10251;
  assign n10374 = n10016 & n10252;
  assign n10375 = n10322 & n10356;
  assign n10376 = ~n10360 & ~n10375;
  assign n10377 = ~n10374 & ~n10376;
  assign n10378 = n10005 & n10377;
  assign n10379 = ~n10005 & ~n10377;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = n10261 & ~n10380;
  assign n10382 = ~n10373 & ~n10381;
  assign n10383 = \[1612]  & n10382;
  assign n10384 = ~\[1612]  & ~Ng2288;
  assign n5706 = ~n10383 & ~n10384;
  assign n10386 = \[1594]  & n10382;
  assign n10387 = ~\[1594]  & ~Ng2291;
  assign n5711 = ~n10386 & ~n10387;
  assign n10389 = Ng853 & n10382;
  assign n10390 = ~Ng853 & ~Ng2294;
  assign n5716 = ~n10389 & ~n10390;
  assign n10392 = Ng2200 & ~n10251;
  assign n10393 = ~n10005 & n10252;
  assign n10394 = n10005 & ~n10252;
  assign n10395 = ~n10393 & ~n10394;
  assign n10396 = n10377 & ~n10395;
  assign n10397 = n10000 & n10396;
  assign n10398 = ~n10000 & ~n10396;
  assign n10399 = ~n10397 & ~n10398;
  assign n10400 = n10261 & ~n10399;
  assign n10401 = ~n10392 & ~n10400;
  assign n10402 = \[1612]  & n10401;
  assign n10403 = ~\[1612]  & ~Ng2333;
  assign n5721 = ~n10402 & ~n10403;
  assign n10405 = \[1594]  & n10401;
  assign n10406 = ~\[1594]  & ~Ng2336;
  assign n5726 = ~n10405 & ~n10406;
  assign n10408 = Ng853 & n10401;
  assign n10409 = ~Ng853 & ~Ng2339;
  assign n5731 = ~n10408 & ~n10409;
  assign n10411 = ~\[1612]  & ~Ng2297;
  assign n10412 = ~n9928 & ~n10251;
  assign n10413 = ~n10260 & ~n10412;
  assign n10414 = ~n10000 & ~n10016;
  assign n10415 = ~n10006 & ~n10414;
  assign n10416 = ~n10395 & ~n10415;
  assign n10417 = ~n10376 & n10416;
  assign n10418 = ~n10057 & n10417;
  assign n10419 = n10057 & ~n10417;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = n10261 & ~n10420;
  assign n10422 = ~n10413 & ~n10421;
  assign n10423 = \[1612]  & ~n10422;
  assign n5736 = ~n10411 & ~n10423;
  assign n10425 = ~\[1594]  & ~Ng2300;
  assign n10426 = \[1594]  & ~n10422;
  assign n5741 = ~n10425 & ~n10426;
  assign n10428 = ~Ng853 & ~Ng2303;
  assign n10429 = Ng853 & ~n10422;
  assign n5746 = ~n10428 & ~n10429;
  assign n10431 = ~\[1612]  & ~Ng2342;
  assign n10432 = ~n9942 & ~n10251;
  assign n10433 = ~n10260 & ~n10432;
  assign n10434 = n10057 & ~n10252;
  assign n10435 = ~n10253 & ~n10434;
  assign n10436 = n10417 & ~n10435;
  assign n10437 = n10052 & n10436;
  assign n10438 = ~n10052 & ~n10436;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = n10261 & n10439;
  assign n10441 = ~n10433 & ~n10440;
  assign n10442 = \[1612]  & ~n10441;
  assign n5751 = ~n10431 & ~n10442;
  assign n10444 = ~\[1594]  & ~Ng2345;
  assign n10445 = \[1594]  & ~n10441;
  assign n5756 = ~n10444 & ~n10445;
  assign n10447 = ~Ng853 & ~Ng2348;
  assign n10448 = Ng853 & ~n10441;
  assign n5761 = ~n10447 & ~n10448;
  assign n10450 = Ng2160 & n5635;
  assign n10451 = Ng2160 & ~n5027;
  assign n10452 = ~n5635 & ~n10451;
  assign n5766 = ~n10450 & ~n10452;
  assign n10454 = Ng2156 & n10450;
  assign n10455 = ~Ng2156 & ~n10450;
  assign n10456 = ~n5642 & ~n10455;
  assign n5771 = ~n10454 & n10456;
  assign n10458 = Ng2151 & n10454;
  assign n10459 = ~Ng2151 & ~n10454;
  assign n10460 = ~n5642 & ~n10459;
  assign n5776 = ~n10458 & n10460;
  assign n10462 = Ng2147 & n10458;
  assign n10463 = ~Ng2147 & ~n10458;
  assign n10464 = ~n5642 & ~n10463;
  assign n5781 = ~n10462 & n10464;
  assign n10466 = Ng2142 & n10462;
  assign n10467 = ~Ng2142 & ~n10462;
  assign n10468 = ~n5642 & ~n10467;
  assign n5786 = ~n10466 & n10468;
  assign n10470 = Ng2138 & n10466;
  assign n10471 = ~Ng2138 & ~n10466;
  assign n10472 = ~n5642 & ~n10471;
  assign n5791 = ~n10470 & n10472;
  assign n10474 = Ng2133 & n10470;
  assign n10475 = ~Ng2133 & ~n10470;
  assign n10476 = ~n5642 & ~n10475;
  assign n5796 = ~n10474 & n10476;
  assign n10478 = Ng2129 & n10474;
  assign n10479 = ~Ng2129 & ~n10474;
  assign n10480 = ~n5642 & ~n10479;
  assign n5801 = ~n10478 & n10480;
  assign n10482 = Ng2124 & n10478;
  assign n10483 = ~Ng2124 & ~n10478;
  assign n10484 = ~n5642 & ~n10483;
  assign n5806 = ~n10482 & n10484;
  assign n10486 = Ng2120 & n10482;
  assign n10487 = ~Ng2120 & ~n10482;
  assign n10488 = ~n10486 & ~n10487;
  assign n5811 = ~n5642 & n10488;
  assign n10490 = n10034 & n10041;
  assign n10491 = n10033 & ~n10041;
  assign n10492 = ~n10028 & n10491;
  assign n10493 = ~n5124 & ~n10492;
  assign n10494 = ~n10490 & ~n10493;
  assign n10495 = \[1612]  & ~n10494;
  assign n10496 = Ng853 & ~Ng11580;
  assign n10497 = \[1612]  & ~Ng11578;
  assign n10498 = \[1594]  & ~Ng11579;
  assign n10499 = ~n10497 & ~n10498;
  assign n10500 = ~n10496 & n10499;
  assign n10501 = Ng853 & ~Ng11586;
  assign n10502 = \[1612]  & ~Ng11584;
  assign n10503 = \[1594]  & ~Ng11585;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = ~n10501 & n10504;
  assign n10506 = Ng853 & ~Ng11583;
  assign n10507 = \[1612]  & ~Ng11581;
  assign n10508 = \[1594]  & ~Ng11582;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n10506 & n10509;
  assign n10511 = n10505 & ~n10510;
  assign n10512 = Ng853 & ~Ng11589;
  assign n10513 = \[1612]  & ~Ng11587;
  assign n10514 = \[1594]  & ~Ng11588;
  assign n10515 = ~n10513 & ~n10514;
  assign n10516 = ~n10512 & n10515;
  assign n10517 = ~n10511 & n10516;
  assign n10518 = ~n10500 & n10517;
  assign n10519 = ~Pg3229 & n10511;
  assign n10520 = Pg3229 & ~n10516;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = ~n10518 & n10521;
  assign n10523 = n10495 & ~n10522;
  assign n10524 = ~Ng11578 & ~n10495;
  assign n5829 = ~n10523 & ~n10524;
  assign n10526 = \[1594]  & ~n10494;
  assign n10527 = ~n10522 & n10526;
  assign n10528 = ~Ng11579 & ~n10526;
  assign n5834 = ~n10527 & ~n10528;
  assign n10530 = Ng853 & ~n10494;
  assign n10531 = ~n10522 & n10530;
  assign n10532 = ~Ng11580 & ~n10530;
  assign n5839 = ~n10531 & ~n10532;
  assign n10534 = ~Pg3229 & ~n10500;
  assign n10535 = Pg3229 & n10500;
  assign n10536 = ~n10534 & ~n10535;
  assign n10537 = ~n10505 & n10536;
  assign n10538 = ~n10511 & ~n10537;
  assign n10539 = n10495 & ~n10538;
  assign n10540 = ~Ng11581 & ~n10495;
  assign n5844 = ~n10539 & ~n10540;
  assign n10542 = n10526 & n10538;
  assign n10543 = Ng11582 & ~n10526;
  assign n5849 = n10542 | n10543;
  assign n10545 = ~Ng11583 & ~n10530;
  assign n10546 = n10530 & ~n10538;
  assign n5854 = ~n10545 & ~n10546;
  assign n10548 = n10510 & n10516;
  assign n10549 = n10536 & ~n10548;
  assign n10550 = n10510 & ~n10536;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = n10495 & n10551;
  assign n10553 = ~Ng11584 & ~n10495;
  assign n5859 = ~n10552 & ~n10553;
  assign n10555 = n10526 & ~n10551;
  assign n10556 = Ng11585 & ~n10526;
  assign n5864 = n10555 | n10556;
  assign n10558 = n10530 & n10551;
  assign n10559 = ~Ng11586 & ~n10530;
  assign n5869 = ~n10558 & ~n10559;
  assign n10561 = n10505 & n10550;
  assign n10562 = n10495 & ~n10561;
  assign n10563 = Ng11587 & ~n10495;
  assign n5874 = n10562 | n10563;
  assign n10565 = n10526 & ~n10561;
  assign n10566 = Ng11588 & ~n10526;
  assign n5879 = n10565 | n10566;
  assign n10568 = n10530 & ~n10561;
  assign n10569 = Ng11589 & ~n10530;
  assign n5884 = n10568 | n10569;
  assign n10571 = ~n9942 & n9987;
  assign n10572 = ~n9928 & n10571;
  assign n10573 = Ng853 & Ng2498;
  assign n10574 = \[1612]  & Ng2492;
  assign n10575 = \[1594]  & Ng2495;
  assign n10576 = ~n10574 & ~n10575;
  assign n6134 = n10573 | ~n10576;
  assign n10578 = ~n10248 & ~n6134;
  assign n10579 = n10572 & n10578;
  assign n10580 = ~n10572 & n6134;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = Ng853 & Ng2489;
  assign n10583 = \[1612]  & Ng2483;
  assign n10584 = \[1594]  & Ng2486;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = ~n10582 & n10585;
  assign n10587 = Ng2257 & n10586;
  assign n10588 = ~n10581 & n10587;
  assign n10589 = Ng853 & ~Ng2501;
  assign n10590 = \[1612]  & ~Ng2502;
  assign n10591 = \[1594]  & ~Ng2503;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = ~n10589 & n10592;
  assign n10594 = ~n10581 & n10593;
  assign n10595 = Ng2257 & ~n10594;
  assign n10596 = ~n10586 & ~n10595;
  assign n10597 = ~n10588 & ~n10596;
  assign n10598 = \[1612]  & n10597;
  assign n10599 = ~\[1612]  & ~Ng2483;
  assign n5889 = ~n10598 & ~n10599;
  assign n10601 = \[1594]  & n10597;
  assign n10602 = ~\[1594]  & ~Ng2486;
  assign n5894 = ~n10601 & ~n10602;
  assign n10604 = Ng853 & n10597;
  assign n10605 = ~Ng853 & ~Ng2489;
  assign n5899 = ~n10604 & ~n10605;
  assign n10607 = ~\[1612]  & Ng2492;
  assign n10608 = Ng2257 & ~n10586;
  assign n10609 = ~n10593 & n10608;
  assign n10610 = n6134 & ~n10609;
  assign n10611 = ~n10248 & ~n10609;
  assign n10612 = n10572 & ~n10611;
  assign n10613 = ~n10610 & ~n10612;
  assign n10614 = \[1612]  & ~n10613;
  assign n5904 = n10607 | n10614;
  assign n10616 = ~\[1594]  & Ng2495;
  assign n10617 = \[1594]  & ~n10613;
  assign n5909 = n10616 | n10617;
  assign n10619 = ~Ng853 & Ng2498;
  assign n10620 = Ng853 & ~n10613;
  assign n5914 = n10619 | n10620;
  assign n10622 = n10594 & n10608;
  assign n10623 = \[1612]  & n10622;
  assign n10624 = \[1612]  & n10588;
  assign n10625 = ~Ng2502 & ~n10624;
  assign n5919 = ~n10623 & ~n10625;
  assign n10627 = \[1594]  & n10622;
  assign n10628 = \[1594]  & n10588;
  assign n10629 = ~Ng2503 & ~n10628;
  assign n5924 = ~n10627 & ~n10629;
  assign n10631 = Ng853 & n10622;
  assign n10632 = Ng853 & n10588;
  assign n10633 = ~Ng2501 & ~n10632;
  assign n5929 = ~n10631 & ~n10633;
  assign n10635 = ~\[1612]  & Ng2504;
  assign n10636 = Ng853 & ~Ng2253;
  assign n10637 = \[1612]  & ~Ng2254;
  assign n10638 = \[1594]  & ~Ng2255;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = ~n10636 & n10639;
  assign n10641 = n9987 & ~n10640;
  assign n10642 = Ng2257 & n10641;
  assign n10643 = Ng853 & Ng2510;
  assign n10644 = \[1612]  & Ng2504;
  assign n10645 = \[1594]  & Ng2507;
  assign n10646 = ~n10644 & ~n10645;
  assign n10647 = ~n10643 & n10646;
  assign n10648 = ~Ng2257 & ~n10647;
  assign n10649 = ~n10642 & ~n10648;
  assign n10650 = \[1612]  & ~n10649;
  assign n5934 = n10635 | n10650;
  assign n10652 = ~\[1594]  & Ng2507;
  assign n10653 = \[1594]  & ~n10649;
  assign n5939 = n10652 | n10653;
  assign n10655 = ~Ng853 & Ng2510;
  assign n10656 = Ng853 & ~n10649;
  assign n5944 = n10655 | n10656;
  assign n10658 = ~\[1612]  & ~Ng2513;
  assign n10659 = Ng853 & Ng2519;
  assign n10660 = \[1612]  & Ng2513;
  assign n10661 = \[1594]  & Ng2516;
  assign n10662 = ~n10660 & ~n10661;
  assign n10663 = ~n10659 & n10662;
  assign n10664 = Ng853 & ~Ng2522;
  assign n10665 = \[1612]  & ~Ng2523;
  assign n10666 = \[1594]  & ~Ng2524;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = ~n10664 & n10667;
  assign n10669 = n10641 & n10663;
  assign n10670 = ~n10647 & ~n10669;
  assign n10671 = ~n10641 & ~n10663;
  assign n10672 = n10647 & ~n10671;
  assign n10673 = Ng2257 & ~n10672;
  assign n10674 = ~n10670 & n10673;
  assign n10675 = ~n10668 & n10674;
  assign n10676 = n10663 & n10675;
  assign n10677 = ~n10663 & ~n10675;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = \[1612]  & n10678;
  assign n5949 = ~n10658 & ~n10679;
  assign n10681 = ~\[1594]  & ~Ng2516;
  assign n10682 = \[1594]  & n10678;
  assign n5954 = ~n10681 & ~n10682;
  assign n10684 = ~Ng853 & ~Ng2519;
  assign n10685 = Ng853 & n10678;
  assign n5959 = ~n10684 & ~n10685;
  assign n10687 = n10668 & n10674;
  assign n10688 = \[1612]  & n10687;
  assign n10689 = n10647 & ~n10669;
  assign n10690 = ~n10647 & ~n10671;
  assign n10691 = Ng2257 & ~n10690;
  assign n10692 = ~n10689 & n10691;
  assign n10693 = \[1612]  & n10692;
  assign n10694 = ~Ng2523 & ~n10693;
  assign n5964 = ~n10688 & ~n10694;
  assign n10696 = \[1594]  & n10687;
  assign n10697 = \[1594]  & n10692;
  assign n10698 = ~Ng2524 & ~n10697;
  assign n5969 = ~n10696 & ~n10698;
  assign n10700 = Ng853 & n10687;
  assign n10701 = Ng853 & n10692;
  assign n10702 = ~Ng2522 & ~n10701;
  assign n5974 = ~n10700 & ~n10702;
  assign n10704 = ~\[1612]  & ~Ng2387;
  assign n10705 = ~n10033 & ~n10041;
  assign n10706 = ~n10075 & ~n10705;
  assign n10707 = ~n10141 & ~n10706;
  assign n10708 = ~n10252 & ~n10707;
  assign n10709 = ~n10247 & ~n10708;
  assign n10710 = \[1612]  & ~n10709;
  assign n5979 = ~n10704 & ~n10710;
  assign n10712 = ~\[1594]  & ~Ng2388;
  assign n10713 = \[1594]  & ~n10709;
  assign n5984 = ~n10712 & ~n10713;
  assign n10715 = ~Ng853 & ~Ng2389;
  assign n10716 = Ng853 & ~n10709;
  assign n5989 = ~n10715 & ~n10716;
  assign n10718 = ~\[1612]  & ~Ng2390;
  assign n10719 = n10141 & n10239;
  assign n10720 = n10028 & ~n10110;
  assign n10721 = ~n10095 & n10113;
  assign n10722 = n10120 & n10721;
  assign n10723 = n10089 & n10722;
  assign n10724 = n10127 & n10723;
  assign n10725 = n10082 & n10724;
  assign n10726 = ~n10101 & ~n10725;
  assign n10727 = Ng2257 & ~n10726;
  assign n10728 = n10720 & ~n10727;
  assign n10729 = ~n10239 & ~n10248;
  assign n10730 = ~n10028 & n10729;
  assign n10731 = ~n10728 & ~n10730;
  assign n10732 = ~n10719 & ~n10731;
  assign n10733 = n10073 & ~n10732;
  assign n10734 = n10102 & ~n10725;
  assign n10735 = n10720 & n10734;
  assign n10736 = ~n10041 & ~n10140;
  assign n10737 = ~n10735 & n10736;
  assign n10738 = ~n10034 & ~n10247;
  assign n10739 = ~n10491 & n10738;
  assign n10740 = ~n10737 & n10739;
  assign n10741 = ~n10733 & n10740;
  assign n10742 = \[1612]  & ~n10741;
  assign n5994 = ~n10718 & ~n10742;
  assign n10744 = ~\[1594]  & ~Ng2391;
  assign n10745 = \[1594]  & ~n10741;
  assign n5999 = ~n10744 & ~n10745;
  assign n10747 = ~Ng853 & ~Ng2392;
  assign n10748 = Ng853 & ~n10741;
  assign n6004 = ~n10747 & ~n10748;
  assign n10750 = ~\[1612]  & ~Ng2393;
  assign n10751 = ~n10041 & n10727;
  assign n10752 = Ng2257 & n10041;
  assign n10753 = n10141 & n10752;
  assign n10754 = n10075 & ~n10753;
  assign n10755 = ~n10751 & n10754;
  assign n10756 = ~n10028 & n10734;
  assign n10757 = n10705 & n10756;
  assign n10758 = ~n10755 & ~n10757;
  assign n10759 = ~n10247 & ~n10758;
  assign n10760 = \[1612]  & ~n10759;
  assign n6009 = ~n10750 & ~n10760;
  assign n10762 = ~\[1594]  & ~Ng2394;
  assign n10763 = \[1594]  & ~n10759;
  assign n6014 = ~n10762 & ~n10763;
  assign n10765 = ~Ng853 & ~Ng2395;
  assign n10766 = Ng853 & ~n10759;
  assign n6019 = ~n10765 & ~n10766;
  assign n10768 = ~n10074 & ~n10726;
  assign n10769 = n5019_1 & ~n10768;
  assign n10770 = Ng2397 & ~n10769;
  assign n10771 = ~n10143 & n10233;
  assign n10772 = n10769 & ~n10771;
  assign n6024 = n10770 | n10772;
  assign n10774 = n5023 & ~n10768;
  assign n10775 = n10771 & n10774;
  assign n10776 = ~Ng2398 & ~n10774;
  assign n6029 = ~n10775 & ~n10776;
  assign n10778 = n5027 & ~n10768;
  assign n10779 = Ng2396 & ~n10778;
  assign n10780 = ~n10771 & n10778;
  assign n6034 = n10779 | n10780;
  assign n10782 = n10233 & n10246;
  assign n10783 = n5019_1 & ~n10782;
  assign n10784 = Ng2478 & ~n5019_1;
  assign n6039 = n10783 | n10784;
  assign n10786 = n5023 & ~n10782;
  assign n10787 = Ng2479 & ~n5023;
  assign n6044 = n10786 | n10787;
  assign n10789 = n5027 & ~n10782;
  assign n10790 = Ng2477 & ~n5027;
  assign n6049 = n10789 | n10790;
  assign n10792 = ~Ng2374 & Ng2373;
  assign n10793 = ~\[1594]  & Ng2380;
  assign n10794 = \[1594]  & n4632;
  assign n10795 = Ng2374 & ~n10794;
  assign n10796 = ~n10793 & n10795;
  assign n6139 = ~n10792 & ~n10796;
  assign n10798 = ~Ng2138 & n10016;
  assign n10799 = Ng2138 & ~n10016;
  assign n10800 = ~n10798 & ~n10799;
  assign n10801 = Ng2151 & ~n10046;
  assign n10802 = ~Ng2151 & n10046;
  assign n10803 = ~n10801 & ~n10802;
  assign n10804 = ~Ng2129 & ~n10000;
  assign n10805 = ~Ng2120 & ~n10052;
  assign n10806 = ~n10804 & ~n10805;
  assign n10807 = Ng2133 & n10005;
  assign n10808 = n10806 & ~n10807;
  assign n10809 = ~n10803 & n10808;
  assign n10810 = ~n10800 & n10809;
  assign n10811 = ~Ng2124 & ~n10057;
  assign n10812 = Ng2142 & n10011;
  assign n10813 = ~n10811 & ~n10812;
  assign n10814 = ~Ng2156 & ~n10069;
  assign n10815 = Ng2156 & n10069;
  assign n10816 = ~n10814 & ~n10815;
  assign n10817 = ~Ng2142 & ~n10011;
  assign n10818 = Ng2120 & n10052;
  assign n10819 = ~n10817 & ~n10818;
  assign n10820 = n10816 & n10819;
  assign n10821 = Ng2124 & n10057;
  assign n10822 = ~Ng2133 & ~n10005;
  assign n10823 = ~n10821 & ~n10822;
  assign n10824 = Ng2160 & n10023;
  assign n10825 = n10823 & ~n10824;
  assign n10826 = n10820 & n10825;
  assign n10827 = n10813 & n10826;
  assign n10828 = ~Ng2160 & ~n10023;
  assign n10829 = Ng2129 & n10000;
  assign n10830 = ~n10828 & ~n10829;
  assign n10831 = n10493 & n10830;
  assign n10832 = ~Ng2147 & n10064;
  assign n10833 = Ng2147 & ~n10064;
  assign n10834 = ~n10832 & ~n10833;
  assign n10835 = n10831 & ~n10834;
  assign n10836 = n10827 & n10835;
  assign n10837 = n10810 & n10836;
  assign n6144 = ~n10072 & ~n10837;
  assign n10839 = ~Ng1315 & Ng2628;
  assign n6245 = n6033 | n10839;
  assign n10841 = Ng1315 & Ng2628;
  assign n10842 = ~Ng1315 & ~Ng2631;
  assign n6250 = ~n10841 & ~n10842;
  assign n10844 = Ng1315 & Ng2631;
  assign n10845 = ~Ng1315 & Ng2584;
  assign n6255 = n10844 | n10845;
  assign n10847 = Ng1315 & Ng2647;
  assign n10848 = \[1605]  & Ng2643;
  assign n10849 = \[1603]  & Ng2645;
  assign n10850 = ~n10848 & ~n10849;
  assign n6260 = ~n10847 & n10850;
  assign n10852 = ~\[1612]  & Ng2561;
  assign n10853 = \[1612]  & ~n10663;
  assign n6327 = n10852 | n10853;
  assign n10855 = ~\[1594]  & Ng2562;
  assign n10856 = \[1594]  & ~n10663;
  assign n6332 = n10855 | n10856;
  assign n10858 = ~Ng853 & Ng2563;
  assign n10859 = Ng853 & ~n10663;
  assign n6337 = n10858 | n10859;
  assign n10861 = ~\[1612]  & ~Ng11593;
  assign n10862 = \[1612]  & ~n10492;
  assign n6342 = ~n10861 & ~n10862;
  assign n10864 = ~\[1594]  & ~Ng11596;
  assign n10865 = \[1594]  & ~n10492;
  assign n6346 = ~n10864 & ~n10865;
  assign n10867 = ~Ng853 & ~Ng11597;
  assign n10868 = Ng853 & ~n10492;
  assign n6350 = ~n10867 & ~n10868;
  assign n10870 = ~\[1612]  & ~Ng2552;
  assign n10871 = \[1612]  & ~n10074;
  assign n6354 = ~n10870 & ~n10871;
  assign n10873 = ~\[1594]  & ~Ng2553;
  assign n10874 = \[1594]  & ~n10074;
  assign n6359 = ~n10873 & ~n10874;
  assign n10876 = ~Ng853 & ~Ng2554;
  assign n10877 = Ng853 & ~n10074;
  assign n6364 = ~n10876 & ~n10877;
  assign n10879 = ~\[1612]  & ~Ng2555;
  assign n10880 = \[1612]  & n6134;
  assign n6369 = ~n10879 & ~n10880;
  assign n10882 = ~\[1594]  & ~Ng2559;
  assign n10883 = \[1594]  & n6134;
  assign n6374 = ~n10882 & ~n10883;
  assign n10885 = ~Ng853 & ~Ng2539;
  assign n10886 = Ng853 & n6134;
  assign n6379 = ~n10885 & ~n10886;
  assign n10888 = ~\[1612]  & ~Ng11598;
  assign n10889 = \[1612]  & ~n10490;
  assign n6384 = ~n10888 & ~n10889;
  assign n10891 = ~\[1594]  & ~Ng11594;
  assign n10892 = \[1594]  & ~n10490;
  assign n6388 = ~n10891 & ~n10892;
  assign n10894 = ~Ng853 & ~Ng11595;
  assign n10895 = Ng853 & ~n10490;
  assign n6392 = ~n10894 & ~n10895;
  assign n10897 = Ng1315 & Ng2564;
  assign n10898 = \[1605]  & Ng2639;
  assign n10899 = \[1603]  & Ng2641;
  assign n10900 = ~n10898 & ~n10899;
  assign n6396 = ~n10897 & n10900;
  assign n10902 = \[1605]  & ~Ng2554;
  assign n10903 = \[1603]  & ~Ng2552;
  assign n10904 = Ng1315 & ~Ng2553;
  assign n10905 = ~n10903 & ~n10904;
  assign n6409 = ~n10902 & n10905;
  assign n10907 = \[1605]  & ~Ng2539;
  assign n10908 = \[1603]  & ~Ng2555;
  assign n10909 = Ng1315 & ~Ng2559;
  assign n10910 = ~n10908 & ~n10909;
  assign n6423 = ~n10907 & n10910;
  assign n10912 = \[1605]  & ~Ng2563;
  assign n10913 = \[1603]  & ~Ng2561;
  assign n10914 = Ng1315 & ~Ng2562;
  assign n10915 = ~n10913 & ~n10914;
  assign n6432 = ~n10912 & n10915;
  assign n10917 = Ng1315 & Ng2694;
  assign n10918 = \[1605]  & Ng2688;
  assign n10919 = \[1603]  & Ng2691;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = ~n10917 & n10920;
  assign n10922 = Ng1315 & Ng2571;
  assign n10923 = \[1605]  & Ng2565;
  assign n10924 = \[1603]  & Ng2568;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926 = ~n10922 & n10925;
  assign n10927 = Ng2584 & n10926;
  assign n10928 = ~n10921 & n10927;
  assign n10929 = Ng1315 & Ng2685;
  assign n10930 = \[1605]  & Ng2679;
  assign n10931 = \[1603]  & Ng2682;
  assign n10932 = ~n10930 & ~n10931;
  assign n10933 = ~n10929 & n10932;
  assign n10934 = ~n10926 & ~n10933;
  assign n10935 = ~n6126 & ~n10934;
  assign n6580 = n10928 | n10935;
  assign n10937 = \[1605]  & n6580;
  assign n10938 = ~Ng2650 & ~n10937;
  assign n10939 = Ng1315 & ~Ng2658;
  assign n10940 = \[1605]  & ~Ng2659;
  assign n10941 = \[1603]  & ~Ng2660;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = ~n10939 & n10942;
  assign n10944 = Pg3229 & ~n10943;
  assign n10945 = Ng1315 & ~Ng2655;
  assign n10946 = \[1605]  & ~Ng2656;
  assign n10947 = \[1603]  & ~Ng2657;
  assign n10948 = ~n10946 & ~n10947;
  assign n10949 = ~n10945 & n10948;
  assign n10950 = Ng1315 & ~Ng2652;
  assign n10951 = \[1605]  & ~Ng2653;
  assign n10952 = \[1603]  & ~Ng2654;
  assign n10953 = ~n10951 & ~n10952;
  assign n10954 = ~n10950 & n10953;
  assign n10955 = n10949 & ~n10954;
  assign n10956 = Ng1315 & ~Ng2649;
  assign n10957 = \[1605]  & ~Ng2650;
  assign n10958 = \[1603]  & ~Ng2651;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = ~n10956 & n10959;
  assign n10961 = n10943 & ~n10960;
  assign n10962 = ~n10955 & n10961;
  assign n10963 = ~Pg3229 & n10955;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~n10944 & n10964;
  assign n10966 = n10937 & ~n10965;
  assign n6441 = ~n10938 & ~n10966;
  assign n10968 = \[1603]  & n6580;
  assign n10969 = ~n10965 & n10968;
  assign n10970 = ~Ng2651 & ~n10968;
  assign n6446 = ~n10969 & ~n10970;
  assign n10972 = Ng1315 & n6580;
  assign n10973 = ~n10965 & n10972;
  assign n10974 = ~Ng2649 & ~n10972;
  assign n6451 = ~n10973 & ~n10974;
  assign n10976 = ~Pg3229 & ~n10960;
  assign n10977 = Pg3229 & n10960;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~n10949 & n10978;
  assign n10980 = ~n10955 & ~n10979;
  assign n10981 = n10937 & n10980;
  assign n10982 = Ng2653 & ~n10937;
  assign n6456 = n10981 | n10982;
  assign n10984 = n10968 & n10980;
  assign n10985 = Ng2654 & ~n10968;
  assign n6461 = n10984 | n10985;
  assign n10987 = n10972 & n10980;
  assign n10988 = Ng2652 & ~n10972;
  assign n6466 = n10987 | n10988;
  assign n10990 = n10943 & n10954;
  assign n10991 = n10978 & ~n10990;
  assign n10992 = n10954 & ~n10978;
  assign n10993 = ~n10991 & ~n10992;
  assign n10994 = n10937 & ~n10993;
  assign n10995 = Ng2656 & ~n10937;
  assign n6471 = n10994 | n10995;
  assign n10997 = n10968 & ~n10993;
  assign n10998 = Ng2657 & ~n10968;
  assign n6476 = n10997 | n10998;
  assign n11000 = n10972 & ~n10993;
  assign n11001 = Ng2655 & ~n10972;
  assign n6481 = n11000 | n11001;
  assign n11003 = n10949 & n10954;
  assign n11004 = ~n10978 & n11003;
  assign n11005 = n10937 & ~n11004;
  assign n11006 = Ng2659 & ~n10937;
  assign n6486 = n11005 | n11006;
  assign n11008 = n10968 & ~n11004;
  assign n11009 = Ng2660 & ~n10968;
  assign n6491 = n11008 | n11009;
  assign n11011 = n10972 & ~n11004;
  assign n11012 = Ng2658 & ~n10972;
  assign n6496 = n11011 | n11012;
  assign n11014 = ~\[1605]  & ~Ng2661;
  assign n11015 = Ng185 & Ng2598;
  assign n11016 = ~n6260 & n11015;
  assign n11017 = \[1603]  & Ng2664;
  assign n11018 = Ng1315 & Ng2667;
  assign n11019 = \[1605]  & Ng2661;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n11017 & n11020;
  assign n11022 = ~n11016 & n11021;
  assign n11023 = ~n6032 & ~n11022;
  assign n11024 = \[1605]  & ~n11023;
  assign n6501 = ~n11014 & ~n11024;
  assign n11026 = ~\[1603]  & ~Ng2664;
  assign n11027 = \[1603]  & ~n11023;
  assign n6506 = ~n11026 & ~n11027;
  assign n11029 = ~Ng1315 & Ng2667;
  assign n11030 = n6033 & ~n11022;
  assign n6511 = n11029 | n11030;
  assign n11032 = ~\[1605]  & ~Ng2670;
  assign n11033 = Ng185 & Ng2616;
  assign n11034 = ~n6396 & n11033;
  assign n11035 = Ng1315 & Ng2676;
  assign n11036 = \[1603]  & Ng2673;
  assign n11037 = \[1605]  & Ng2670;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = ~n11035 & n11038;
  assign n11040 = ~n11034 & n11039;
  assign n11041 = ~n6032 & ~n11040;
  assign n11042 = \[1605]  & ~n11041;
  assign n6516 = ~n11032 & ~n11042;
  assign n11044 = ~\[1603]  & ~Ng2673;
  assign n11045 = \[1603]  & ~n11041;
  assign n6521 = ~n11044 & ~n11045;
  assign n11047 = ~Ng1315 & Ng2676;
  assign n11048 = n6033 & ~n11040;
  assign n6526 = n11047 | n11048;
  assign n11050 = ~\[1605]  & Ng2688;
  assign n11051 = ~n6032 & ~n10921;
  assign n11052 = ~n11022 & ~n11040;
  assign n11053 = n6032 & ~n11052;
  assign n11054 = Ng1315 & Ng2443;
  assign n11055 = \[1605]  & Ng2439;
  assign n11056 = \[1603]  & Ng2441;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = ~n11054 & n11057;
  assign n11059 = Ng1315 & Ng2428;
  assign n11060 = \[1605]  & Ng2424;
  assign n11061 = \[1603]  & Ng2426;
  assign n11062 = ~n11060 & ~n11061;
  assign n11063 = ~n11059 & n11062;
  assign n11064 = n10949 & n11063;
  assign n11065 = Ng1315 & Ng2458;
  assign n11066 = \[1605]  & Ng2454;
  assign n11067 = \[1603]  & Ng2456;
  assign n11068 = ~n11066 & ~n11067;
  assign n11069 = ~n11065 & n11068;
  assign n11070 = n10960 & ~n11069;
  assign n11071 = ~n11064 & ~n11070;
  assign n11072 = n11058 & ~n11071;
  assign n11073 = ~n10954 & n11072;
  assign n11074 = ~n11058 & ~n11069;
  assign n11075 = ~n10943 & n11074;
  assign n11076 = ~n10949 & n11058;
  assign n11077 = n10990 & n11069;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = Ng1315 & Ng2399;
  assign n11080 = \[1605]  & Ng2469;
  assign n11081 = \[1603]  & Ng2471;
  assign n11082 = ~n11080 & ~n11081;
  assign n11083 = ~n11079 & n11082;
  assign n11084 = ~n11058 & ~n11083;
  assign n11085 = n10949 & n11084;
  assign n11086 = n10954 & n11085;
  assign n11087 = n11078 & ~n11086;
  assign n11088 = n10960 & ~n11087;
  assign n11089 = ~n11075 & ~n11088;
  assign n11090 = ~n11063 & ~n11089;
  assign n11091 = n11003 & n11083;
  assign n11092 = n10990 & n11074;
  assign n11093 = ~n10949 & n11084;
  assign n11094 = ~n10954 & n11069;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = ~n11092 & n11095;
  assign n11097 = n11063 & ~n11096;
  assign n11098 = ~n11091 & ~n11097;
  assign n11099 = ~n10960 & ~n11098;
  assign n11100 = ~n11090 & ~n11099;
  assign n11101 = ~n11073 & n11100;
  assign n11102 = n10943 & ~n11063;
  assign n11103 = n10949 & ~n11102;
  assign n11104 = n11083 & ~n11103;
  assign n11105 = n10949 & ~n11063;
  assign n11106 = ~n10954 & n11063;
  assign n11107 = ~n11105 & ~n11106;
  assign n11108 = n11074 & n11107;
  assign n11109 = ~n11104 & ~n11108;
  assign n11110 = n10960 & ~n11109;
  assign n11111 = n11003 & ~n11058;
  assign n11112 = n10943 & ~n11111;
  assign n11113 = ~n10943 & ~n11083;
  assign n11114 = ~n11069 & ~n11113;
  assign n11115 = ~n11070 & ~n11114;
  assign n11116 = n11063 & n11115;
  assign n11117 = ~n11112 & n11116;
  assign n11118 = ~n11110 & ~n11117;
  assign n11119 = n11069 & ~n11076;
  assign n11120 = ~n11085 & ~n11119;
  assign n11121 = ~n10954 & ~n11120;
  assign n11122 = ~n11063 & n11121;
  assign n11123 = ~n11069 & ~n11103;
  assign n11124 = ~n11107 & ~n11123;
  assign n11125 = ~n10960 & n11058;
  assign n11126 = ~n11124 & n11125;
  assign n11127 = ~n11122 & ~n11126;
  assign n11128 = n11118 & n11127;
  assign n11129 = n11040 & n11128;
  assign n11130 = n11101 & ~n11129;
  assign n11131 = n11053 & n11130;
  assign n11132 = ~n11051 & ~n11131;
  assign n11133 = \[1605]  & ~n11132;
  assign n6531 = n11050 | n11133;
  assign n11135 = ~\[1603]  & Ng2691;
  assign n11136 = \[1603]  & ~n11132;
  assign n6536 = n11135 | n11136;
  assign n11138 = ~Ng1315 & Ng2694;
  assign n11139 = Ng1315 & ~n11132;
  assign n6541 = n11138 | n11139;
  assign n11141 = ~\[1605]  & Ng2679;
  assign n11142 = ~n6032 & ~n10933;
  assign n11143 = n11022 & n11101;
  assign n11144 = n11128 & ~n11143;
  assign n11145 = n11053 & n11144;
  assign n11146 = ~n11142 & ~n11145;
  assign n11147 = \[1605]  & ~n11146;
  assign n6546 = n11141 | n11147;
  assign n11149 = ~\[1603]  & Ng2682;
  assign n11150 = \[1603]  & ~n11146;
  assign n6551 = n11149 | n11150;
  assign n11152 = ~Ng1315 & Ng2685;
  assign n11153 = Ng1315 & ~n11146;
  assign n6556 = n11152 | n11153;
  assign n11155 = ~\[1605]  & ~Ng2565;
  assign n11156 = n10921 & n10927;
  assign n11157 = \[1605]  & ~n11156;
  assign n6561 = ~n11155 & ~n11157;
  assign n11159 = ~\[1603]  & ~Ng2568;
  assign n11160 = \[1603]  & ~n11156;
  assign n6566 = ~n11159 & ~n11160;
  assign n11162 = ~Ng1315 & ~Ng2571;
  assign n11163 = Ng1315 & ~n11156;
  assign n6571 = ~n11162 & ~n11163;
  assign n11165 = Ng2580 & Ng2581;
  assign n11166 = \[1603]  & ~n5078;
  assign n11167 = ~\[1603]  & ~Pg16437;
  assign n11168 = ~Ng2580 & ~n11167;
  assign n11169 = ~n11166 & n11168;
  assign n6585 = n11165 | n11169;
  assign n11171 = Pg3229 & Ng2366;
  assign n11172 = ~Pg3229 & ~Ng2380;
  assign n6633 = ~n11171 & ~n11172;
  assign n11174 = Ng1315 & Ng2584;
  assign n11175 = ~Ng1315 & Ng2704;
  assign n6643 = n11174 | n11175;
  assign n11177 = ~Ng1315 & ~Ng2733;
  assign n6648 = ~n6374_1 & ~n11177;
  assign n11179 = \[1603]  & Ng2704;
  assign n11180 = Ng1315 & ~Ng2733;
  assign n11181 = Ng2714 & n11180;
  assign n11182 = ~Ng2714 & ~n11180;
  assign n11183 = ~n11181 & ~n11182;
  assign n6653 = ~n11179 & n11183;
  assign n11185 = Ng2707 & n11181;
  assign n11186 = ~Ng2707 & ~n11181;
  assign n11187 = ~n11179 & ~n11186;
  assign n6658 = ~n11185 & n11187;
  assign n11189 = Ng2727 & n11185;
  assign n11190 = ~Ng2727 & ~n11185;
  assign n11191 = ~n11179 & ~n11190;
  assign n6663 = ~n11189 & n11191;
  assign n11193 = Ng2720 & n11189;
  assign n11194 = ~Ng2720 & ~n11189;
  assign n11195 = ~n11179 & ~n11194;
  assign n6668 = ~n11193 & n11195;
  assign n11197 = Ng2734 & n11193;
  assign n11198 = ~Ng2734 & ~n11193;
  assign n11199 = ~n11179 & ~n11198;
  assign n6673 = ~n11197 & n11199;
  assign n11201 = Ng2746 & n11197;
  assign n11202 = ~Ng2746 & ~n11197;
  assign n11203 = ~n11179 & ~n11202;
  assign n6678 = ~n11201 & n11203;
  assign n11205 = Ng2740 & n11201;
  assign n11206 = ~Ng2740 & ~n11201;
  assign n11207 = ~n11179 & ~n11206;
  assign n6683 = ~n11205 & n11207;
  assign n11209 = Ng2753 & n11205;
  assign n11210 = ~Ng2753 & ~n11205;
  assign n11211 = ~n11179 & ~n11210;
  assign n6688 = ~n11209 & n11211;
  assign n11213 = Ng2760 & n11209;
  assign n11214 = ~Ng2760 & ~n11209;
  assign n11215 = ~n11179 & ~n11214;
  assign n6693 = ~n11213 & n11215;
  assign n11217 = ~Ng2766 & ~n11213;
  assign n11218 = Ng2766 & n11213;
  assign n11219 = ~n11217 & ~n11218;
  assign n6698 = ~n11179 & n11219;
  assign n11221 = Ng2599 & ~Ng2733;
  assign n11222 = Ng2612 & n11221;
  assign n11223 = \[1605]  & n11222;
  assign n11224 = Ng2773 & ~n11223;
  assign n11225 = ~Ng2714 & n11223;
  assign n6703 = n11224 | n11225;
  assign n11227 = \[1603]  & n11222;
  assign n11228 = Ng2774 & ~n11227;
  assign n11229 = ~Ng2714 & n11227;
  assign n6708 = n11228 | n11229;
  assign n11231 = Ng1315 & n11222;
  assign n11232 = Ng2772 & ~n11231;
  assign n11233 = ~Ng2714 & n11231;
  assign n6713 = n11232 | n11233;
  assign n11235 = Ng2776 & ~n11223;
  assign n11236 = ~Ng2707 & n11223;
  assign n6718 = n11235 | n11236;
  assign n11238 = Ng2777 & ~n11227;
  assign n11239 = ~Ng2707 & n11227;
  assign n6723 = n11238 | n11239;
  assign n11241 = Ng2775 & ~n11231;
  assign n11242 = ~Ng2707 & n11231;
  assign n6728 = n11241 | n11242;
  assign n11244 = Ng2779 & ~n11223;
  assign n11245 = ~Ng2727 & n11223;
  assign n6733 = n11244 | n11245;
  assign n11247 = Ng2780 & ~n11227;
  assign n11248 = ~Ng2727 & n11227;
  assign n6738 = n11247 | n11248;
  assign n11250 = Ng2778 & ~n11231;
  assign n11251 = ~Ng2727 & n11231;
  assign n6743 = n11250 | n11251;
  assign n11253 = Ng2782 & ~n11223;
  assign n11254 = ~Ng2720 & n11223;
  assign n6748 = n11253 | n11254;
  assign n11256 = Ng2783 & ~n11227;
  assign n11257 = ~Ng2720 & n11227;
  assign n6753 = n11256 | n11257;
  assign n11259 = Ng2781 & ~n11231;
  assign n11260 = ~Ng2720 & n11231;
  assign n6758 = n11259 | n11260;
  assign n11262 = Ng2785 & ~n11223;
  assign n11263 = ~Ng2734 & n11223;
  assign n6763 = n11262 | n11263;
  assign n11265 = Ng2786 & ~n11227;
  assign n11266 = ~Ng2734 & n11227;
  assign n6768 = n11265 | n11266;
  assign n11268 = Ng2784 & ~n11231;
  assign n11269 = ~Ng2734 & n11231;
  assign n6773 = n11268 | n11269;
  assign n11271 = Ng2788 & ~n11223;
  assign n11272 = ~Ng2746 & n11223;
  assign n6778 = n11271 | n11272;
  assign n11274 = Ng2789 & ~n11227;
  assign n11275 = ~Ng2746 & n11227;
  assign n6783 = n11274 | n11275;
  assign n11277 = Ng2787 & ~n11231;
  assign n11278 = ~Ng2746 & n11231;
  assign n6788 = n11277 | n11278;
  assign n11280 = Ng2791 & ~n11223;
  assign n11281 = ~Ng2740 & n11223;
  assign n6793 = n11280 | n11281;
  assign n11283 = Ng2792 & ~n11227;
  assign n11284 = ~Ng2740 & n11227;
  assign n6798 = n11283 | n11284;
  assign n11286 = Ng2790 & ~n11231;
  assign n11287 = ~Ng2740 & n11231;
  assign n6803 = n11286 | n11287;
  assign n11289 = Ng2794 & ~n11223;
  assign n11290 = ~Ng2753 & n11223;
  assign n6808 = n11289 | n11290;
  assign n11292 = Ng2795 & ~n11227;
  assign n11293 = ~Ng2753 & n11227;
  assign n6813 = n11292 | n11293;
  assign n11295 = Ng2793 & ~n11231;
  assign n11296 = ~Ng2753 & n11231;
  assign n6818 = n11295 | n11296;
  assign n11298 = Ng2797 & ~n11223;
  assign n11299 = ~Ng2760 & n11223;
  assign n6823 = n11298 | n11299;
  assign n11301 = Ng2798 & ~n11227;
  assign n11302 = ~Ng2760 & n11227;
  assign n6828 = n11301 | n11302;
  assign n11304 = Ng2796 & ~n11231;
  assign n11305 = ~Ng2760 & n11231;
  assign n6833 = n11304 | n11305;
  assign n11307 = Ng2800 & ~n11223;
  assign n11308 = ~Ng2766 & n11223;
  assign n6838 = n11307 | n11308;
  assign n11310 = Ng2801 & ~n11227;
  assign n11311 = ~Ng2766 & n11227;
  assign n6843 = n11310 | n11311;
  assign n11313 = Ng2799 & ~n11231;
  assign n11314 = ~Ng2766 & n11231;
  assign n6848 = n11313 | n11314;
  assign n11316 = \[1605]  & Ng2704;
  assign n11317 = ~Ng2803 & ~n11316;
  assign n11318 = ~n10921 & n11316;
  assign n6853 = ~n11317 & ~n11318;
  assign n11320 = ~Ng2804 & ~n11179;
  assign n11321 = ~n10921 & n11179;
  assign n6858 = ~n11320 & ~n11321;
  assign n11323 = Ng1315 & Ng2704;
  assign n11324 = ~Ng2802 & ~n11323;
  assign n11325 = ~n10921 & n11323;
  assign n6863 = ~n11324 & ~n11325;
  assign n11327 = ~Ng2806 & ~n11316;
  assign n11328 = ~n10933 & n11316;
  assign n6868 = ~n11327 & ~n11328;
  assign n11330 = ~Ng2807 & ~n11179;
  assign n11331 = ~n10933 & n11179;
  assign n6873 = ~n11330 & ~n11331;
  assign n11333 = ~Ng2805 & ~n11323;
  assign n11334 = ~n10933 & n11323;
  assign n6878 = ~n11333 & ~n11334;
  assign n11336 = Ng1315 & ~Ng2781;
  assign n11337 = \[1605]  & ~Ng2782;
  assign n11338 = \[1603]  & ~Ng2783;
  assign n11339 = ~n11337 & ~n11338;
  assign n11340 = ~n11336 & n11339;
  assign n11341 = ~Ng2720 & ~n11340;
  assign n11342 = Ng1315 & ~Ng2775;
  assign n11343 = \[1605]  & ~Ng2776;
  assign n11344 = \[1603]  & ~Ng2777;
  assign n11345 = ~n11343 & ~n11344;
  assign n11346 = ~n11342 & n11345;
  assign n11347 = Ng2707 & n11346;
  assign n11348 = ~Ng2707 & ~n11346;
  assign n11349 = ~n11347 & ~n11348;
  assign n11350 = ~n11341 & n11349;
  assign n11351 = Ng1315 & ~Ng2784;
  assign n11352 = \[1605]  & ~Ng2785;
  assign n11353 = \[1603]  & ~Ng2786;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = ~n11351 & n11354;
  assign n11356 = ~Ng2734 & n11355;
  assign n11357 = Ng2734 & ~n11355;
  assign n11358 = ~n11356 & ~n11357;
  assign n11359 = n11350 & ~n11358;
  assign n11360 = Ng1315 & ~Ng2796;
  assign n11361 = \[1605]  & ~Ng2797;
  assign n11362 = \[1603]  & ~Ng2798;
  assign n11363 = ~n11361 & ~n11362;
  assign n11364 = ~n11360 & n11363;
  assign n11365 = Ng2760 & ~n11364;
  assign n11366 = ~Ng2760 & n11364;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = Ng1315 & ~Ng2772;
  assign n11369 = \[1605]  & ~Ng2773;
  assign n11370 = \[1603]  & ~Ng2774;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = ~n11368 & n11371;
  assign n11373 = ~Ng2714 & n11372;
  assign n11374 = Ng2714 & ~n11372;
  assign n11375 = ~n11373 & ~n11374;
  assign n11376 = ~n11367 & ~n11375;
  assign n11377 = Ng1315 & ~Ng2778;
  assign n11378 = \[1605]  & ~Ng2779;
  assign n11379 = \[1603]  & ~Ng2780;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = ~n11377 & n11380;
  assign n11382 = Ng2727 & n11381;
  assign n11383 = Ng1315 & ~Ng2790;
  assign n11384 = \[1605]  & ~Ng2791;
  assign n11385 = \[1603]  & ~Ng2792;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = ~n11383 & n11386;
  assign n11388 = Ng2740 & n11387;
  assign n11389 = ~Ng2740 & ~n11387;
  assign n11390 = ~n11388 & ~n11389;
  assign n11391 = ~n11382 & n11390;
  assign n11392 = n11376 & n11391;
  assign n11393 = n11359 & n11392;
  assign n11394 = ~Ng2727 & ~n11381;
  assign n11395 = Ng1315 & ~Ng2799;
  assign n11396 = \[1605]  & ~Ng2800;
  assign n11397 = \[1603]  & ~Ng2801;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = ~n11395 & n11398;
  assign n11400 = Ng2766 & n11399;
  assign n11401 = ~Ng2766 & ~n11399;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = ~n11394 & n11402;
  assign n11404 = Ng2720 & n11340;
  assign n11405 = Ng1315 & ~Ng2793;
  assign n11406 = \[1605]  & ~Ng2794;
  assign n11407 = \[1603]  & ~Ng2795;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = ~n11405 & n11408;
  assign n11410 = ~Ng2753 & ~n11409;
  assign n11411 = ~n11404 & ~n11410;
  assign n11412 = Ng2753 & n11409;
  assign n11413 = n11411 & ~n11412;
  assign n11414 = Ng1315 & ~Ng2787;
  assign n11415 = \[1605]  & ~Ng2788;
  assign n11416 = \[1603]  & ~Ng2789;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = ~n11414 & n11417;
  assign n11419 = Ng2746 & ~n11418;
  assign n11420 = ~Ng2746 & n11418;
  assign n11421 = ~n11419 & ~n11420;
  assign n11422 = n11413 & ~n11421;
  assign n11423 = n11403 & n11422;
  assign n11424 = n11393 & n11423;
  assign n11425 = Ng1315 & ~Ng2802;
  assign n11426 = Ng1315 & ~Ng2805;
  assign n11427 = \[1605]  & ~Ng2806;
  assign n11428 = \[1603]  & ~Ng2807;
  assign n11429 = ~n11427 & ~n11428;
  assign n11430 = ~n11426 & n11429;
  assign n11431 = \[1605]  & ~Ng2803;
  assign n11432 = \[1603]  & ~Ng2804;
  assign n11433 = ~n11431 & ~n11432;
  assign n11434 = n11430 & n11433;
  assign n11435 = ~n11425 & n11434;
  assign n11436 = ~n11424 & n11435;
  assign n11437 = n11223 & n11436;
  assign n11438 = Ng2809 & ~n11223;
  assign n6883 = n11437 | n11438;
  assign n11440 = n11227 & n11436;
  assign n11441 = Ng2810 & ~n11227;
  assign n6888 = n11440 | n11441;
  assign n11443 = n11231 & n11436;
  assign n11444 = Ng2808 & ~n11231;
  assign n6893 = n11443 | n11444;
  assign n11446 = ~Ng2812 & ~n11223;
  assign n6898 = ~n11316 & ~n11446;
  assign n11448 = ~Ng2813 & ~n11227;
  assign n6903 = ~n11179 & ~n11448;
  assign n11450 = ~Ng2811 & ~n11231;
  assign n6908 = ~n11323 & ~n11450;
  assign n6913 = ~Pg3234 & Ng13475;
  assign n6918 = ~Pg3234 & Ng3054;
  assign n6923 = Pg3234 | Ng3079;
  assign n11455 = ~Ng510 & ~Ng525;
  assign n11456 = ~Ng557 & ~n11455;
  assign n11457 = ~Ng557 & ~Ng525;
  assign n11458 = ~Ng510 & ~n11457;
  assign n11459 = ~n11456 & n11458;
  assign n11460 = ~Ng738 & \[1605] ;
  assign n11461 = ~Ng739 & \[1603] ;
  assign n11462 = ~Ng737 & Ng1315;
  assign n11463 = ~n11461 & ~n11462;
  assign n11464 = ~n11460 & n11463;
  assign n11465 = n6616 & ~n11464;
  assign n11466 = ~n6553 & n11465;
  assign n11467 = ~n6562 & ~n6570;
  assign n11468 = n6538 & n11467;
  assign n11469 = n11466 & n11468;
  assign n11470 = n6579 & ~n6607;
  assign n11471 = n6597 & n11470;
  assign n11472 = ~n6544 & ~n6628_1;
  assign n11473 = n11471 & n11472;
  assign n11474 = n11469 & n11473;
  assign n11475 = n6585_1 & n11474;
  assign n11476 = ~Ng734 & Ng1315;
  assign n11477 = ~Ng736 & \[1603] ;
  assign n11478 = ~Ng735 & \[1605] ;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 = ~n11476 & n11479;
  assign n11481 = ~n11475 & n11480;
  assign n11482 = ~Pg563 & ~Ng559;
  assign n11483 = ~n4984_1 & n11482;
  assign n11484 = ~n1898_1 & n11483;
  assign n11485 = Ng8284 & n11484;
  assign n11486 = ~n11481 & n11485;
  assign n11487 = n11459 & ~n11486;
  assign n11488 = n11458 & n11484;
  assign n11489 = ~Ng529 & n11488;
  assign n11490 = n6131 & ~n6585_1;
  assign n11491 = ~n6131 & n6585_1;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = n11485 & n11492;
  assign n11494 = Ng510 & n11493;
  assign n11495 = n11456 & ~n11494;
  assign n11496 = ~n11489 & n11495;
  assign n6927 = n11487 | n11496;
  assign n11498 = n11459 & ~n11484;
  assign n11499 = Ng8284 & n11459;
  assign n11500 = ~n11481 & n11499;
  assign n11501 = ~n11498 & ~n11500;
  assign n11502 = ~Ng530 & n11488;
  assign n11503 = ~n6116 & ~n6538;
  assign n11504 = n6116 & n6538;
  assign n11505 = ~n11503 & ~n11504;
  assign n11506 = n11485 & ~n11505;
  assign n11507 = Ng510 & n11506;
  assign n11508 = n11456 & ~n11507;
  assign n11509 = ~n11502 & n11508;
  assign n6932 = ~n11501 | n11509;
  assign n11511 = ~Ng531 & n11488;
  assign n11512 = n6131 & n6579;
  assign n11513 = ~n6131 & ~n6579;
  assign n11514 = ~n11512 & ~n11513;
  assign n11515 = n11485 & ~n11514;
  assign n11516 = Ng510 & n11515;
  assign n11517 = n11456 & ~n11516;
  assign n11518 = ~n11511 & n11517;
  assign n6937 = ~n11501 | n11518;
  assign n11520 = ~Ng532 & n11488;
  assign n11521 = ~n6116 & n6597;
  assign n11522 = ~n6116 & ~n11475;
  assign n11523 = ~n6597 & ~n11522;
  assign n11524 = n11485 & ~n11523;
  assign n11525 = ~n11521 & n11524;
  assign n11526 = Ng510 & n11525;
  assign n11527 = n11456 & ~n11526;
  assign n11528 = ~n11520 & n11527;
  assign n6942 = n11487 | n11528;
  assign n11530 = ~Ng533 & n11488;
  assign n11531 = ~n6570 & ~n11475;
  assign n11532 = n6131 & n11531;
  assign n11533 = ~n6131 & ~n11531;
  assign n11534 = ~n11532 & ~n11533;
  assign n11535 = n11485 & n11534;
  assign n11536 = Ng510 & n11535;
  assign n11537 = n11456 & ~n11536;
  assign n11538 = ~n11530 & n11537;
  assign n6947 = n11498 | n11538;
  assign n11540 = ~Ng534 & n11488;
  assign n11541 = ~n6562 & ~n11475;
  assign n11542 = n6116 & n11541;
  assign n11543 = ~n6116 & ~n11541;
  assign n11544 = ~n11542 & ~n11543;
  assign n11545 = n11485 & n11544;
  assign n11546 = Ng510 & n11545;
  assign n11547 = n11456 & ~n11546;
  assign n11548 = ~n11540 & n11547;
  assign n6952 = n11498 | n11548;
  assign n11550 = ~n6544 & ~n11475;
  assign n11551 = ~n6131 & n11550;
  assign n11552 = n6131 & ~n11550;
  assign n11553 = ~n11551 & ~n11552;
  assign n11554 = n11485 & ~n11553;
  assign n11555 = n11459 & ~n11554;
  assign n11556 = ~Ng536 & n11488;
  assign n11557 = ~n6607 & ~n11475;
  assign n11558 = ~n6131 & n11557;
  assign n11559 = n6131 & ~n11557;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = n11485 & ~n11560;
  assign n11562 = Ng510 & n11561;
  assign n11563 = n11456 & ~n11562;
  assign n11564 = ~n11556 & n11563;
  assign n6957 = n11555 | n11564;
  assign n11566 = ~n6553 & ~n11475;
  assign n11567 = ~n6116 & n11566;
  assign n11568 = n6116 & ~n11566;
  assign n11569 = ~n11567 & ~n11568;
  assign n11570 = n11485 & ~n11569;
  assign n11571 = n11459 & ~n11570;
  assign n11572 = ~Ng537 & n11488;
  assign n11573 = ~n6116 & n6616;
  assign n11574 = ~n6616 & ~n11522;
  assign n11575 = n11485 & ~n11574;
  assign n11576 = ~n11573 & n11575;
  assign n11577 = Ng510 & n11576;
  assign n11578 = n11456 & ~n11577;
  assign n11579 = ~n11572 & n11578;
  assign n6962 = n11571 | n11579;
  assign n11581 = n11554 & n11569;
  assign n11582 = n11553 & n11570;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = Ng557 & ~n11583;
  assign n11585 = ~Pg3229 & ~Ng541;
  assign n11586 = Pg3229 & ~Ng538;
  assign n11587 = ~Ng557 & ~n11586;
  assign n11588 = n11488 & n11587;
  assign n11589 = ~n11585 & n11588;
  assign n11590 = ~n11584 & ~n11589;
  assign n11591 = n11493 & n11505;
  assign n11592 = ~n11492 & n11506;
  assign n11593 = ~n11591 & ~n11592;
  assign n11594 = ~n11515 & ~n11593;
  assign n11595 = n11515 & n11593;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = n11576 & n11596;
  assign n11598 = ~n11576 & ~n11596;
  assign n11599 = ~n11597 & ~n11598;
  assign n11600 = ~n11561 & n11599;
  assign n11601 = n11561 & ~n11599;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = n11535 & ~n11544;
  assign n11604 = ~n11534 & n11545;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = ~n11525 & ~n11605;
  assign n11607 = n11525 & n11605;
  assign n11608 = ~n11606 & ~n11607;
  assign n11609 = n11602 & ~n11608;
  assign n11610 = ~n11602 & n11608;
  assign n11611 = ~n11609 & ~n11610;
  assign n11612 = Ng510 & n11611;
  assign n6967 = ~n11590 | n11612;
  assign n11614 = ~Ng1196 & ~Ng1211;
  assign n11615 = ~Ng1243 & ~n11614;
  assign n11616 = ~Ng1243 & ~Ng1211;
  assign n11617 = ~Ng1196 & ~n11616;
  assign n11618 = ~n11615 & n11617;
  assign n11619 = ~n8174 & n8197;
  assign n11620 = n8153 & n11619;
  assign n11621 = \[1605]  & ~Ng1424;
  assign n11622 = \[1603]  & ~Ng1425;
  assign n11623 = Ng1315 & ~Ng1423;
  assign n11624 = ~n11622 & ~n11623;
  assign n11625 = ~n11621 & n11624;
  assign n11626 = n8168 & ~n11625;
  assign n11627 = ~n8217 & n11626;
  assign n11628 = ~n8140 & ~n8207;
  assign n11629 = n8146 & n11628;
  assign n11630 = n11627 & n11629;
  assign n11631 = ~n8162 & ~n8230;
  assign n11632 = n8183 & n11631;
  assign n11633 = n11630 & n11632;
  assign n11634 = n11620 & n11633;
  assign n11635 = Ng1315 & ~Ng1420;
  assign n11636 = \[1603]  & ~Ng1422;
  assign n11637 = \[1605]  & ~Ng1421;
  assign n11638 = ~n11636 & ~n11637;
  assign n11639 = ~n11635 & n11638;
  assign n11640 = ~n11634 & n11639;
  assign n11641 = ~Pg1249 & ~n3404_1;
  assign n11642 = ~Ng1245 & n11641;
  assign n11643 = Ng8293 & n11642;
  assign n11644 = ~n11640 & n11643;
  assign n11645 = n11618 & ~n11644;
  assign n11646 = n11617 & n11642;
  assign n11647 = ~Ng1215 & n11646;
  assign n11648 = ~n7734 & ~n8197;
  assign n11649 = n7734 & n8197;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = n11643 & ~n11650;
  assign n11652 = Ng1196 & n11651;
  assign n11653 = n11615 & ~n11652;
  assign n11654 = ~n11647 & n11653;
  assign n6972 = n11645 | n11654;
  assign n11656 = n11618 & ~n11642;
  assign n11657 = Ng8293 & n11618;
  assign n11658 = ~n11640 & n11657;
  assign n11659 = ~n11656 & ~n11658;
  assign n11660 = ~Ng1216 & n11646;
  assign n11661 = ~n7722 & ~n8146;
  assign n11662 = n7722 & n8146;
  assign n11663 = ~n11661 & ~n11662;
  assign n11664 = n11643 & ~n11663;
  assign n11665 = Ng1196 & n11664;
  assign n11666 = n11615 & ~n11665;
  assign n11667 = ~n11660 & n11666;
  assign n6977 = ~n11659 | n11667;
  assign n11669 = ~Ng1217 & n11646;
  assign n11670 = ~n7734 & n8183;
  assign n11671 = n7734 & ~n8183;
  assign n11672 = ~n11670 & ~n11671;
  assign n11673 = n11643 & n11672;
  assign n11674 = Ng1196 & n11673;
  assign n11675 = n11615 & ~n11674;
  assign n11676 = ~n11669 & n11675;
  assign n6982 = ~n11659 | n11676;
  assign n11678 = ~Ng1218 & n11646;
  assign n11679 = n7722 & n8168;
  assign n11680 = ~n7722 & ~n8168;
  assign n11681 = ~n11679 & ~n11680;
  assign n11682 = n11643 & ~n11681;
  assign n11683 = Ng1196 & n11682;
  assign n11684 = n11615 & ~n11683;
  assign n11685 = ~n11678 & n11684;
  assign n6987 = n11645 | n11685;
  assign n11687 = ~Ng1219 & n11646;
  assign n11688 = ~n8162 & ~n11634;
  assign n11689 = ~n7734 & n11688;
  assign n11690 = n7734 & ~n11688;
  assign n11691 = ~n11689 & ~n11690;
  assign n11692 = n11643 & ~n11691;
  assign n11693 = Ng1196 & n11692;
  assign n11694 = n11615 & ~n11693;
  assign n11695 = ~n11687 & n11694;
  assign n6992 = n11656 | n11695;
  assign n11697 = ~Ng1220 & n11646;
  assign n11698 = ~n8174 & ~n11634;
  assign n11699 = n7722 & n11698;
  assign n11700 = ~n7722 & ~n11698;
  assign n11701 = ~n11699 & ~n11700;
  assign n11702 = n11643 & n11701;
  assign n11703 = Ng1196 & n11702;
  assign n11704 = n11615 & ~n11703;
  assign n11705 = ~n11697 & n11704;
  assign n6997 = n11656 | n11705;
  assign n11707 = ~n8207 & ~n11634;
  assign n11708 = n7734 & n11707;
  assign n11709 = ~n7734 & ~n11707;
  assign n11710 = ~n11708 & ~n11709;
  assign n11711 = n11643 & n11710;
  assign n11712 = n11618 & ~n11711;
  assign n11713 = ~Ng1222 & n11646;
  assign n11714 = ~n8140 & ~n11634;
  assign n11715 = n7734 & n11714;
  assign n11716 = ~n7734 & ~n11714;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = n11643 & n11717;
  assign n11719 = Ng1196 & n11718;
  assign n11720 = n11615 & ~n11719;
  assign n11721 = ~n11713 & n11720;
  assign n7002 = n11712 | n11721;
  assign n11723 = ~n8217 & ~n11634;
  assign n11724 = ~n7722 & n11723;
  assign n11725 = n7722 & ~n11723;
  assign n11726 = ~n11724 & ~n11725;
  assign n11727 = n11643 & ~n11726;
  assign n11728 = n11618 & ~n11727;
  assign n11729 = ~Ng1223 & n11646;
  assign n11730 = ~n7722 & ~n8153;
  assign n11731 = n7722 & n8153;
  assign n11732 = ~n11730 & ~n11731;
  assign n11733 = n11643 & ~n11732;
  assign n11734 = Ng1196 & n11733;
  assign n11735 = n11615 & ~n11734;
  assign n11736 = ~n11729 & n11735;
  assign n7007 = n11728 | n11736;
  assign n11738 = ~Pg3229 & Ng1227;
  assign n11739 = Pg3229 & Ng1224;
  assign n11740 = ~n11738 & ~n11739;
  assign n11741 = n11646 & ~n11740;
  assign n11742 = ~Ng1243 & ~n11741;
  assign n11743 = n11711 & n11726;
  assign n11744 = ~n11710 & n11727;
  assign n11745 = Ng1243 & ~n11744;
  assign n11746 = ~n11743 & n11745;
  assign n11747 = ~n11742 & ~n11746;
  assign n11748 = n11718 & n11732;
  assign n11749 = ~n11717 & n11733;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = n11650 & n11664;
  assign n11752 = n11651 & n11663;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = n11682 & ~n11753;
  assign n11755 = ~n11682 & n11753;
  assign n11756 = ~n11754 & ~n11755;
  assign n11757 = ~n11750 & n11756;
  assign n11758 = n11750 & ~n11756;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = n11692 & ~n11701;
  assign n11761 = n11691 & n11702;
  assign n11762 = ~n11760 & ~n11761;
  assign n11763 = n11673 & n11762;
  assign n11764 = ~n11673 & ~n11762;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = ~n11759 & n11765;
  assign n11767 = n11759 & ~n11765;
  assign n11768 = Ng1196 & ~n11767;
  assign n11769 = ~n11766 & n11768;
  assign n7012 = n11747 | n11769;
  assign n11771 = ~Ng1890 & ~Ng1905;
  assign n11772 = ~Ng1937 & ~n11771;
  assign n11773 = ~Ng1937 & ~Ng1905;
  assign n11774 = ~Ng1890 & ~n11773;
  assign n11775 = ~n11772 & n11774;
  assign n11776 = ~Ng1939 & ~n4911;
  assign n11777 = ~Pg1943 & n11776;
  assign n11778 = \[1603]  & ~Ng2116;
  assign n11779 = ~n9783 & ~n9817;
  assign n11780 = \[1605]  & ~Ng2118;
  assign n11781 = \[1603]  & ~Ng2119;
  assign n11782 = Ng1315 & ~Ng2117;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = ~n11780 & n11783;
  assign n11785 = n9767 & ~n11784;
  assign n11786 = ~n9760 & n11785;
  assign n11787 = n9745 & n9754;
  assign n11788 = ~n9804 & n11787;
  assign n11789 = n11786 & n11788;
  assign n11790 = n9776 & n9793;
  assign n11791 = ~n9739 & n11790;
  assign n11792 = ~n9829 & n11791;
  assign n11793 = n11789 & n11792;
  assign n11794 = n11779 & n11793;
  assign n11795 = \[1605]  & ~Ng2115;
  assign n11796 = Ng1315 & ~Ng2114;
  assign n11797 = ~n11795 & ~n11796;
  assign n11798 = ~n11794 & n11797;
  assign n11799 = ~n11778 & n11798;
  assign n11800 = Ng8302 & ~n11799;
  assign n11801 = n11777 & n11800;
  assign n11802 = n11775 & ~n11801;
  assign n11803 = n11774 & n11777;
  assign n11804 = ~Ng1909 & n11803;
  assign n11805 = Ng8302 & n11777;
  assign n11806 = ~n9332 & n9776;
  assign n11807 = ~n9332 & ~n11794;
  assign n11808 = ~n9776 & ~n11807;
  assign n11809 = ~n11806 & ~n11808;
  assign n11810 = n11805 & n11809;
  assign n11811 = Ng1890 & n11810;
  assign n11812 = n11772 & ~n11811;
  assign n11813 = ~n11804 & n11812;
  assign n7017 = n11802 | n11813;
  assign n11815 = n11777 & ~n11800;
  assign n11816 = n11775 & ~n11815;
  assign n11817 = ~Ng1910 & n11803;
  assign n11818 = ~n9320 & ~n11794;
  assign n11819 = ~n9767 & ~n11818;
  assign n11820 = ~n9320 & n9767;
  assign n11821 = ~n11819 & ~n11820;
  assign n11822 = n11805 & n11821;
  assign n11823 = Ng1890 & n11822;
  assign n11824 = n11772 & ~n11823;
  assign n11825 = ~n11817 & n11824;
  assign n7022 = n11816 | n11825;
  assign n11827 = ~Ng1911 & n11803;
  assign n11828 = ~n9745 & ~n11807;
  assign n11829 = ~n9332 & n9745;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = n11805 & n11830;
  assign n11832 = Ng1890 & n11831;
  assign n11833 = n11772 & ~n11832;
  assign n11834 = ~n11827 & n11833;
  assign n7027 = n11816 | n11834;
  assign n11836 = ~Ng1912 & n11803;
  assign n11837 = ~n9793 & ~n11818;
  assign n11838 = ~n9320 & n9793;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = n11805 & n11839;
  assign n11841 = Ng1890 & n11840;
  assign n11842 = n11772 & ~n11841;
  assign n11843 = ~n11836 & n11842;
  assign n7032 = n11802 | n11843;
  assign n11845 = n11775 & ~n11777;
  assign n11846 = ~Ng1913 & n11803;
  assign n11847 = ~n9760 & ~n11794;
  assign n11848 = n9332 & n11847;
  assign n11849 = ~n9332 & ~n11847;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = n11805 & n11850;
  assign n11852 = Ng1890 & n11851;
  assign n11853 = n11772 & ~n11852;
  assign n11854 = ~n11846 & n11853;
  assign n7037 = n11845 | n11854;
  assign n11856 = ~Ng1914 & n11803;
  assign n11857 = ~n9817 & ~n11794;
  assign n11858 = ~n9320 & ~n11857;
  assign n11859 = n9320 & n11857;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = n11805 & n11860;
  assign n11862 = Ng1890 & n11861;
  assign n11863 = n11772 & ~n11862;
  assign n11864 = ~n11856 & n11863;
  assign n7042 = n11845 | n11864;
  assign n11866 = ~n9739 & ~n11794;
  assign n11867 = n9332 & n11866;
  assign n11868 = ~n9332 & ~n11866;
  assign n11869 = ~n11867 & ~n11868;
  assign n11870 = n11805 & n11869;
  assign n11871 = n11775 & ~n11870;
  assign n11872 = ~Ng1916 & n11803;
  assign n11873 = ~n9783 & ~n11794;
  assign n11874 = ~n9332 & ~n11873;
  assign n11875 = n9332 & n11873;
  assign n11876 = ~n11874 & ~n11875;
  assign n11877 = n11805 & n11876;
  assign n11878 = Ng1890 & n11877;
  assign n11879 = n11772 & ~n11878;
  assign n11880 = ~n11872 & n11879;
  assign n7047 = n11871 | n11880;
  assign n11882 = ~n9804 & ~n11794;
  assign n11883 = n9320 & n11882;
  assign n11884 = ~n9320 & ~n11882;
  assign n11885 = ~n11883 & ~n11884;
  assign n11886 = n11805 & n11885;
  assign n11887 = n11775 & ~n11886;
  assign n11888 = ~Ng1917 & n11803;
  assign n11889 = ~n9754 & ~n11818;
  assign n11890 = ~n9320 & n9754;
  assign n11891 = ~n11889 & ~n11890;
  assign n11892 = n11805 & n11891;
  assign n11893 = Ng1890 & n11892;
  assign n11894 = n11772 & ~n11893;
  assign n11895 = ~n11888 & n11894;
  assign n7052 = n11887 | n11895;
  assign n11897 = ~n11869 & n11886;
  assign n11898 = n11870 & ~n11885;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = Ng1937 & ~n11899;
  assign n11901 = ~Pg3229 & Ng1921;
  assign n11902 = Pg3229 & Ng1918;
  assign n11903 = ~n11901 & ~n11902;
  assign n11904 = n11803 & ~n11903;
  assign n11905 = ~Ng1937 & n11904;
  assign n11906 = ~n11900 & ~n11905;
  assign n11907 = ~n11830 & n11840;
  assign n11908 = n11831 & ~n11839;
  assign n11909 = ~n11907 & ~n11908;
  assign n11910 = n11810 & ~n11821;
  assign n11911 = ~n11809 & n11822;
  assign n11912 = ~n11910 & ~n11911;
  assign n11913 = n11909 & n11912;
  assign n11914 = ~n11909 & ~n11912;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 = n11877 & ~n11891;
  assign n11917 = ~n11876 & n11892;
  assign n11918 = ~n11916 & ~n11917;
  assign n11919 = n11851 & ~n11860;
  assign n11920 = ~n11850 & n11861;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = ~n11918 & n11921;
  assign n11923 = n11918 & ~n11921;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = ~n11915 & n11924;
  assign n11926 = n11915 & ~n11924;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = Ng1890 & n11927;
  assign n7057 = ~n11906 | n11928;
  assign n11930 = ~Ng2584 & ~Ng2599;
  assign n11931 = ~Ng2631 & ~n11930;
  assign n11932 = ~Ng2631 & ~Ng2599;
  assign n11933 = ~Ng2584 & ~n11932;
  assign n11934 = ~n11931 & n11933;
  assign n11935 = ~Pg2637 & ~n6418;
  assign n11936 = ~Ng2633 & n11935;
  assign n11937 = \[1603]  & ~Ng2810;
  assign n11938 = n11372 & ~n11399;
  assign n11939 = ~n11346 & n11938;
  assign n11940 = \[1605]  & ~Ng2812;
  assign n11941 = \[1603]  & ~Ng2813;
  assign n11942 = Ng1315 & ~Ng2811;
  assign n11943 = ~n11941 & ~n11942;
  assign n11944 = ~n11940 & n11943;
  assign n11945 = n11355 & ~n11944;
  assign n11946 = n11409 & n11945;
  assign n11947 = ~n11364 & ~n11381;
  assign n11948 = n11387 & n11947;
  assign n11949 = n11946 & n11948;
  assign n11950 = ~n11340 & ~n11430;
  assign n11951 = n11418 & n11950;
  assign n11952 = n11949 & n11951;
  assign n11953 = n11939 & n11952;
  assign n11954 = \[1605]  & ~Ng2809;
  assign n11955 = Ng1315 & ~Ng2808;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = ~n11953 & n11956;
  assign n11958 = ~n11937 & n11957;
  assign n11959 = Ng8311 & ~n11958;
  assign n11960 = n11936 & n11959;
  assign n11961 = n11934 & ~n11960;
  assign n11962 = n11933 & n11936;
  assign n11963 = ~Ng2603 & n11962;
  assign n11964 = Ng8311 & n11936;
  assign n11965 = n10933 & ~n11409;
  assign n11966 = ~n10933 & n11409;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = n11964 & n11967;
  assign n11969 = Ng2584 & n11968;
  assign n11970 = n11931 & ~n11969;
  assign n11971 = ~n11963 & n11970;
  assign n7062 = n11961 | n11971;
  assign n11973 = n11936 & ~n11959;
  assign n11974 = n11934 & ~n11973;
  assign n11975 = ~Ng2604 & n11962;
  assign n11976 = ~n10921 & ~n11387;
  assign n11977 = n10921 & n11387;
  assign n11978 = ~n11976 & ~n11977;
  assign n11979 = n11964 & ~n11978;
  assign n11980 = Ng2584 & n11979;
  assign n11981 = n11931 & ~n11980;
  assign n11982 = ~n11975 & n11981;
  assign n7067 = n11974 | n11982;
  assign n11984 = ~Ng2605 & n11962;
  assign n11985 = ~n10933 & ~n11418;
  assign n11986 = n10933 & n11418;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = n11964 & ~n11987;
  assign n11989 = Ng2584 & n11988;
  assign n11990 = n11931 & ~n11989;
  assign n11991 = ~n11984 & n11990;
  assign n7072 = n11974 | n11991;
  assign n11993 = ~Ng2606 & n11962;
  assign n11994 = n10921 & ~n11355;
  assign n11995 = ~n10921 & n11355;
  assign n11996 = ~n11994 & ~n11995;
  assign n11997 = n11964 & n11996;
  assign n11998 = Ng2584 & n11997;
  assign n11999 = n11931 & ~n11998;
  assign n12000 = ~n11993 & n11999;
  assign n7077 = n11961 | n12000;
  assign n12002 = n11934 & ~n11936;
  assign n12003 = ~Ng2607 & n11962;
  assign n12004 = ~n11340 & ~n11953;
  assign n12005 = n10933 & n12004;
  assign n12006 = ~n10933 & ~n12004;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = n11964 & n12007;
  assign n12009 = Ng2584 & n12008;
  assign n12010 = n11931 & ~n12009;
  assign n12011 = ~n12003 & n12010;
  assign n7082 = n12002 | n12011;
  assign n12013 = ~Ng2608 & n11962;
  assign n12014 = ~n11381 & ~n11953;
  assign n12015 = n10921 & n12014;
  assign n12016 = ~n10921 & ~n12014;
  assign n12017 = ~n12015 & ~n12016;
  assign n12018 = n11964 & n12017;
  assign n12019 = Ng2584 & n12018;
  assign n12020 = n11931 & ~n12019;
  assign n12021 = ~n12013 & n12020;
  assign n7087 = n12002 | n12021;
  assign n12023 = ~n11399 & ~n11953;
  assign n12024 = n10933 & n12023;
  assign n12025 = ~n10933 & ~n12023;
  assign n12026 = ~n12024 & ~n12025;
  assign n12027 = n11964 & n12026;
  assign n12028 = n11934 & ~n12027;
  assign n12029 = ~Ng2610 & n11962;
  assign n12030 = ~n11346 & ~n11953;
  assign n12031 = n10933 & n12030;
  assign n12032 = ~n10933 & ~n12030;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = n11964 & n12033;
  assign n12035 = Ng2584 & n12034;
  assign n12036 = n11931 & ~n12035;
  assign n12037 = ~n12029 & n12036;
  assign n7092 = n12028 | n12037;
  assign n12039 = ~n11364 & ~n11953;
  assign n12040 = n10921 & n12039;
  assign n12041 = ~n10921 & ~n12039;
  assign n12042 = ~n12040 & ~n12041;
  assign n12043 = n11964 & n12042;
  assign n12044 = n11934 & ~n12043;
  assign n12045 = ~Ng2611 & n11962;
  assign n12046 = n10921 & ~n11372;
  assign n12047 = ~n10921 & n11372;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = n11964 & n12048;
  assign n12050 = Ng2584 & n12049;
  assign n12051 = n11931 & ~n12050;
  assign n12052 = ~n12045 & n12051;
  assign n7097 = n12044 | n12052;
  assign n12054 = n12027 & ~n12042;
  assign n12055 = ~n12026 & n12043;
  assign n12056 = ~n12054 & ~n12055;
  assign n12057 = Ng2631 & ~n12056;
  assign n12058 = ~Pg3229 & Ng2615;
  assign n12059 = Pg3229 & Ng2612;
  assign n12060 = ~n12058 & ~n12059;
  assign n12061 = n11962 & ~n12060;
  assign n12062 = ~Ng2631 & n12061;
  assign n12063 = ~n12057 & ~n12062;
  assign n12064 = ~n12033 & n12049;
  assign n12065 = n12034 & ~n12048;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = n12008 & ~n12017;
  assign n12068 = ~n12007 & n12018;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = ~n12066 & n12069;
  assign n12071 = n12066 & ~n12069;
  assign n12072 = ~n12070 & ~n12071;
  assign n12073 = n11987 & n11997;
  assign n12074 = n11988 & ~n11996;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = n11968 & n11978;
  assign n12077 = ~n11967 & n11979;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = ~n12075 & n12078;
  assign n12080 = n12075 & ~n12078;
  assign n12081 = ~n12079 & ~n12080;
  assign n12082 = ~n12072 & ~n12081;
  assign n12083 = n12072 & n12081;
  assign n12084 = ~n12082 & ~n12083;
  assign n12085 = Ng2584 & n12084;
  assign n7102 = ~n12063 | n12085;
  assign n12087 = Ng13475 & Ng2993;
  assign n12088 = ~Ng13475 & ~Ng2993;
  assign n12089 = ~Pg3234 & ~n12088;
  assign n7107 = ~n12087 & n12089;
  assign n12091 = Ng2998 & n12087;
  assign n12092 = ~Ng2998 & ~n12087;
  assign n12093 = Ng13475 & n6028;
  assign n12094 = ~n12092 & ~n12093;
  assign n12095 = ~n12091 & n12094;
  assign n7112 = Pg3234 | n12095;
  assign n12097 = ~Pg3234 & ~n12093;
  assign n12098 = ~Ng3006 & ~n12091;
  assign n12099 = Ng3006 & n12091;
  assign n12100 = ~n12098 & ~n12099;
  assign n7117 = n12097 & n12100;
  assign n12102 = ~Ng3002 & ~n12099;
  assign n12103 = Ng3002 & n12099;
  assign n12104 = ~n12102 & ~n12103;
  assign n7122 = n12097 & n12104;
  assign n12106 = Ng3013 & n12103;
  assign n12107 = ~Ng3013 & ~n12103;
  assign n12108 = n12097 & ~n12107;
  assign n7127 = ~n12106 & n12108;
  assign n12110 = Ng3010 & n12106;
  assign n12111 = ~Ng3010 & ~n12106;
  assign n12112 = n12097 & ~n12111;
  assign n7132 = ~n12110 & n12112;
  assign n12114 = ~Ng3024 & ~n12110;
  assign n12115 = Ng3024 & n12110;
  assign n12116 = ~n12114 & ~n12115;
  assign n7137 = n12097 & n12116;
  assign n12118 = Ng3018 & n12093;
  assign n12119 = ~Ng3018 & ~n12093;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = ~Ng3028 & ~Ng3036;
  assign n12122 = Ng3032 & n12118;
  assign n12123 = n12121 & n12122;
  assign n12124 = ~Pg3234 & ~n12123;
  assign n7142 = n12120 | ~n12124;
  assign n12126 = ~Ng3028 & ~n12118;
  assign n12127 = Ng3028 & n12118;
  assign n12128 = ~n12126 & ~n12127;
  assign n7147 = n12124 & n12128;
  assign n12130 = Ng3036 & n12127;
  assign n12131 = ~Ng3036 & ~n12127;
  assign n12132 = ~n12130 & ~n12131;
  assign n7152 = n12124 & n12132;
  assign n12134 = ~Ng3032 & ~n12130;
  assign n12135 = Ng3032 & n12130;
  assign n12136 = ~n12134 & ~n12135;
  assign n7157 = n12124 & n12136;
  assign n12138 = Ng3062 & Ng2987;
  assign n12139 = Ng3043 & ~Ng2987;
  assign n7173 = n12138 | n12139;
  assign n12141 = Ng3063 & Ng2987;
  assign n12142 = Ng3044 & ~Ng2987;
  assign n7177 = n12141 | n12142;
  assign n12144 = Ng3064 & Ng2987;
  assign n12145 = Ng3045 & ~Ng2987;
  assign n7181 = n12144 | n12145;
  assign n12147 = Ng3065 & Ng2987;
  assign n12148 = Ng3046 & ~Ng2987;
  assign n7185 = n12147 | n12148;
  assign n12150 = Ng3066 & Ng2987;
  assign n12151 = Ng3047 & ~Ng2987;
  assign n7189 = n12150 | n12151;
  assign n12153 = Ng3067 & Ng2987;
  assign n12154 = Ng3048 & ~Ng2987;
  assign n7193 = n12153 | n12154;
  assign n12156 = Ng3068 & Ng2987;
  assign n12157 = Ng3049 & ~Ng2987;
  assign n7197 = n12156 | n12157;
  assign n12159 = Ng3069 & Ng2987;
  assign n12160 = Ng3050 & ~Ng2987;
  assign n7201 = n12159 | n12160;
  assign n12162 = Ng3070 & Ng2987;
  assign n12163 = Ng3051 & ~Ng2987;
  assign n7205 = n12162 | n12163;
  assign n12165 = ~Pg3231 & Ng3120;
  assign n12166 = ~Pg8270 & Pg8271;
  assign n12167 = Pg8270 & ~Pg8271;
  assign n12168 = ~n12166 & ~n12167;
  assign n12169 = Pg8275 & Pg8274;
  assign n12170 = ~Pg8275 & ~Pg8274;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = n12168 & n12171;
  assign n12173 = ~n12168 & ~n12171;
  assign n12174 = ~n12172 & ~n12173;
  assign n12175 = ~Pg8268 & Pg8269;
  assign n12176 = Pg8268 & ~Pg8269;
  assign n12177 = ~n12175 & ~n12176;
  assign n12178 = Pg8273 & Pg8272;
  assign n12179 = ~Pg8273 & ~Pg8272;
  assign n12180 = ~n12178 & ~n12179;
  assign n12181 = ~n12177 & n12180;
  assign n12182 = n12177 & ~n12180;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = n12174 & n12183;
  assign n12185 = ~n12174 & ~n12183;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~n12165 & ~n12186;
  assign n12188 = n12165 & n12186;
  assign n7210 = n12187 | n12188;
  assign n12190 = Ng3083 & ~n12186;
  assign n12191 = ~Ng3083 & n12186;
  assign n7214 = ~n12190 & ~n12191;
  assign n12193 = Ng3071 & Ng2987;
  assign n12194 = Ng3052 & ~Ng2987;
  assign n7219 = n12193 | n12194;
  assign n12196 = Ng3072 & Ng2987;
  assign n12197 = Ng3053 & ~Ng2987;
  assign n7223 = n12196 | n12197;
  assign n12199 = Ng3073 & Ng2987;
  assign n12200 = Ng3055 & ~Ng2987;
  assign n7227 = n12199 | n12200;
  assign n12202 = Ng3074 & Ng2987;
  assign n12203 = Ng3056 & ~Ng2987;
  assign n7231 = n12202 | n12203;
  assign n12205 = Ng3075 & Ng2987;
  assign n12206 = Ng3057 & ~Ng2987;
  assign n7235 = n12205 | n12206;
  assign n12208 = Ng3076 & Ng2987;
  assign n12209 = Ng3058 & ~Ng2987;
  assign n7239 = n12208 | n12209;
  assign n12211 = Ng3077 & Ng2987;
  assign n12212 = Ng3059 & ~Ng2987;
  assign n7243 = n12211 | n12212;
  assign n12214 = Ng3078 & Ng2987;
  assign n12215 = Ng3060 & ~Ng2987;
  assign n7247 = n12214 | n12215;
  assign n12217 = Ng2997 & Ng2987;
  assign n12218 = Ng3061 & ~Ng2987;
  assign n7251 = n12217 | n12218;
  assign n12220 = ~Pg8261 & Pg8259;
  assign n12221 = Pg8261 & ~Pg8259;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = Pg8266 & Pg8265;
  assign n12224 = ~Pg8266 & ~Pg8265;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = n12222 & n12225;
  assign n12227 = ~n12222 & ~n12225;
  assign n12228 = ~n12226 & ~n12227;
  assign n12229 = ~Pg8263 & Pg8260;
  assign n12230 = Pg8263 & ~Pg8260;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = Pg8264 & Pg8262;
  assign n12233 = ~Pg8264 & ~Pg8262;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = ~n12231 & n12234;
  assign n12236 = n12231 & ~n12234;
  assign n12237 = ~n12235 & ~n12236;
  assign n12238 = n12228 & n12237;
  assign n12239 = ~n12228 & ~n12237;
  assign n12240 = ~n12238 & ~n12239;
  assign n12241 = Ng2990 & ~n12240;
  assign n12242 = ~Ng2990 & n12240;
  assign n7256 = ~n12241 & ~n12242;
  assign n12244 = ~n12165 & ~n12240;
  assign n12245 = n12165 & n12240;
  assign n7261 = n12244 | n12245;
  assign Pg27380 = ~n894_1;
  assign Pg26135 = ~n854_1;
  assign Pg25435 = ~n864_1;
  assign Pg24734 = ~n869_1;
  assign n1534 = ~Ng125;
  assign n1543 = ~Ng121;
  assign n1552_1 = ~Ng117;
  assign n1561_1 = ~Ng113;
  assign n1570_1 = ~Ng109;
  assign n1579_1 = ~Ng105;
  assign n1588 = ~Ng101;
  assign n1597_1 = ~Ng97;
  assign n2073 = ~Ng451;
  assign n2078_1 = ~Ng453;
  assign n2083_1 = ~Ng279;
  assign n2088_1 = ~Ng281;
  assign n2093_1 = ~Ng283;
  assign n2098 = ~Ng285;
  assign n2103 = ~Ng287;
  assign n2108_1 = ~Ng289;
  assign n2118 = ~Ng291;
  assign n3040 = ~Ng813;
  assign n3049_1 = ~Ng809;
  assign n3058_1 = ~Ng805;
  assign n3067_1 = ~Ng801;
  assign n3076_1 = ~Ng797;
  assign n3085_1 = ~Ng793;
  assign n3094_1 = ~Ng789;
  assign n3103_1 = ~Ng785;
  assign n3579_1 = ~Ng1138;
  assign n3584_1 = ~Ng1140;
  assign n3589_1 = ~Ng966;
  assign n3594_1 = ~Ng968;
  assign n3599_1 = ~Ng970;
  assign n3604_1 = ~Ng972;
  assign n3609_1 = ~Ng974;
  assign n3614_1 = ~Ng976;
  assign n3624_1 = ~Ng978;
  assign n4547 = ~Ng1506;
  assign n4556 = ~Ng1501;
  assign n4565 = ~Ng1496;
  assign n4574 = ~Ng1491;
  assign n4583 = ~Ng1486;
  assign n4592 = ~Ng1481;
  assign n4601 = ~Ng1476;
  assign n4610 = ~Ng1471;
  assign n5086 = ~Ng1832;
  assign n5091 = ~Ng1834;
  assign n5096 = ~Ng1660;
  assign n5101 = ~Ng1662;
  assign n5106 = ~Ng1664;
  assign n5111 = ~Ng1666;
  assign n5116 = ~Ng1668;
  assign n5121 = ~Ng1670;
  assign n5131 = ~Ng1672;
  assign n6054 = ~Ng2200;
  assign n6063 = ~Ng2195;
  assign n6072 = ~Ng2190;
  assign n6081 = ~Ng2185;
  assign n6090 = ~Ng2180;
  assign n6099 = ~Ng2175;
  assign n6108 = ~Ng2170;
  assign n6117 = ~Ng2165;
  assign n6593 = ~Ng2526;
  assign n6598 = ~Ng2528;
  assign n6603 = ~Ng2354;
  assign n6608 = ~Ng2356;
  assign n6613 = ~Ng2358;
  assign n6618 = ~Ng2360;
  assign n6623 = ~Ng2362;
  assign n6628 = ~Ng2364;
  assign n6638 = ~Ng2366;
  assign Pg25420 = Pg25442;
  assign Pg8167 = \[1594] ;
  assign Pg8106 = \[1605] ;
  assign Pg8087 = \[1612] ;
  assign Pg8082 = \[1594] ;
  assign Pg8030 = \[1603] ;
  assign Pg8012 = \[1612] ;
  assign Pg8007 = \[1594] ;
  assign Pg7961 = \[1612] ;
  assign Pg7956 = \[1594] ;
  assign Pg7909 = \[1612] ;
  assign Pg7487 = \[1603] ;
  assign Pg7425 = \[1605] ;
  assign Pg7390 = \[1603] ;
  assign Pg7357 = \[1603] ;
  assign Pg7302 = \[1605] ;
  assign Pg7264 = \[1594] ;
  assign Pg7229 = \[1605] ;
  assign Pg7194 = \[1603] ;
  assign Pg7161 = \[1603] ;
  assign Pg7084 = \[1594] ;
  assign Pg7052 = \[1605] ;
  assign Pg7014 = \[1594] ;
  assign Pg6979 = \[1605] ;
  assign Pg6944 = \[1603] ;
  assign Pg6911 = \[1603] ;
  assign Pg6837 = \[1612] ;
  assign Pg6782 = \[1594] ;
  assign Pg6750 = \[1605] ;
  assign Pg6712 = \[1594] ;
  assign Pg6677 = \[1605] ;
  assign Pg6642 = \[1603] ;
  assign Pg6573 = \[1612] ;
  assign Pg6518 = \[1594] ;
  assign Pg6485 = \[1605] ;
  assign Pg6447 = \[1594] ;
  assign Pg6368 = \[1612] ;
  assign Pg6313 = \[1594] ;
  assign Pg6231 = \[1612] ;
  assign Pg5796 = \[1603] ;
  assign Pg5747 = \[1605] ;
  assign Pg5738 = \[1603] ;
  assign Pg5695 = \[1605] ;
  assign Pg5686 = \[1603] ;
  assign Pg5657 = \[1605] ;
  assign Pg5648 = \[1603] ;
  assign Pg5637 = \[1609] ;
  assign Pg5629 = \[1605] ;
  assign Pg5612 = \[1609] ;
  assign Pg5595 = \[1609] ;
  assign Pg5555 = \[1612] ;
  assign Pg5549 = \[1609] ;
  assign Pg5511 = \[1612] ;
  assign Pg5472 = \[1612] ;
  assign Pg5437 = \[1612] ;
  assign n271_1 = Pg51;
  assign n354_1 = Pg8021;
  assign n363_1 = Pg3212;
  assign n367_1 = Pg3228;
  assign n371_1 = Pg3227;
  assign n375_1 = Pg3226;
  assign n379_1 = Pg3225;
  assign n383_1 = Pg3224;
  assign n387_1 = Pg3223;
  assign n391_1 = Pg3222;
  assign n395_1 = Pg3221;
  assign n399_1 = Pg3232;
  assign n403_1 = Pg3220;
  assign n407_1 = Pg3219;
  assign n411_1 = Pg3218;
  assign n415 = Pg3217;
  assign n419_1 = Pg3216;
  assign n423_1 = Pg3215;
  assign n427 = Pg3214;
  assign n431_1 = Pg3213;
  assign n484 = Pg8251;
  assign n492_1 = Pg4090;
  assign n500 = Pg4323;
  assign n508_1 = Pg4590;
  assign n516_1 = Pg6225;
  assign n524_1 = Pg6442;
  assign n532_1 = Pg6895;
  assign n540_1 = Pg7334;
  assign n548_1 = Pg7519;
  assign n556_1 = Pg8249;
  assign n564_1 = Pg4088;
  assign n572_1 = Pg4321;
  assign n580_1 = Pg8023;
  assign n588 = Pg8175;
  assign n596_1 = Pg3993;
  assign n604_1 = Pg4200;
  assign n612_1 = Pg4450;
  assign n620_1 = Pg8096;
  assign n849_1 = Pg24734;
  assign n859_1 = Pg25442;
  assign n873_1 = Pg26104;
  assign n877_1 = Pg25435;
  assign n881_1 = Pg27380;
  assign n885_1 = Pg26149;
  assign n889_1 = Pg26135;
  assign n1538_1 = Ng450;
  assign n1547_1 = Ng452;
  assign n1556_1 = Ng454;
  assign n1565_1 = Ng280;
  assign n1574 = Ng282;
  assign n1583 = Ng284;
  assign n1592 = Ng286;
  assign n1601 = Ng288;
  assign n1605_1 = Ng13407;
  assign n1609_1 = Ng290;
  assign n1628_1 = Ng11497;
  assign n1632 = Ng342;
  assign n1636_1 = Ng11498;
  assign n1640_1 = Ng350;
  assign n1644_1 = Ng11499;
  assign n1648_1 = Ng352;
  assign n1652_1 = Ng11500;
  assign n1656_1 = Ng357;
  assign n1660 = Ng11501;
  assign n1664_1 = Ng365;
  assign n1668 = Ng11502;
  assign n1672 = Ng367;
  assign n1676_1 = Ng11503;
  assign n1680 = Ng372;
  assign n1684 = Ng11504;
  assign n1688_1 = Ng380;
  assign n1692_1 = Ng11505;
  assign n1696_1 = Ng382;
  assign n1700_1 = Ng11506;
  assign n1704_1 = Ng387;
  assign n1708 = Ng11507;
  assign n1712 = Ng395;
  assign n1716_1 = Ng11508;
  assign n1720_1 = Ng397;
  assign n1744_1 = Ng513;
  assign n1748 = Ng523;
  assign n1753_1 = Ng11512;
  assign n1757_1 = Ng564;
  assign n1762_1 = Ng11515;
  assign n1766_1 = Ng570;
  assign n1771_1 = Ng11516;
  assign n1775_1 = Ng572;
  assign n1780_1 = Ng11517;
  assign n1784_1 = Ng574;
  assign n1789_1 = Ng11513;
  assign n1793 = Ng566;
  assign n1798 = Ng11514;
  assign n1802_1 = Ng568;
  assign n1880_1 = Ng528;
  assign n1884_1 = Ng535;
  assign n1893_1 = Ng543;
  assign n1907_1 = Ng549;
  assign n1916_1 = Ng558;
  assign n2055_1 = Ng8284;
  assign n2068_1 = Pg16297;
  assign n2392 = Ng13457;
  assign n2396_1 = \[1612] ;
  assign n2400_1 = \[1594] ;
  assign n3044_1 = Ng1137;
  assign n3053_1 = Ng1139;
  assign n3062_1 = Ng1141;
  assign n3071_1 = Ng967;
  assign n3080_1 = Ng969;
  assign n3089_1 = Ng971;
  assign n3098_1 = Ng973;
  assign n3107 = Ng975;
  assign n3111_1 = Ng13423;
  assign n3115_1 = Ng977;
  assign n3134 = Ng11524;
  assign n3138_1 = Ng1029;
  assign n3142_1 = Ng11525;
  assign n3146_1 = Ng1037;
  assign n3150 = Ng11526;
  assign n3154_1 = Ng1039;
  assign n3158_1 = Ng11527;
  assign n3162_1 = Ng1044;
  assign n3166 = Ng11528;
  assign n3170_1 = Ng1052;
  assign n3174_1 = Ng11529;
  assign n3178_1 = Ng1054;
  assign n3182_1 = Ng11530;
  assign n3186_1 = Ng1059;
  assign n3190_1 = Ng11531;
  assign n3194_1 = Ng1067;
  assign n3198_1 = Ng11532;
  assign n3202_1 = Ng1069;
  assign n3206_1 = Ng11533;
  assign n3210_1 = Ng1074;
  assign n3214_1 = Ng11534;
  assign n3218_1 = Ng1082;
  assign n3222_1 = Ng11535;
  assign n3226_1 = Ng1084;
  assign n3250_1 = Ng1199;
  assign n3254_1 = Ng1209;
  assign n3259_1 = Ng11539;
  assign n3263_1 = Ng1250;
  assign n3268_1 = Ng11542;
  assign n3272_1 = Ng1256;
  assign n3277_1 = Ng11543;
  assign n3281_1 = Ng1258;
  assign n3286_1 = Ng11544;
  assign n3290_1 = Ng1260;
  assign n3295_1 = Ng11540;
  assign n3299_1 = Ng1252;
  assign n3304_1 = Ng11541;
  assign n3308_1 = Ng1254;
  assign n3386_1 = Ng1214;
  assign n3390_1 = Ng1221;
  assign n3399_1 = Ng1229;
  assign n3413_1 = Ng1235;
  assign n3422_1 = Ng1244;
  assign n3561_1 = Ng8293;
  assign n3574_1 = Pg16355;
  assign n3629_1 = Ng13475;
  assign n3633_1 = \[1605] ;
  assign n3637_1 = \[1603] ;
  assign n4551 = Ng1831;
  assign n4560 = Ng1833;
  assign n4569 = Ng1835;
  assign n4578 = Ng1661;
  assign n4587 = Ng1663;
  assign n4596 = Ng1665;
  assign n4605 = Ng1667;
  assign n4614 = Ng1669;
  assign n4618 = Ng13439;
  assign n4622 = Ng1671;
  assign n4641 = Ng11551;
  assign n4645 = Ng1723;
  assign n4649 = Ng11552;
  assign n4653 = Ng1731;
  assign n4657 = Ng11553;
  assign n4661 = Ng1733;
  assign n4665 = Ng11554;
  assign n4669 = Ng1738;
  assign n4673 = Ng11555;
  assign n4677 = Ng1746;
  assign n4681 = Ng11556;
  assign n4685 = Ng1748;
  assign n4689 = Ng11557;
  assign n4693 = Ng1753;
  assign n4697 = Ng11558;
  assign n4701 = Ng1761;
  assign n4705 = Ng11559;
  assign n4709 = Ng1763;
  assign n4713 = Ng11560;
  assign n4717 = Ng1768;
  assign n4721 = Ng11561;
  assign n4725 = Ng1776;
  assign n4729 = Ng11562;
  assign n4733 = Ng1778;
  assign n4757 = Ng1893;
  assign n4761 = Ng1903;
  assign n4766 = Ng11566;
  assign n4770 = Ng1944;
  assign n4775 = Ng11569;
  assign n4779 = Ng1950;
  assign n4784 = Ng11570;
  assign n4788 = Ng1952;
  assign n4793 = Ng11571;
  assign n4797 = Ng1954;
  assign n4802 = Ng11567;
  assign n4806 = Ng1946;
  assign n4811 = Ng11568;
  assign n4815 = Ng1948;
  assign n4893_1 = Ng1908;
  assign n4897_1 = Ng1915;
  assign n4906_1 = Ng1923;
  assign n4920 = Ng1929;
  assign n4929 = Ng1938;
  assign n5068 = Ng8302;
  assign n5081 = Pg16399;
  assign n5820 = Ng2256;
  assign n5824 = \[1609] ;
  assign n6058 = Ng2525;
  assign n6067 = Ng2527;
  assign n6076 = Ng2529;
  assign n6085 = Ng2355;
  assign n6094 = Ng2357;
  assign n6103 = Ng2359;
  assign n6112 = Ng2361;
  assign n6121 = Ng2363;
  assign n6125 = Ng13455;
  assign n6129 = Ng2365;
  assign n6148 = Ng11578;
  assign n6152 = Ng2417;
  assign n6156 = Ng11579;
  assign n6160 = Ng2425;
  assign n6164 = Ng11580;
  assign n6168 = Ng2427;
  assign n6172 = Ng11581;
  assign n6176 = Ng2432;
  assign n6180 = Ng11582;
  assign n6184 = Ng2440;
  assign n6188 = Ng11583;
  assign n6192 = Ng2442;
  assign n6196 = Ng11584;
  assign n6200 = Ng2447;
  assign n6204 = Ng11585;
  assign n6208 = Ng2455;
  assign n6212 = Ng11586;
  assign n6216 = Ng2457;
  assign n6220 = Ng11587;
  assign n6224 = Ng2462;
  assign n6228 = Ng11588;
  assign n6232 = Ng2470;
  assign n6236 = Ng11589;
  assign n6240 = Ng2472;
  assign n6264 = Ng2587;
  assign n6268 = Ng2597;
  assign n6273 = Ng11593;
  assign n6277 = Ng2638;
  assign n6282 = Ng11596;
  assign n6286 = Ng2644;
  assign n6291 = Ng11597;
  assign n6295 = Ng2646;
  assign n6300 = Ng11598;
  assign n6304 = Ng2648;
  assign n6309 = Ng11594;
  assign n6313 = Ng2640;
  assign n6318 = Ng11595;
  assign n6322 = Ng2642;
  assign n6400 = Ng2602;
  assign n6404 = Ng2609;
  assign n6413 = Ng2617;
  assign n6427 = Ng2623;
  assign n6436 = Ng2632;
  assign n6575 = Ng8311;
  assign n6588 = Pg16437;
  assign n7161 = Pg3234;
  assign n7164 = Pg5388;
  assign n7168 = Pg16496;
  always @ (posedge clock) begin
    Pg8021 <= n271_1;
    Ng2817 <= n275_1;
    Ng2933 <= n280;
    Ng13457 <= n285_1;
    Ng2883 <= n290_1;
    Ng2888 <= n295_1;
    Ng2896 <= n300_1;
    Ng2892 <= n305_1;
    Ng2903 <= n310_1;
    Ng2900 <= n315;
    Ng2908 <= n320_1;
    Ng2912 <= n325_1;
    Ng2917 <= n330_1;
    Ng2924 <= n335_1;
    Ng2920 <= n340_1;
    Ng2984 <= n345_1;
    Ng2985 <= n350_1;
    Ng2929 <= n354_1;
    Ng2879 <= n359_1;
    Ng2934 <= n363_1;
    Ng2935 <= n367_1;
    Ng2938 <= n371_1;
    Ng2941 <= n375_1;
    Ng2944 <= n379_1;
    Ng2947 <= n383_1;
    Ng2953 <= n387_1;
    Ng2956 <= n391_1;
    Ng2959 <= n395_1;
    Ng2962 <= n399_1;
    Ng2963 <= n403_1;
    Ng2966 <= n407_1;
    Ng2969 <= n411_1;
    Ng2972 <= n415;
    Ng2975 <= n419_1;
    Ng2978 <= n423_1;
    Ng2981 <= n427;
    Ng2874 <= n431_1;
    Ng1506 <= n436;
    Ng1501 <= n441_1;
    Ng1496 <= n446_1;
    Ng1491 <= n451;
    Ng1486 <= n456;
    Ng1481 <= n461_1;
    Ng1476 <= n466_1;
    Ng1471 <= n471_1;
    Ng13439 <= n476_1;
    Pg8251 <= n481;
    Ng813 <= n484;
    Pg4090 <= n489;
    Ng809 <= n492_1;
    Pg4323 <= n497_1;
    Ng805 <= n500;
    Pg4590 <= n505_1;
    Ng801 <= n508_1;
    Pg6225 <= n513_1;
    Ng797 <= n516_1;
    Pg6442 <= n521_1;
    Ng793 <= n524_1;
    Pg6895 <= n529_1;
    Ng789 <= n532_1;
    Pg7334 <= n537_1;
    Ng785 <= n540_1;
    Pg7519 <= n545_1;
    Ng13423 <= n548_1;
    Pg8249 <= n553_1;
    Ng125 <= n556_1;
    Pg4088 <= n561_1;
    Ng121 <= n564_1;
    Pg4321 <= n569_1;
    Ng117 <= n572_1;
    Pg8023 <= n577_1;
    Ng113 <= n580_1;
    Pg8175 <= n585_1;
    Ng109 <= n588;
    Pg3993 <= n593;
    Ng105 <= n596_1;
    Pg4200 <= n601_1;
    Ng101 <= n604_1;
    Pg4450 <= n609_1;
    Ng97 <= n612_1;
    Pg8096 <= n617_1;
    Ng13407 <= n620_1;
    Ng2200 <= n625_1;
    Ng2195 <= n630;
    Ng2190 <= n635_1;
    Ng2185 <= n640_1;
    Ng2180 <= n645_1;
    Ng2175 <= n650;
    Ng2170 <= n655;
    Ng2165 <= n660;
    Ng13455 <= n665_1;
    Ng3210 <= n670;
    Ng3211 <= n675_1;
    Ng3084 <= n680;
    Ng3085 <= n685_1;
    Ng3086 <= n690;
    Ng3087 <= n695_1;
    Ng3091 <= n700_1;
    Ng3092 <= n705_1;
    Ng3093 <= n710_1;
    Ng3094 <= n715_1;
    Ng3095 <= n720;
    Ng3096 <= n725;
    Ng3097 <= n730_1;
    Ng3098 <= n735_1;
    Ng3099 <= n740_1;
    Ng3100 <= n745_1;
    Ng3101 <= n750_1;
    Ng3102 <= n755_1;
    Ng3103 <= n760_1;
    Ng3104 <= n765_1;
    Ng3105 <= n770_1;
    Ng3106 <= n775_1;
    Ng3107 <= n780_1;
    Ng3108 <= n785_1;
    Ng3155 <= n790_1;
    Ng3158 <= n795_1;
    Ng3161 <= n800_1;
    Ng3164 <= n805_1;
    Ng3167 <= n810_1;
    Ng3170 <= n815_1;
    Ng3173 <= n820;
    Ng3176 <= n825_1;
    Ng3179 <= n830_1;
    Ng3182 <= n835_1;
    Ng3185 <= n840_1;
    Ng3088 <= n845_1;
    Ng3191 <= n849_1;
    Ng3128 <= n854_1;
    Ng3126 <= n859_1;
    Ng3125 <= n864_1;
    Ng3123 <= n869_1;
    Ng3120 <= n873_1;
    Ng3110 <= n877_1;
    Ng3139 <= n881_1;
    Ng3135 <= n885_1;
    Ng3147 <= n889_1;
    Ng185 <= n894_1;
    Ng130 <= n899_1;
    Ng131 <= n904_1;
    Ng129 <= n909_1;
    Ng133 <= n914_1;
    Ng134 <= n919_1;
    Ng132 <= n924_1;
    Ng142 <= n929_1;
    Ng143 <= n934;
    Ng141 <= n939_1;
    Ng145 <= n944_1;
    Ng146 <= n949_1;
    Ng144 <= n954_1;
    Ng148 <= n959_1;
    Ng149 <= n964_1;
    Ng147 <= n969_1;
    Ng151 <= n974_1;
    Ng152 <= n979_1;
    Ng150 <= n984_1;
    Ng154 <= n989_1;
    Ng155 <= n994_1;
    Ng153 <= n999_1;
    Ng157 <= n1004_1;
    Ng158 <= n1009_1;
    Ng156 <= n1014;
    Ng160 <= n1019_1;
    Ng161 <= n1024_1;
    Ng159 <= n1029;
    Ng163 <= n1034_1;
    Ng164 <= n1039_1;
    Ng162 <= n1044;
    Ng169 <= n1049;
    Ng170 <= n1054_1;
    Ng168 <= n1059_1;
    Ng172 <= n1064_1;
    Ng173 <= n1069;
    Ng171 <= n1074_1;
    Ng175 <= n1079;
    Ng176 <= n1084_1;
    Ng174 <= n1089_1;
    Ng178 <= n1094_1;
    Ng179 <= n1099_1;
    Ng177 <= n1104_1;
    Ng186 <= n1109_1;
    Ng189 <= n1114;
    Ng192 <= n1119_1;
    Ng231 <= n1124_1;
    Ng234 <= n1129_1;
    Ng237 <= n1134_1;
    Ng195 <= n1139_1;
    Ng198 <= n1144_1;
    Ng201 <= n1149_1;
    Ng240 <= n1154_1;
    Ng243 <= n1159_1;
    Ng246 <= n1164;
    Ng204 <= n1169_1;
    Ng207 <= n1174_1;
    Ng210 <= n1179_1;
    Ng249 <= n1184_1;
    Ng252 <= n1189_1;
    Ng255 <= n1194;
    Ng213 <= n1199_1;
    Ng216 <= n1204_1;
    Ng219 <= n1209_1;
    Ng258 <= n1214_1;
    Ng261 <= n1219_1;
    Ng264 <= n1224_1;
    Ng222 <= n1229_1;
    Ng225 <= n1234_1;
    Ng228 <= n1239_1;
    Ng267 <= n1244_1;
    Ng270 <= n1249_1;
    Ng273 <= n1254_1;
    Ng92 <= n1259_1;
    Ng88 <= n1264_1;
    Ng83 <= n1269;
    Ng79 <= n1274;
    Ng74 <= n1279;
    Ng70 <= n1284_1;
    Ng65 <= n1289;
    Ng61 <= n1294;
    Ng56 <= n1299;
    Ng52 <= n1304;
    Ng11497 <= n1309;
    Ng11498 <= n1314_1;
    Ng11499 <= n1319;
    Ng11500 <= n1324_1;
    Ng11501 <= n1329_1;
    Ng11502 <= n1334_1;
    Ng11503 <= n1339_1;
    Ng11504 <= n1344_1;
    Ng11505 <= n1349_1;
    Ng11506 <= n1354;
    Ng11507 <= n1359;
    Ng11508 <= n1364;
    Ng408 <= n1369;
    Ng411 <= n1374_1;
    Ng414 <= n1379;
    Ng417 <= n1384_1;
    Ng420 <= n1389_1;
    Ng423 <= n1394_1;
    Ng427 <= n1399_1;
    Ng428 <= n1404_1;
    Ng426 <= n1409_1;
    Ng429 <= n1414;
    Ng432 <= n1419;
    Ng435 <= n1424_1;
    Ng438 <= n1429_1;
    Ng441 <= n1434;
    Ng444 <= n1439_1;
    Ng448 <= n1444_1;
    Ng449 <= n1449;
    Ng447 <= n1454;
    Ng312 <= n1459_1;
    Ng313 <= n1464;
    Ng314 <= n1469_1;
    Ng315 <= n1474_1;
    Ng316 <= n1479_1;
    Ng317 <= n1484_1;
    Ng318 <= n1489;
    Ng319 <= n1494_1;
    Ng320 <= n1499;
    Ng322 <= n1504;
    Ng323 <= n1509_1;
    Ng321 <= n1514_1;
    Ng403 <= n1519_1;
    Ng404 <= n1524_1;
    Ng402 <= n1529_1;
    Ng450 <= n1534;
    Ng451 <= n1538_1;
    Ng452 <= n1543;
    Ng453 <= n1547_1;
    Ng454 <= n1552_1;
    Ng279 <= n1556_1;
    Ng280 <= n1561_1;
    Ng281 <= n1565_1;
    Ng282 <= n1570_1;
    Ng283 <= n1574;
    Ng284 <= n1579_1;
    Ng285 <= n1583;
    Ng286 <= n1588;
    Ng287 <= n1592;
    Ng288 <= n1597_1;
    Ng289 <= n1601;
    Ng290 <= n1605_1;
    Ng291 <= n1609_1;
    Ng299 <= n1614_1;
    Ng305 <= n1619_1;
    Ng298 <= n1624_1;
    Ng342 <= n1628_1;
    Ng349 <= n1632;
    Ng350 <= n1636_1;
    Ng351 <= n1640_1;
    Ng352 <= n1644_1;
    Ng353 <= n1648_1;
    Ng357 <= n1652_1;
    Ng364 <= n1656_1;
    Ng365 <= n1660;
    Ng366 <= n1664_1;
    Ng367 <= n1668;
    Ng368 <= n1672;
    Ng372 <= n1676_1;
    Ng379 <= n1680;
    Ng380 <= n1684;
    Ng381 <= n1688_1;
    Ng382 <= n1692_1;
    Ng383 <= n1696_1;
    Ng387 <= n1700_1;
    Ng394 <= n1704_1;
    Ng395 <= n1708;
    Ng396 <= n1712;
    Ng397 <= n1716_1;
    Ng324 <= n1720_1;
    Ng554 <= n1725;
    Ng557 <= n1730;
    Ng510 <= n1735_1;
    Ng513 <= n1740;
    Ng523 <= n1744_1;
    Ng524 <= n1748;
    Ng564 <= n1753_1;
    Ng569 <= n1757_1;
    Ng570 <= n1762_1;
    Ng571 <= n1766_1;
    Ng572 <= n1771_1;
    Ng573 <= n1775_1;
    Ng574 <= n1780_1;
    Ng565 <= n1784_1;
    Ng566 <= n1789_1;
    Ng567 <= n1793;
    Ng568 <= n1798;
    Ng489 <= n1802_1;
    Ng486 <= n1807_1;
    Ng487 <= n1812_1;
    Ng488 <= n1817_1;
    Ng11512 <= n1822_1;
    Ng11515 <= n1826_1;
    Ng11516 <= n1830_1;
    Ng477 <= n1834_1;
    Ng478 <= n1839;
    Ng479 <= n1844_1;
    Ng480 <= n1849_1;
    Ng484 <= n1854;
    Ng464 <= n1859_1;
    Ng11517 <= n1864_1;
    Ng11513 <= n1868_1;
    Ng11514 <= n1872_1;
    Ng528 <= n1876_1;
    Ng535 <= n1880_1;
    Ng542 <= n1884_1;
    Ng543 <= n1889_1;
    Ng544 <= n1893_1;
    Ng548 <= n1898_1;
    Ng549 <= n1903;
    Ng8284 <= n1907_1;
    Ng558 <= n1912_1;
    Ng559 <= n1916_1;
    Ng576 <= n1921;
    Ng577 <= n1926_1;
    Ng575 <= n1931;
    Ng579 <= n1936_1;
    Ng580 <= n1941_1;
    Ng578 <= n1946_1;
    Ng582 <= n1951_1;
    Ng583 <= n1956_1;
    Ng581 <= n1961;
    Ng585 <= n1966_1;
    Ng586 <= n1971;
    Ng584 <= n1976_1;
    Ng587 <= n1981;
    Ng590 <= n1986;
    Ng593 <= n1991_1;
    Ng596 <= n1996_1;
    Ng599 <= n2001;
    Ng602 <= n2006_1;
    Ng614 <= n2011_1;
    Ng617 <= n2016;
    Ng620 <= n2021_1;
    Ng605 <= n2026_1;
    Ng608 <= n2031_1;
    Ng611 <= n2036_1;
    Ng490 <= n2041_1;
    Ng493 <= n2046;
    Ng496 <= n2051_1;
    Ng506 <= n2055_1;
    Ng507 <= n2060_1;
    Pg16297 <= n2065;
    Ng525 <= n2068_1;
    Ng529 <= n2073;
    Ng530 <= n2078_1;
    Ng531 <= n2083_1;
    Ng532 <= n2088_1;
    Ng533 <= n2093_1;
    Ng534 <= n2098;
    Ng536 <= n2103;
    Ng537 <= n2108_1;
    Ng538 <= n2113_1;
    Ng541 <= n2118;
    Ng630 <= n2123_1;
    Ng659 <= n2128;
    Ng640 <= n2133;
    Ng633 <= n2138_1;
    Ng653 <= n2143_1;
    Ng646 <= n2148_1;
    Ng660 <= n2153_1;
    Ng672 <= n2158_1;
    Ng666 <= n2163_1;
    Ng679 <= n2168_1;
    Ng686 <= n2173_1;
    Ng692 <= n2178_1;
    Ng699 <= n2183_1;
    Ng700 <= n2188;
    Ng698 <= n2193;
    Ng702 <= n2198_1;
    Ng703 <= n2203_1;
    Ng701 <= n2208_1;
    Ng705 <= n2213;
    Ng706 <= n2218;
    Ng704 <= n2223_1;
    Ng708 <= n2228;
    Ng709 <= n2233_1;
    Ng707 <= n2238;
    Ng711 <= n2243_1;
    Ng712 <= n2248;
    Ng710 <= n2253_1;
    Ng714 <= n2258;
    Ng715 <= n2263;
    Ng713 <= n2268;
    Ng717 <= n2273;
    Ng718 <= n2278_1;
    Ng716 <= n2283;
    Ng720 <= n2288;
    Ng721 <= n2293;
    Ng719 <= n2298;
    Ng723 <= n2303;
    Ng724 <= n2308;
    Ng722 <= n2313;
    Ng726 <= n2318;
    Ng727 <= n2323_1;
    Ng725 <= n2328;
    Ng729 <= n2333;
    Ng730 <= n2338;
    Ng728 <= n2343;
    Ng732 <= n2348;
    Ng733 <= n2353;
    Ng731 <= n2358_1;
    Ng735 <= n2363;
    Ng736 <= n2368;
    Ng734 <= n2373;
    Ng738 <= n2378;
    Ng739 <= n2383;
    Ng737 <= n2388;
    \[1612]  <= n2392;
    \[1594]  <= n2396_1;
    Ng853 <= n2400_1;
    Ng818 <= n2405;
    Ng819 <= n2410;
    Ng817 <= n2415;
    Ng821 <= n2420;
    Ng822 <= n2425_1;
    Ng820 <= n2430_1;
    Ng830 <= n2435;
    Ng831 <= n2440;
    Ng829 <= n2445;
    Ng833 <= n2450_1;
    Ng834 <= n2455_1;
    Ng832 <= n2460_1;
    Ng836 <= n2465;
    Ng837 <= n2470;
    Ng835 <= n2475;
    Ng839 <= n2480;
    Ng840 <= n2485;
    Ng838 <= n2490;
    Ng842 <= n2495_1;
    Ng843 <= n2500_1;
    Ng841 <= n2505_1;
    Ng845 <= n2510_1;
    Ng846 <= n2515_1;
    Ng844 <= n2520_1;
    Ng848 <= n2525;
    Ng849 <= n2530;
    Ng847 <= n2535;
    Ng851 <= n2540;
    Ng852 <= n2545_1;
    Ng850 <= n2550;
    Ng857 <= n2555;
    Ng858 <= n2560_1;
    Ng856 <= n2565;
    Ng860 <= n2570;
    Ng861 <= n2575_1;
    Ng859 <= n2580;
    Ng863 <= n2585;
    Ng864 <= n2590;
    Ng862 <= n2595_1;
    Ng866 <= n2600;
    Ng867 <= n2605;
    Ng865 <= n2610;
    Ng873 <= n2615;
    Ng876 <= n2620_1;
    Ng879 <= n2625;
    Ng918 <= n2630;
    Ng921 <= n2635;
    Ng924 <= n2640;
    Ng882 <= n2645;
    Ng885 <= n2650;
    Ng888 <= n2655;
    Ng927 <= n2660;
    Ng930 <= n2665;
    Ng933 <= n2670;
    Ng891 <= n2675;
    Ng894 <= n2680_1;
    Ng897 <= n2685;
    Ng936 <= n2690;
    Ng939 <= n2695_1;
    Ng942 <= n2700;
    Ng900 <= n2705_1;
    Ng903 <= n2710_1;
    Ng906 <= n2715_1;
    Ng945 <= n2720;
    Ng948 <= n2725_1;
    Ng951 <= n2730_1;
    Ng909 <= n2735_1;
    Ng912 <= n2740_1;
    Ng915 <= n2745_1;
    Ng954 <= n2750_1;
    Ng957 <= n2755_1;
    Ng960 <= n2760_1;
    Ng780 <= n2765_1;
    Ng776 <= n2770_1;
    Ng771 <= n2775_1;
    Ng767 <= n2780_1;
    Ng762 <= n2785_1;
    Ng758 <= n2790_1;
    Ng753 <= n2795_1;
    Ng749 <= n2800_1;
    Ng744 <= n2805_1;
    Ng740 <= n2810_1;
    Ng11524 <= n2815_1;
    Ng11525 <= n2820_1;
    Ng11526 <= n2825_1;
    Ng11527 <= n2830_1;
    Ng11528 <= n2835;
    Ng11529 <= n2840_1;
    Ng11530 <= n2845_1;
    Ng11531 <= n2850_1;
    Ng11532 <= n2855_1;
    Ng11533 <= n2860_1;
    Ng11534 <= n2865_1;
    Ng11535 <= n2870_1;
    Ng1095 <= n2875_1;
    Ng1098 <= n2880_1;
    Ng1101 <= n2885_1;
    Ng1104 <= n2890_1;
    Ng1107 <= n2895_1;
    Ng1110 <= n2900_1;
    Ng1114 <= n2905_1;
    Ng1115 <= n2910_1;
    Ng1113 <= n2915_1;
    Ng1116 <= n2920_1;
    Ng1119 <= n2925_1;
    Ng1122 <= n2930_1;
    Ng1125 <= n2935_1;
    Ng1128 <= n2940_1;
    Ng1131 <= n2945_1;
    Ng1135 <= n2950_1;
    Ng1136 <= n2955_1;
    Ng1134 <= n2960_1;
    Ng999 <= n2965_1;
    Ng1000 <= n2970_1;
    Ng1001 <= n2975_1;
    Ng1002 <= n2980_1;
    Ng1003 <= n2985_1;
    Ng1004 <= n2990_1;
    Ng1005 <= n2995_1;
    Ng1006 <= n3000_1;
    Ng1007 <= n3005_1;
    Ng1009 <= n3010_1;
    Ng1010 <= n3015;
    Ng1008 <= n3020_1;
    Ng1090 <= n3025;
    Ng1091 <= n3030_1;
    Ng1089 <= n3035_1;
    Ng1137 <= n3040;
    Ng1138 <= n3044_1;
    Ng1139 <= n3049_1;
    Ng1140 <= n3053_1;
    Ng1141 <= n3058_1;
    Ng966 <= n3062_1;
    Ng967 <= n3067_1;
    Ng968 <= n3071_1;
    Ng969 <= n3076_1;
    Ng970 <= n3080_1;
    Ng971 <= n3085_1;
    Ng972 <= n3089_1;
    Ng973 <= n3094_1;
    Ng974 <= n3098_1;
    Ng975 <= n3103_1;
    Ng976 <= n3107;
    Ng977 <= n3111_1;
    Ng978 <= n3115_1;
    Ng986 <= n3120_1;
    Ng992 <= n3125_1;
    Ng985 <= n3130_1;
    Ng1029 <= n3134;
    Ng1036 <= n3138_1;
    Ng1037 <= n3142_1;
    Ng1038 <= n3146_1;
    Ng1039 <= n3150;
    Ng1040 <= n3154_1;
    Ng1044 <= n3158_1;
    Ng1051 <= n3162_1;
    Ng1052 <= n3166;
    Ng1053 <= n3170_1;
    Ng1054 <= n3174_1;
    Ng1055 <= n3178_1;
    Ng1059 <= n3182_1;
    Ng1066 <= n3186_1;
    Ng1067 <= n3190_1;
    Ng1068 <= n3194_1;
    Ng1069 <= n3198_1;
    Ng1070 <= n3202_1;
    Ng1074 <= n3206_1;
    Ng1081 <= n3210_1;
    Ng1082 <= n3214_1;
    Ng1083 <= n3218_1;
    Ng1084 <= n3222_1;
    Ng1011 <= n3226_1;
    Ng1240 <= n3231_1;
    Ng1243 <= n3236_1;
    Ng1196 <= n3241_1;
    Ng1199 <= n3246_1;
    Ng1209 <= n3250_1;
    Ng1210 <= n3254_1;
    Ng1250 <= n3259_1;
    Ng1255 <= n3263_1;
    Ng1256 <= n3268_1;
    Ng1257 <= n3272_1;
    Ng1258 <= n3277_1;
    Ng1259 <= n3281_1;
    Ng1260 <= n3286_1;
    Ng1251 <= n3290_1;
    Ng1252 <= n3295_1;
    Ng1253 <= n3299_1;
    Ng1254 <= n3304_1;
    Ng1176 <= n3308_1;
    Ng1173 <= n3313_1;
    Ng1174 <= n3318_1;
    Ng1175 <= n3323_1;
    Ng11539 <= n3328_1;
    Ng11542 <= n3332_1;
    Ng11543 <= n3336_1;
    Ng1164 <= n3340_1;
    Ng1165 <= n3345_1;
    Ng1166 <= n3350_1;
    Ng1167 <= n3355_1;
    Ng1171 <= n3360_1;
    Ng1151 <= n3365_1;
    Ng11544 <= n3370_1;
    Ng11540 <= n3374_1;
    Ng11541 <= n3378_1;
    Ng1214 <= n3382_1;
    Ng1221 <= n3386_1;
    Ng1228 <= n3390_1;
    Ng1229 <= n3395_1;
    Ng1230 <= n3399_1;
    Ng1234 <= n3404_1;
    Ng1235 <= n3409_1;
    Ng8293 <= n3413_1;
    Ng1244 <= n3418_1;
    Ng1245 <= n3422_1;
    Ng1262 <= n3427_1;
    Ng1263 <= n3432_1;
    Ng1261 <= n3437_1;
    Ng1265 <= n3442_1;
    Ng1266 <= n3447_1;
    Ng1264 <= n3452_1;
    Ng1268 <= n3457_1;
    Ng1269 <= n3462_1;
    Ng1267 <= n3467_1;
    Ng1271 <= n3472_1;
    Ng1272 <= n3477_1;
    Ng1270 <= n3482_1;
    Ng1273 <= n3487_1;
    Ng1276 <= n3492_1;
    Ng1279 <= n3497_1;
    Ng1282 <= n3502_1;
    Ng1285 <= n3507_1;
    Ng1288 <= n3512_1;
    Ng1300 <= n3517_1;
    Ng1303 <= n3522_1;
    Ng1306 <= n3527_1;
    Ng1291 <= n3532_1;
    Ng1294 <= n3537_1;
    Ng1297 <= n3542_1;
    Ng1177 <= n3547_1;
    Ng1180 <= n3552_1;
    Ng1183 <= n3557_1;
    Ng1192 <= n3561_1;
    Ng1193 <= n3566_1;
    Pg16355 <= n3571_1;
    Ng1211 <= n3574_1;
    Ng1215 <= n3579_1;
    Ng1216 <= n3584_1;
    Ng1217 <= n3589_1;
    Ng1218 <= n3594_1;
    Ng1219 <= n3599_1;
    Ng1220 <= n3604_1;
    Ng1222 <= n3609_1;
    Ng1223 <= n3614_1;
    Ng1224 <= n3619_1;
    Ng1227 <= n3624_1;
    \[1605]  <= n3629_1;
    \[1603]  <= n3633_1;
    Ng1315 <= n3637_1;
    Ng1316 <= n3642_1;
    Ng1345 <= n3647_1;
    Ng1326 <= n3652_1;
    Ng1319 <= n3657_1;
    Ng1339 <= n3662_1;
    Ng1332 <= n3667_1;
    Ng1346 <= n3672_1;
    Ng1358 <= n3677_1;
    Ng1352 <= n3682_1;
    Ng1365 <= n3687_1;
    Ng1372 <= n3692_1;
    Ng1378 <= n3697_1;
    Ng1385 <= n3702_1;
    Ng1386 <= n3707_1;
    Ng1384 <= n3712_1;
    Ng1388 <= n3717_1;
    Ng1389 <= n3722_1;
    Ng1387 <= n3727_1;
    Ng1391 <= n3732_1;
    Ng1392 <= n3737_1;
    Ng1390 <= n3742_1;
    Ng1394 <= n3747;
    Ng1395 <= n3752_1;
    Ng1393 <= n3757;
    Ng1397 <= n3762_1;
    Ng1398 <= n3767;
    Ng1396 <= n3772_1;
    Ng1400 <= n3777;
    Ng1401 <= n3782;
    Ng1399 <= n3787_1;
    Ng1403 <= n3792_1;
    Ng1404 <= n3797;
    Ng1402 <= n3802_1;
    Ng1406 <= n3807_1;
    Ng1407 <= n3812;
    Ng1405 <= n3817;
    Ng1409 <= n3822_1;
    Ng1410 <= n3827;
    Ng1408 <= n3832_1;
    Ng1412 <= n3837;
    Ng1413 <= n3842_1;
    Ng1411 <= n3847_1;
    Ng1415 <= n3852_1;
    Ng1416 <= n3857_1;
    Ng1414 <= n3862_1;
    Ng1418 <= n3867;
    Ng1419 <= n3872_1;
    Ng1417 <= n3877_1;
    Ng1421 <= n3882;
    Ng1422 <= n3887;
    Ng1420 <= n3892_1;
    Ng1424 <= n3897_1;
    Ng1425 <= n3902;
    Ng1423 <= n3907_1;
    Ng1512 <= n3912_1;
    Ng1513 <= n3917;
    Ng1511 <= n3922;
    Ng1515 <= n3927;
    Ng1516 <= n3932_1;
    Ng1514 <= n3937;
    Ng1524 <= n3942_1;
    Ng1525 <= n3947;
    Ng1523 <= n3952;
    Ng1527 <= n3957_1;
    Ng1528 <= n3962;
    Ng1526 <= n3967;
    Ng1530 <= n3972;
    Ng1531 <= n3977;
    Ng1529 <= n3982;
    Ng1533 <= n3987;
    Ng1534 <= n3992;
    Ng1532 <= n3997_1;
    Ng1536 <= n4002_1;
    Ng1537 <= n4007_1;
    Ng1535 <= n4012;
    Ng1539 <= n4017;
    Ng1540 <= n4022_1;
    Ng1538 <= n4027;
    Ng1542 <= n4032_1;
    Ng1543 <= n4037_1;
    Ng1541 <= n4042;
    Ng1545 <= n4047;
    Ng1546 <= n4052;
    Ng1544 <= n4057_1;
    Ng1551 <= n4062_1;
    Ng1552 <= n4067;
    Ng1550 <= n4072_1;
    Ng1554 <= n4077;
    Ng1555 <= n4082;
    Ng1553 <= n4087;
    Ng1557 <= n4092;
    Ng1558 <= n4097;
    Ng1556 <= n4102_1;
    Ng1560 <= n4107_1;
    Ng1561 <= n4112_1;
    Ng1559 <= n4117;
    Ng1567 <= n4122_1;
    Ng1570 <= n4127_1;
    Ng1573 <= n4132_1;
    Ng1612 <= n4137_1;
    Ng1615 <= n4142_1;
    Ng1618 <= n4147_1;
    Ng1576 <= n4152;
    Ng1579 <= n4157;
    Ng1582 <= n4162;
    Ng1621 <= n4167_1;
    Ng1624 <= n4172;
    Ng1627 <= n4177;
    Ng1585 <= n4182;
    Ng1588 <= n4187_1;
    Ng1591 <= n4192;
    Ng1630 <= n4197_1;
    Ng1633 <= n4202;
    Ng1636 <= n4207;
    Ng1594 <= n4212_1;
    Ng1597 <= n4217_1;
    Ng1600 <= n4222;
    Ng1639 <= n4227;
    Ng1642 <= n4232;
    Ng1645 <= n4237;
    Ng1603 <= n4242;
    Ng1606 <= n4247;
    Ng1609 <= n4252_1;
    Ng1648 <= n4257_1;
    Ng1651 <= n4262;
    Ng1654 <= n4267;
    Ng1466 <= n4272;
    Ng1462 <= n4277;
    Ng1457 <= n4282;
    Ng1453 <= n4287;
    Ng1448 <= n4292;
    Ng1444 <= n4297;
    Ng1439 <= n4302;
    Ng1435 <= n4307;
    Ng1430 <= n4312;
    Ng1426 <= n4317;
    Ng11551 <= n4322_1;
    Ng11552 <= n4327;
    Ng11553 <= n4332_1;
    Ng11554 <= n4337_1;
    Ng11555 <= n4342;
    Ng11556 <= n4347_1;
    Ng11557 <= n4352_1;
    Ng11558 <= n4357_1;
    Ng11559 <= n4362_1;
    Ng11560 <= n4367;
    Ng11561 <= n4372;
    Ng11562 <= n4377;
    Ng1789 <= n4382;
    Ng1792 <= n4387;
    Ng1795 <= n4392;
    Ng1798 <= n4397;
    Ng1801 <= n4402;
    Ng1804 <= n4407;
    Ng1808 <= n4412;
    Ng1809 <= n4417;
    Ng1807 <= n4422;
    Ng1810 <= n4427;
    Ng1813 <= n4432;
    Ng1816 <= n4437;
    Ng1819 <= n4442_1;
    Ng1822 <= n4447_1;
    Ng1825 <= n4452_1;
    Ng1829 <= n4457;
    Ng1830 <= n4462;
    Ng1828 <= n4467;
    Ng1693 <= n4472;
    Ng1694 <= n4477;
    Ng1695 <= n4482;
    Ng1696 <= n4487;
    Ng1697 <= n4492;
    Ng1698 <= n4497;
    Ng1699 <= n4502;
    Ng1700 <= n4507;
    Ng1701 <= n4512;
    Ng1703 <= n4517;
    Ng1704 <= n4522;
    Ng1702 <= n4527;
    Ng1784 <= n4532;
    Ng1785 <= n4537;
    Ng1783 <= n4542;
    Ng1831 <= n4547;
    Ng1832 <= n4551;
    Ng1833 <= n4556;
    Ng1834 <= n4560;
    Ng1835 <= n4565;
    Ng1660 <= n4569;
    Ng1661 <= n4574;
    Ng1662 <= n4578;
    Ng1663 <= n4583;
    Ng1664 <= n4587;
    Ng1665 <= n4592;
    Ng1666 <= n4596;
    Ng1667 <= n4601;
    Ng1668 <= n4605;
    Ng1669 <= n4610;
    Ng1670 <= n4614;
    Ng1671 <= n4618;
    Ng1672 <= n4622;
    Ng1680 <= n4627;
    Ng1686 <= n4632;
    Ng1679 <= n4637;
    Ng1723 <= n4641;
    Ng1730 <= n4645;
    Ng1731 <= n4649;
    Ng1732 <= n4653;
    Ng1733 <= n4657;
    Ng1734 <= n4661;
    Ng1738 <= n4665;
    Ng1745 <= n4669;
    Ng1746 <= n4673;
    Ng1747 <= n4677;
    Ng1748 <= n4681;
    Ng1749 <= n4685;
    Ng1753 <= n4689;
    Ng1760 <= n4693;
    Ng1761 <= n4697;
    Ng1762 <= n4701;
    Ng1763 <= n4705;
    Ng1764 <= n4709;
    Ng1768 <= n4713;
    Ng1775 <= n4717;
    Ng1776 <= n4721;
    Ng1777 <= n4725;
    Ng1778 <= n4729;
    Ng1705 <= n4733;
    Ng1934 <= n4738;
    Ng1937 <= n4743;
    Ng1890 <= n4748;
    Ng1893 <= n4753;
    Ng1903 <= n4757;
    Ng1904 <= n4761;
    Ng1944 <= n4766;
    Ng1949 <= n4770;
    Ng1950 <= n4775;
    Ng1951 <= n4779;
    Ng1952 <= n4784;
    Ng1953 <= n4788;
    Ng1954 <= n4793;
    Ng1945 <= n4797;
    Ng1946 <= n4802;
    Ng1947 <= n4806;
    Ng1948 <= n4811;
    Ng1870 <= n4815;
    Ng1867 <= n4820;
    Ng1868 <= n4825;
    Ng1869 <= n4830;
    Ng11566 <= n4835;
    Ng11569 <= n4839;
    Ng11570 <= n4843;
    Ng1858 <= n4847;
    Ng1859 <= n4852;
    Ng1860 <= n4857;
    Ng1861 <= n4862;
    Ng1865 <= n4867;
    Ng1845 <= n4872_1;
    Ng11571 <= n4877;
    Ng11567 <= n4881;
    Ng11568 <= n4885;
    Ng1908 <= n4889;
    Ng1915 <= n4893_1;
    Ng1922 <= n4897_1;
    Ng1923 <= n4902;
    Ng1924 <= n4906_1;
    Ng1928 <= n4911;
    Ng1929 <= n4916;
    Ng8302 <= n4920;
    Ng1938 <= n4925;
    Ng1939 <= n4929;
    Ng1956 <= n4934;
    Ng1957 <= n4939;
    Ng1955 <= n4944;
    Ng1959 <= n4949;
    Ng1960 <= n4954;
    Ng1958 <= n4959;
    Ng1962 <= n4964;
    Ng1963 <= n4969;
    Ng1961 <= n4974;
    Ng1965 <= n4979;
    Ng1966 <= n4984;
    Ng1964 <= n4989;
    Ng1967 <= n4994;
    Ng1970 <= n4999;
    Ng1973 <= n5004;
    Ng1976 <= n5009;
    Ng1979 <= n5014;
    Ng1982 <= n5019;
    Ng1994 <= n5024;
    Ng1997 <= n5029;
    Ng2000 <= n5034;
    Ng1985 <= n5039;
    Ng1988 <= n5044;
    Ng1991 <= n5049;
    Ng1871 <= n5054;
    Ng1874 <= n5059;
    Ng1877 <= n5064;
    Ng1886 <= n5068;
    Ng1887 <= n5073;
    Pg16399 <= n5078;
    Ng1905 <= n5081;
    Ng1909 <= n5086;
    Ng1910 <= n5091;
    Ng1911 <= n5096;
    Ng1912 <= n5101;
    Ng1913 <= n5106;
    Ng1914 <= n5111;
    Ng1916 <= n5116;
    Ng1917 <= n5121;
    Ng1918 <= n5126;
    Ng1921 <= n5131;
    Ng2010 <= n5136;
    Ng2039 <= n5141;
    Ng2020 <= n5146;
    Ng2013 <= n5151;
    Ng2033 <= n5156;
    Ng2026 <= n5161;
    Ng2040 <= n5166;
    Ng2052 <= n5171;
    Ng2046 <= n5176;
    Ng2059 <= n5181;
    Ng2066 <= n5186;
    Ng2072 <= n5191;
    Ng2079 <= n5196;
    Ng2080 <= n5201;
    Ng2078 <= n5206;
    Ng2082 <= n5211;
    Ng2083 <= n5216;
    Ng2081 <= n5221;
    Ng2085 <= n5226;
    Ng2086 <= n5231;
    Ng2084 <= n5236;
    Ng2088 <= n5241;
    Ng2089 <= n5246;
    Ng2087 <= n5251;
    Ng2091 <= n5256;
    Ng2092 <= n5261;
    Ng2090 <= n5266;
    Ng2094 <= n5271;
    Ng2095 <= n5276;
    Ng2093 <= n5281;
    Ng2097 <= n5286;
    Ng2098 <= n5291;
    Ng2096 <= n5296;
    Ng2100 <= n5301;
    Ng2101 <= n5306;
    Ng2099 <= n5311;
    Ng2103 <= n5316;
    Ng2104 <= n5321;
    Ng2102 <= n5326;
    Ng2106 <= n5331;
    Ng2107 <= n5336;
    Ng2105 <= n5341;
    Ng2109 <= n5346;
    Ng2110 <= n5351;
    Ng2108 <= n5356;
    Ng2112 <= n5361;
    Ng2113 <= n5366;
    Ng2111 <= n5371;
    Ng2115 <= n5376;
    Ng2116 <= n5381;
    Ng2114 <= n5386;
    Ng2118 <= n5391;
    Ng2119 <= n5396;
    Ng2117 <= n5401;
    Ng2206 <= n5406;
    Ng2207 <= n5411;
    Ng2205 <= n5416;
    Ng2209 <= n5421;
    Ng2210 <= n5426;
    Ng2208 <= n5431;
    Ng2218 <= n5436;
    Ng2219 <= n5441;
    Ng2217 <= n5446;
    Ng2221 <= n5451;
    Ng2222 <= n5456;
    Ng2220 <= n5461;
    Ng2224 <= n5466;
    Ng2225 <= n5471;
    Ng2223 <= n5476;
    Ng2227 <= n5481;
    Ng2228 <= n5486;
    Ng2226 <= n5491;
    Ng2230 <= n5496;
    Ng2231 <= n5501;
    Ng2229 <= n5506;
    Ng2233 <= n5511;
    Ng2234 <= n5516;
    Ng2232 <= n5521;
    Ng2236 <= n5526;
    Ng2237 <= n5531;
    Ng2235 <= n5536;
    Ng2239 <= n5541;
    Ng2240 <= n5546;
    Ng2238 <= n5551;
    Ng2245 <= n5556;
    Ng2246 <= n5561;
    Ng2244 <= n5566;
    Ng2248 <= n5571;
    Ng2249 <= n5576;
    Ng2247 <= n5581;
    Ng2251 <= n5586;
    Ng2252 <= n5591;
    Ng2250 <= n5596;
    Ng2254 <= n5601;
    Ng2255 <= n5606;
    Ng2253 <= n5611;
    Ng2261 <= n5616;
    Ng2264 <= n5621;
    Ng2267 <= n5626;
    Ng2306 <= n5631;
    Ng2309 <= n5636;
    Ng2312 <= n5641;
    Ng2270 <= n5646;
    Ng2273 <= n5651;
    Ng2276 <= n5656;
    Ng2315 <= n5661;
    Ng2318 <= n5666;
    Ng2321 <= n5671;
    Ng2279 <= n5676;
    Ng2282 <= n5681;
    Ng2285 <= n5686;
    Ng2324 <= n5691;
    Ng2327 <= n5696;
    Ng2330 <= n5701;
    Ng2288 <= n5706;
    Ng2291 <= n5711;
    Ng2294 <= n5716;
    Ng2333 <= n5721;
    Ng2336 <= n5726;
    Ng2339 <= n5731;
    Ng2297 <= n5736;
    Ng2300 <= n5741;
    Ng2303 <= n5746;
    Ng2342 <= n5751;
    Ng2345 <= n5756;
    Ng2348 <= n5761;
    Ng2160 <= n5766;
    Ng2156 <= n5771;
    Ng2151 <= n5776;
    Ng2147 <= n5781;
    Ng2142 <= n5786;
    Ng2138 <= n5791;
    Ng2133 <= n5796;
    Ng2129 <= n5801;
    Ng2124 <= n5806;
    Ng2120 <= n5811;
    Ng2256 <= n5816;
    \[1609]  <= n5820;
    Ng2257 <= n5824;
    Ng11578 <= n5829;
    Ng11579 <= n5834;
    Ng11580 <= n5839;
    Ng11581 <= n5844;
    Ng11582 <= n5849;
    Ng11583 <= n5854;
    Ng11584 <= n5859;
    Ng11585 <= n5864;
    Ng11586 <= n5869;
    Ng11587 <= n5874;
    Ng11588 <= n5879;
    Ng11589 <= n5884;
    Ng2483 <= n5889;
    Ng2486 <= n5894;
    Ng2489 <= n5899;
    Ng2492 <= n5904;
    Ng2495 <= n5909;
    Ng2498 <= n5914;
    Ng2502 <= n5919;
    Ng2503 <= n5924;
    Ng2501 <= n5929;
    Ng2504 <= n5934;
    Ng2507 <= n5939;
    Ng2510 <= n5944;
    Ng2513 <= n5949;
    Ng2516 <= n5954;
    Ng2519 <= n5959;
    Ng2523 <= n5964;
    Ng2524 <= n5969;
    Ng2522 <= n5974;
    Ng2387 <= n5979;
    Ng2388 <= n5984;
    Ng2389 <= n5989;
    Ng2390 <= n5994;
    Ng2391 <= n5999;
    Ng2392 <= n6004;
    Ng2393 <= n6009;
    Ng2394 <= n6014;
    Ng2395 <= n6019;
    Ng2397 <= n6024;
    Ng2398 <= n6029;
    Ng2396 <= n6034;
    Ng2478 <= n6039;
    Ng2479 <= n6044;
    Ng2477 <= n6049;
    Ng2525 <= n6054;
    Ng2526 <= n6058;
    Ng2527 <= n6063;
    Ng2528 <= n6067;
    Ng2529 <= n6072;
    Ng2354 <= n6076;
    Ng2355 <= n6081;
    Ng2356 <= n6085;
    Ng2357 <= n6090;
    Ng2358 <= n6094;
    Ng2359 <= n6099;
    Ng2360 <= n6103;
    Ng2361 <= n6108;
    Ng2362 <= n6112;
    Ng2363 <= n6117;
    Ng2364 <= n6121;
    Ng2365 <= n6125;
    Ng2366 <= n6129;
    Ng2374 <= n6134;
    Ng2380 <= n6139;
    Ng2373 <= n6144;
    Ng2417 <= n6148;
    Ng2424 <= n6152;
    Ng2425 <= n6156;
    Ng2426 <= n6160;
    Ng2427 <= n6164;
    Ng2428 <= n6168;
    Ng2432 <= n6172;
    Ng2439 <= n6176;
    Ng2440 <= n6180;
    Ng2441 <= n6184;
    Ng2442 <= n6188;
    Ng2443 <= n6192;
    Ng2447 <= n6196;
    Ng2454 <= n6200;
    Ng2455 <= n6204;
    Ng2456 <= n6208;
    Ng2457 <= n6212;
    Ng2458 <= n6216;
    Ng2462 <= n6220;
    Ng2469 <= n6224;
    Ng2470 <= n6228;
    Ng2471 <= n6232;
    Ng2472 <= n6236;
    Ng2399 <= n6240;
    Ng2628 <= n6245;
    Ng2631 <= n6250;
    Ng2584 <= n6255;
    Ng2587 <= n6260;
    Ng2597 <= n6264;
    Ng2598 <= n6268;
    Ng2638 <= n6273;
    Ng2643 <= n6277;
    Ng2644 <= n6282;
    Ng2645 <= n6286;
    Ng2646 <= n6291;
    Ng2647 <= n6295;
    Ng2648 <= n6300;
    Ng2639 <= n6304;
    Ng2640 <= n6309;
    Ng2641 <= n6313;
    Ng2642 <= n6318;
    Ng2564 <= n6322;
    Ng2561 <= n6327;
    Ng2562 <= n6332;
    Ng2563 <= n6337;
    Ng11593 <= n6342;
    Ng11596 <= n6346;
    Ng11597 <= n6350;
    Ng2552 <= n6354;
    Ng2553 <= n6359;
    Ng2554 <= n6364;
    Ng2555 <= n6369;
    Ng2559 <= n6374;
    Ng2539 <= n6379;
    Ng11598 <= n6384;
    Ng11594 <= n6388;
    Ng11595 <= n6392;
    Ng2602 <= n6396;
    Ng2609 <= n6400;
    Ng2616 <= n6404;
    Ng2617 <= n6409;
    Ng2618 <= n6413;
    Ng2622 <= n6418;
    Ng2623 <= n6423;
    Ng8311 <= n6427;
    Ng2632 <= n6432;
    Ng2633 <= n6436;
    Ng2650 <= n6441;
    Ng2651 <= n6446;
    Ng2649 <= n6451;
    Ng2653 <= n6456;
    Ng2654 <= n6461;
    Ng2652 <= n6466;
    Ng2656 <= n6471;
    Ng2657 <= n6476;
    Ng2655 <= n6481;
    Ng2659 <= n6486;
    Ng2660 <= n6491;
    Ng2658 <= n6496;
    Ng2661 <= n6501;
    Ng2664 <= n6506;
    Ng2667 <= n6511;
    Ng2670 <= n6516;
    Ng2673 <= n6521;
    Ng2676 <= n6526;
    Ng2688 <= n6531;
    Ng2691 <= n6536;
    Ng2694 <= n6541;
    Ng2679 <= n6546;
    Ng2682 <= n6551;
    Ng2685 <= n6556;
    Ng2565 <= n6561;
    Ng2568 <= n6566;
    Ng2571 <= n6571;
    Ng2580 <= n6575;
    Ng2581 <= n6580;
    Pg16437 <= n6585;
    Ng2599 <= n6588;
    Ng2603 <= n6593;
    Ng2604 <= n6598;
    Ng2605 <= n6603;
    Ng2606 <= n6608;
    Ng2607 <= n6613;
    Ng2608 <= n6618;
    Ng2610 <= n6623;
    Ng2611 <= n6628;
    Ng2612 <= n6633;
    Ng2615 <= n6638;
    Ng2704 <= n6643;
    Ng2733 <= n6648;
    Ng2714 <= n6653;
    Ng2707 <= n6658;
    Ng2727 <= n6663;
    Ng2720 <= n6668;
    Ng2734 <= n6673;
    Ng2746 <= n6678;
    Ng2740 <= n6683;
    Ng2753 <= n6688;
    Ng2760 <= n6693;
    Ng2766 <= n6698;
    Ng2773 <= n6703;
    Ng2774 <= n6708;
    Ng2772 <= n6713;
    Ng2776 <= n6718;
    Ng2777 <= n6723;
    Ng2775 <= n6728;
    Ng2779 <= n6733;
    Ng2780 <= n6738;
    Ng2778 <= n6743;
    Ng2782 <= n6748;
    Ng2783 <= n6753;
    Ng2781 <= n6758;
    Ng2785 <= n6763;
    Ng2786 <= n6768;
    Ng2784 <= n6773;
    Ng2788 <= n6778;
    Ng2789 <= n6783;
    Ng2787 <= n6788;
    Ng2791 <= n6793;
    Ng2792 <= n6798;
    Ng2790 <= n6803;
    Ng2794 <= n6808;
    Ng2795 <= n6813;
    Ng2793 <= n6818;
    Ng2797 <= n6823;
    Ng2798 <= n6828;
    Ng2796 <= n6833;
    Ng2800 <= n6838;
    Ng2801 <= n6843;
    Ng2799 <= n6848;
    Ng2803 <= n6853;
    Ng2804 <= n6858;
    Ng2802 <= n6863;
    Ng2806 <= n6868;
    Ng2807 <= n6873;
    Ng2805 <= n6878;
    Ng2809 <= n6883;
    Ng2810 <= n6888;
    Ng2808 <= n6893;
    Ng2812 <= n6898;
    Ng2813 <= n6903;
    Ng2811 <= n6908;
    Ng3054 <= n6913;
    Ng3079 <= n6918;
    Ng13475 <= n6923;
    Ng3043 <= n6927;
    Ng3044 <= n6932;
    Ng3045 <= n6937;
    Ng3046 <= n6942;
    Ng3047 <= n6947;
    Ng3048 <= n6952;
    Ng3049 <= n6957;
    Ng3050 <= n6962;
    Ng3051 <= n6967;
    Ng3052 <= n6972;
    Ng3053 <= n6977;
    Ng3055 <= n6982;
    Ng3056 <= n6987;
    Ng3057 <= n6992;
    Ng3058 <= n6997;
    Ng3059 <= n7002;
    Ng3060 <= n7007;
    Ng3061 <= n7012;
    Ng3062 <= n7017;
    Ng3063 <= n7022;
    Ng3064 <= n7027;
    Ng3065 <= n7032;
    Ng3066 <= n7037;
    Ng3067 <= n7042;
    Ng3068 <= n7047;
    Ng3069 <= n7052;
    Ng3070 <= n7057;
    Ng3071 <= n7062;
    Ng3072 <= n7067;
    Ng3073 <= n7072;
    Ng3074 <= n7077;
    Ng3075 <= n7082;
    Ng3076 <= n7087;
    Ng3077 <= n7092;
    Ng3078 <= n7097;
    Ng2997 <= n7102;
    Ng2993 <= n7107;
    Ng2998 <= n7112;
    Ng3006 <= n7117;
    Ng3002 <= n7122;
    Ng3013 <= n7127;
    Ng3010 <= n7132;
    Ng3024 <= n7137;
    Ng3018 <= n7142;
    Ng3028 <= n7147;
    Ng3036 <= n7152;
    Ng3032 <= n7157;
    Pg5388 <= n7161;
    Ng2986 <= n7164;
    Ng2987 <= n7168;
    Pg8275 <= n7173;
    Pg8274 <= n7177;
    Pg8273 <= n7181;
    Pg8272 <= n7185;
    Pg8268 <= n7189;
    Pg8269 <= n7193;
    Pg8270 <= n7197;
    Pg8271 <= n7201;
    Ng3083 <= n7205;
    Pg8267 <= n7210;
    Ng2992 <= n7214;
    Pg8266 <= n7219;
    Pg8265 <= n7223;
    Pg8264 <= n7227;
    Pg8262 <= n7231;
    Pg8263 <= n7235;
    Pg8260 <= n7239;
    Pg8261 <= n7243;
    Pg8259 <= n7247;
    Ng2990 <= n7251;
    Ng2991 <= n7256;
    Pg8258 <= n7261;
  end
endmodule


