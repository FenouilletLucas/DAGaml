// Benchmark "frg1" written by ABC on Tue May 16 16:07:49 2017

module frg1 ( 
    c0, a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w,
    x, y, z, a0, b0,
    d0, e0, f0  );
  input  c0, a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0;
  output d0, e0, f0;
  wire n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n579, n580, n581, n582,
    n584, n585, n586, n587;
  assign n32 = ~c & ~r;
  assign n33 = ~v & n32;
  assign n34 = ~z & n33;
  assign n35 = ~q & n34;
  assign n36 = ~y & n35;
  assign n37 = a & n36;
  assign n38 = ~o & n37;
  assign n39 = ~p & n38;
  assign n40 = ~s & n39;
  assign n41 = ~t & n40;
  assign n42 = ~u & n41;
  assign n43 = ~w & n42;
  assign n44 = ~x & n43;
  assign n45 = ~c & e;
  assign n46 = ~r & n45;
  assign n47 = ~v & n46;
  assign n48 = ~z & n47;
  assign n49 = ~q & n48;
  assign n50 = ~y & n49;
  assign n51 = ~o & n50;
  assign n52 = ~p & n51;
  assign n53 = ~s & n52;
  assign n54 = ~t & n53;
  assign n55 = ~u & n54;
  assign n56 = ~w & n55;
  assign n57 = ~x & n56;
  assign n58 = ~q & n33;
  assign n59 = a & n58;
  assign n60 = ~o & n59;
  assign n61 = ~p & n60;
  assign n62 = ~s & n61;
  assign n63 = ~t & n62;
  assign n64 = ~u & n63;
  assign n65 = ~m & n64;
  assign n66 = ~q & n47;
  assign n67 = ~o & n66;
  assign n68 = ~p & n67;
  assign n69 = ~s & n68;
  assign n70 = ~t & n69;
  assign n71 = ~u & n70;
  assign n72 = ~m & n71;
  assign n73 = ~z & n32;
  assign n74 = ~k & n73;
  assign n75 = ~q & n74;
  assign n76 = ~y & n75;
  assign n77 = a & n76;
  assign n78 = ~o & n77;
  assign n79 = ~p & n78;
  assign n80 = ~w & n79;
  assign n81 = ~x & n80;
  assign n82 = ~z & n46;
  assign n83 = ~k & n82;
  assign n84 = ~q & n83;
  assign n85 = ~y & n84;
  assign n86 = ~o & n85;
  assign n87 = ~p & n86;
  assign n88 = ~w & n87;
  assign n89 = ~x & n88;
  assign n90 = ~c & ~h;
  assign n91 = ~r & n90;
  assign n92 = ~v & n91;
  assign n93 = ~z & n92;
  assign n94 = a & n93;
  assign n95 = ~p & n94;
  assign n96 = ~s & n95;
  assign n97 = ~t & n96;
  assign n98 = ~x & n97;
  assign n99 = ~h & n45;
  assign n100 = ~r & n99;
  assign n101 = ~v & n100;
  assign n102 = ~z & n101;
  assign n103 = ~p & n102;
  assign n104 = ~s & n103;
  assign n105 = ~t & n104;
  assign n106 = ~x & n105;
  assign n107 = a & ~c;
  assign n108 = ~o & n107;
  assign n109 = ~p & n108;
  assign n110 = ~s & n109;
  assign n111 = ~t & n110;
  assign n112 = ~w & n111;
  assign n113 = ~x & n112;
  assign n114 = ~i & n113;
  assign n115 = ~o & n45;
  assign n116 = ~p & n115;
  assign n117 = ~s & n116;
  assign n118 = ~t & n117;
  assign n119 = ~w & n118;
  assign n120 = ~x & n119;
  assign n121 = ~i & n120;
  assign n122 = a & n92;
  assign n123 = ~p & n122;
  assign n124 = ~s & n123;
  assign n125 = ~t & n124;
  assign n126 = ~m & n125;
  assign n127 = ~p & n101;
  assign n128 = ~s & n127;
  assign n129 = ~t & n128;
  assign n130 = ~m & n129;
  assign n131 = ~c & ~j;
  assign n132 = ~r & n131;
  assign n133 = ~v & n132;
  assign n134 = ~z & n133;
  assign n135 = ~q & n134;
  assign n136 = ~y & n135;
  assign n137 = a & n136;
  assign n138 = ~u & n137;
  assign n139 = ~j & n45;
  assign n140 = ~r & n139;
  assign n141 = ~v & n140;
  assign n142 = ~z & n141;
  assign n143 = ~q & n142;
  assign n144 = ~y & n143;
  assign n145 = ~u & n144;
  assign n146 = ~m & n111;
  assign n147 = ~i & n146;
  assign n148 = ~m & n118;
  assign n149 = ~i & n148;
  assign n150 = a & n90;
  assign n151 = ~p & n150;
  assign n152 = ~s & n151;
  assign n153 = ~t & n152;
  assign n154 = ~m & n153;
  assign n155 = ~i & n154;
  assign n156 = ~p & n99;
  assign n157 = ~s & n156;
  assign n158 = ~t & n157;
  assign n159 = ~m & n158;
  assign n160 = ~i & n159;
  assign n161 = ~c & ~k;
  assign n162 = a & n161;
  assign n163 = ~o & n162;
  assign n164 = ~p & n163;
  assign n165 = ~w & n164;
  assign n166 = ~x & n165;
  assign n167 = ~i & n166;
  assign n168 = ~k & n45;
  assign n169 = ~o & n168;
  assign n170 = ~p & n169;
  assign n171 = ~w & n170;
  assign n172 = ~x & n171;
  assign n173 = ~i & n172;
  assign n174 = ~x & n153;
  assign n175 = ~i & n174;
  assign n176 = ~x & n158;
  assign n177 = ~i & n176;
  assign n178 = ~q & n133;
  assign n179 = a & n178;
  assign n180 = ~u & n179;
  assign n181 = ~m & n180;
  assign n182 = ~q & n141;
  assign n183 = ~u & n182;
  assign n184 = ~m & n183;
  assign n185 = ~k & n32;
  assign n186 = ~q & n185;
  assign n187 = a & n186;
  assign n188 = ~o & n187;
  assign n189 = ~p & n188;
  assign n190 = ~m & n189;
  assign n191 = ~k & n46;
  assign n192 = ~q & n191;
  assign n193 = ~o & n192;
  assign n194 = ~p & n193;
  assign n195 = ~m & n194;
  assign n196 = ~z & n91;
  assign n197 = ~k & n196;
  assign n198 = a & n197;
  assign n199 = ~p & n198;
  assign n200 = ~x & n199;
  assign n201 = ~z & n100;
  assign n202 = ~k & n201;
  assign n203 = ~p & n202;
  assign n204 = ~x & n203;
  assign n205 = ~c & ~g;
  assign n206 = ~q & n205;
  assign n207 = ~y & n206;
  assign n208 = a & n207;
  assign n209 = ~o & n208;
  assign n210 = ~u & n209;
  assign n211 = ~w & n210;
  assign n212 = ~g & n45;
  assign n213 = ~q & n212;
  assign n214 = ~y & n213;
  assign n215 = ~o & n214;
  assign n216 = ~u & n215;
  assign n217 = ~w & n216;
  assign n218 = ~k & n205;
  assign n219 = ~q & n218;
  assign n220 = ~y & n219;
  assign n221 = a & n220;
  assign n222 = ~o & n221;
  assign n223 = ~w & n222;
  assign n224 = ~k & n212;
  assign n225 = ~q & n224;
  assign n226 = ~y & n225;
  assign n227 = ~o & n226;
  assign n228 = ~w & n227;
  assign n229 = ~z & n132;
  assign n230 = ~k & n229;
  assign n231 = ~q & n230;
  assign n232 = ~y & n231;
  assign n233 = a & n232;
  assign n234 = ~z & n140;
  assign n235 = ~k & n234;
  assign n236 = ~q & n235;
  assign n237 = ~y & n236;
  assign n238 = ~c & ~z;
  assign n239 = ~y & n238;
  assign n240 = a & n239;
  assign n241 = ~w & n240;
  assign n242 = ~x & n241;
  assign n243 = ~n & n242;
  assign n244 = ~z & n45;
  assign n245 = ~y & n244;
  assign n246 = ~w & n245;
  assign n247 = ~x & n246;
  assign n248 = ~n & n247;
  assign n249 = ~c & ~v;
  assign n250 = a & n249;
  assign n251 = ~s & n250;
  assign n252 = ~t & n251;
  assign n253 = ~u & n252;
  assign n254 = ~l & n253;
  assign n255 = ~v & n45;
  assign n256 = ~s & n255;
  assign n257 = ~t & n256;
  assign n258 = ~u & n257;
  assign n259 = ~l & n258;
  assign n260 = ~v & n90;
  assign n261 = a & n260;
  assign n262 = ~s & n261;
  assign n263 = ~t & n262;
  assign n264 = ~l & n263;
  assign n265 = ~v & n99;
  assign n266 = ~s & n265;
  assign n267 = ~t & n266;
  assign n268 = ~l & n267;
  assign n269 = ~m & n164;
  assign n270 = ~i & n269;
  assign n271 = ~m & n170;
  assign n272 = ~i & n271;
  assign n273 = ~k & n90;
  assign n274 = a & n273;
  assign n275 = ~p & n274;
  assign n276 = ~m & n275;
  assign n277 = ~i & n276;
  assign n278 = ~k & n99;
  assign n279 = ~p & n278;
  assign n280 = ~m & n279;
  assign n281 = ~i & n280;
  assign n282 = ~x & n275;
  assign n283 = ~i & n282;
  assign n284 = ~x & n279;
  assign n285 = ~i & n284;
  assign n286 = a & n206;
  assign n287 = ~o & n286;
  assign n288 = ~u & n287;
  assign n289 = ~m & n288;
  assign n290 = ~o & n213;
  assign n291 = ~u & n290;
  assign n292 = ~m & n291;
  assign n293 = ~g & n131;
  assign n294 = ~q & n293;
  assign n295 = a & n294;
  assign n296 = ~u & n295;
  assign n297 = ~m & n296;
  assign n298 = ~g & n139;
  assign n299 = ~q & n298;
  assign n300 = ~u & n299;
  assign n301 = ~m & n300;
  assign n302 = ~k & n91;
  assign n303 = a & n302;
  assign n304 = ~p & n303;
  assign n305 = ~m & n304;
  assign n306 = ~k & n100;
  assign n307 = ~p & n306;
  assign n308 = ~m & n307;
  assign n309 = a & n219;
  assign n310 = ~o & n309;
  assign n311 = ~m & n310;
  assign n312 = ~o & n225;
  assign n313 = ~m & n312;
  assign n314 = ~k & n293;
  assign n315 = ~q & n314;
  assign n316 = a & n315;
  assign n317 = ~m & n316;
  assign n318 = ~k & n132;
  assign n319 = ~q & n318;
  assign n320 = a & n319;
  assign n321 = ~m & n320;
  assign n322 = ~j & n90;
  assign n323 = ~r & n322;
  assign n324 = ~k & n323;
  assign n325 = a & n324;
  assign n326 = ~m & n325;
  assign n327 = ~v & n323;
  assign n328 = a & n327;
  assign n329 = ~m & n328;
  assign n330 = ~k & n298;
  assign n331 = ~q & n330;
  assign n332 = ~m & n331;
  assign n333 = ~k & n140;
  assign n334 = ~q & n333;
  assign n335 = ~m & n334;
  assign n336 = ~j & n99;
  assign n337 = ~r & n336;
  assign n338 = ~k & n337;
  assign n339 = ~m & n338;
  assign n340 = ~v & n337;
  assign n341 = ~m & n340;
  assign n342 = ~y & n294;
  assign n343 = a & n342;
  assign n344 = ~u & n343;
  assign n345 = ~y & n299;
  assign n346 = ~u & n345;
  assign n347 = ~y & n315;
  assign n348 = a & n347;
  assign n349 = ~z & n323;
  assign n350 = ~k & n349;
  assign n351 = a & n350;
  assign n352 = ~z & n327;
  assign n353 = a & n352;
  assign n354 = ~y & n331;
  assign n355 = ~z & n337;
  assign n356 = ~k & n355;
  assign n357 = ~z & n340;
  assign n358 = ~w & n107;
  assign n359 = ~x & n358;
  assign n360 = ~i & n359;
  assign n361 = ~n & n360;
  assign n362 = ~w & n45;
  assign n363 = ~x & n362;
  assign n364 = ~i & n363;
  assign n365 = ~n & n364;
  assign n366 = ~x & n150;
  assign n367 = ~i & n366;
  assign n368 = ~n & n367;
  assign n369 = ~x & n99;
  assign n370 = ~i & n369;
  assign n371 = ~n & n370;
  assign n372 = a & n205;
  assign n373 = ~w & n372;
  assign n374 = ~i & n373;
  assign n375 = ~n & n374;
  assign n376 = ~w & n212;
  assign n377 = ~i & n376;
  assign n378 = ~n & n377;
  assign n379 = ~z & n90;
  assign n380 = a & n379;
  assign n381 = ~x & n380;
  assign n382 = ~n & n381;
  assign n383 = ~z & n99;
  assign n384 = ~x & n383;
  assign n385 = ~n & n384;
  assign n386 = ~y & n205;
  assign n387 = a & n386;
  assign n388 = ~w & n387;
  assign n389 = ~n & n388;
  assign n390 = ~y & n212;
  assign n391 = ~w & n390;
  assign n392 = ~n & n391;
  assign n393 = ~y & n293;
  assign n394 = a & n393;
  assign n395 = ~n & n394;
  assign n396 = ~z & n131;
  assign n397 = ~y & n396;
  assign n398 = a & n397;
  assign n399 = ~n & n398;
  assign n400 = ~z & n322;
  assign n401 = a & n400;
  assign n402 = ~n & n401;
  assign n403 = ~y & n298;
  assign n404 = ~n & n403;
  assign n405 = ~z & n139;
  assign n406 = ~y & n405;
  assign n407 = ~n & n406;
  assign n408 = ~z & n336;
  assign n409 = ~n & n408;
  assign n410 = ~s & n107;
  assign n411 = ~t & n410;
  assign n412 = ~i & n411;
  assign n413 = ~l & n412;
  assign n414 = ~s & n45;
  assign n415 = ~t & n414;
  assign n416 = ~i & n415;
  assign n417 = ~l & n416;
  assign n418 = ~v & n131;
  assign n419 = a & n418;
  assign n420 = ~u & n419;
  assign n421 = ~l & n420;
  assign n422 = ~v & n139;
  assign n423 = ~u & n422;
  assign n424 = ~l & n423;
  assign n425 = ~v & n322;
  assign n426 = a & n425;
  assign n427 = ~l & n426;
  assign n428 = ~v & n336;
  assign n429 = ~l & n428;
  assign n430 = ~o & n372;
  assign n431 = ~m & n430;
  assign n432 = ~i & n431;
  assign n433 = ~o & n212;
  assign n434 = ~m & n433;
  assign n435 = ~i & n434;
  assign n436 = ~w & n430;
  assign n437 = ~i & n436;
  assign n438 = ~w & n433;
  assign n439 = ~i & n438;
  assign n440 = ~i & n372;
  assign n441 = ~l & n440;
  assign n442 = ~i & n212;
  assign n443 = ~l & n442;
  assign n444 = ~u & n372;
  assign n445 = ~l & n444;
  assign n446 = ~u & n212;
  assign n447 = ~l & n446;
  assign n448 = ~c & ~e;
  assign n449 = ~a & n448;
  assign n450 = ~c0 & n449;
  assign n451 = ~l & n107;
  assign n452 = ~n & n451;
  assign n453 = ~l & n45;
  assign n454 = ~n & n453;
  assign n455 = ~m & n107;
  assign n456 = ~n & n455;
  assign n457 = ~m & n45;
  assign n458 = ~n & n457;
  assign n459 = ~l & n162;
  assign n460 = ~l & n168;
  assign n461 = a & n131;
  assign n462 = ~i & n461;
  assign n463 = ~i & n139;
  assign n464 = ~g & n90;
  assign n465 = a & n464;
  assign n466 = ~g & n99;
  assign n467 = ~b & c;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n465 & n468;
  assign n470 = ~n463 & n469;
  assign n471 = ~n462 & n470;
  assign n472 = ~n460 & n471;
  assign n473 = ~n459 & n472;
  assign n474 = ~n458 & n473;
  assign n475 = ~n456 & n474;
  assign n476 = ~n454 & n475;
  assign n477 = ~n452 & n476;
  assign n478 = ~n450 & n477;
  assign n479 = ~n447 & n478;
  assign n480 = ~n445 & n479;
  assign n481 = ~n443 & n480;
  assign n482 = ~n441 & n481;
  assign n483 = ~n439 & n482;
  assign n484 = ~n437 & n483;
  assign n485 = ~n435 & n484;
  assign n486 = ~n432 & n485;
  assign n487 = ~n429 & n486;
  assign n488 = ~n427 & n487;
  assign n489 = ~n424 & n488;
  assign n490 = ~n421 & n489;
  assign n491 = ~n417 & n490;
  assign n492 = ~n413 & n491;
  assign n493 = ~n409 & n492;
  assign n494 = ~n407 & n493;
  assign n495 = ~n404 & n494;
  assign n496 = ~n402 & n495;
  assign n497 = ~n399 & n496;
  assign n498 = ~n395 & n497;
  assign n499 = ~n392 & n498;
  assign n500 = ~n389 & n499;
  assign n501 = ~n385 & n500;
  assign n502 = ~n382 & n501;
  assign n503 = ~n378 & n502;
  assign n504 = ~n375 & n503;
  assign n505 = ~n371 & n504;
  assign n506 = ~n368 & n505;
  assign n507 = ~n365 & n506;
  assign n508 = ~n361 & n507;
  assign n509 = ~n357 & n508;
  assign n510 = ~n356 & n509;
  assign n511 = ~n354 & n510;
  assign n512 = ~n353 & n511;
  assign n513 = ~n351 & n512;
  assign n514 = ~n348 & n513;
  assign n515 = ~n346 & n514;
  assign n516 = ~n344 & n515;
  assign n517 = ~n341 & n516;
  assign n518 = ~n339 & n517;
  assign n519 = ~n335 & n518;
  assign n520 = ~n332 & n519;
  assign n521 = ~n329 & n520;
  assign n522 = ~n326 & n521;
  assign n523 = ~n321 & n522;
  assign n524 = ~n317 & n523;
  assign n525 = ~n313 & n524;
  assign n526 = ~n311 & n525;
  assign n527 = ~n308 & n526;
  assign n528 = ~n305 & n527;
  assign n529 = ~n301 & n528;
  assign n530 = ~n297 & n529;
  assign n531 = ~n292 & n530;
  assign n532 = ~n289 & n531;
  assign n533 = ~n285 & n532;
  assign n534 = ~n283 & n533;
  assign n535 = ~n281 & n534;
  assign n536 = ~n277 & n535;
  assign n537 = ~n272 & n536;
  assign n538 = ~n270 & n537;
  assign n539 = ~n268 & n538;
  assign n540 = ~n264 & n539;
  assign n541 = ~n259 & n540;
  assign n542 = ~n254 & n541;
  assign n543 = ~n248 & n542;
  assign n544 = ~n243 & n543;
  assign n545 = ~n237 & n544;
  assign n546 = ~n233 & n545;
  assign n547 = ~n228 & n546;
  assign n548 = ~n223 & n547;
  assign n549 = ~n217 & n548;
  assign n550 = ~n211 & n549;
  assign n551 = ~n204 & n550;
  assign n552 = ~n200 & n551;
  assign n553 = ~n195 & n552;
  assign n554 = ~n190 & n553;
  assign n555 = ~n184 & n554;
  assign n556 = ~n181 & n555;
  assign n557 = ~n177 & n556;
  assign n558 = ~n175 & n557;
  assign n559 = ~n173 & n558;
  assign n560 = ~n167 & n559;
  assign n561 = ~n160 & n560;
  assign n562 = ~n155 & n561;
  assign n563 = ~n149 & n562;
  assign n564 = ~n147 & n563;
  assign n565 = ~n145 & n564;
  assign n566 = ~n138 & n565;
  assign n567 = ~n130 & n566;
  assign n568 = ~n126 & n567;
  assign n569 = ~n121 & n568;
  assign n570 = ~n114 & n569;
  assign n571 = ~n106 & n570;
  assign n572 = ~n98 & n571;
  assign n573 = ~n89 & n572;
  assign n574 = ~n81 & n573;
  assign n575 = ~n72 & n574;
  assign n576 = ~n65 & n575;
  assign n577 = ~n57 & n576;
  assign d0 = n44 | ~n577;
  assign n579 = e & f;
  assign n580 = f & ~a0;
  assign n581 = ~a & ~c;
  assign n582 = ~n580 & n581;
  assign e0 = n579 | ~n582;
  assign n584 = c & ~e;
  assign n585 = ~e & ~b0;
  assign n586 = a & ~e;
  assign n587 = ~n585 & ~n586;
  assign f0 = n584 | ~n587;
endmodule


