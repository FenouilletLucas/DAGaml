// Benchmark "x1" written by ABC on Tue May 16 16:07:53 2017

module x1 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0,
    a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2, i1, i2,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0;
  output a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2, i1,
    i2, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1;
  wire n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n147, n148, n149, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1336, n1337, n1339, n1340, n1341, n1342,
    n1343, n1345, n1346, n1347, n1348, n1349;
  assign n87 = ~j & ~r;
  assign n88 = ~v & n87;
  assign n89 = a0 & n88;
  assign n90 = ~b & r0;
  assign n91 = ~b & f0;
  assign n92 = ~b & a0;
  assign n93 = ~l & a0;
  assign n94 = m & a0;
  assign n95 = n & a0;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~n93 & n96;
  assign n98 = ~n92 & n97;
  assign n99 = ~n91 & n98;
  assign n100 = ~n90 & n99;
  assign a1 = n89 | ~n100;
  assign a2 = f0 | r0;
  assign n103 = ~a & b;
  assign n104 = ~j & n103;
  assign n105 = ~m & n104;
  assign n106 = ~n & n105;
  assign n107 = v & n106;
  assign n108 = ~k & n107;
  assign n109 = l & n108;
  assign n110 = a0 & n109;
  assign n111 = j & n103;
  assign n112 = ~m & n111;
  assign n113 = ~n & n112;
  assign n114 = ~k & n113;
  assign n115 = l & n114;
  assign n116 = a0 & n115;
  assign n117 = k0 & n107;
  assign n118 = c & j;
  assign n119 = ~w & n118;
  assign n120 = g0 & n119;
  assign n121 = o0 & t0;
  assign n122 = ~n120 & ~n121;
  assign n123 = ~n117 & n122;
  assign n124 = ~n116 & n123;
  assign b1 = n110 | ~n124;
  assign n126 = ~a & ~e;
  assign n127 = ~g & n126;
  assign n128 = ~m & n127;
  assign n129 = o & n128;
  assign n130 = p & n129;
  assign n131 = ~u & n130;
  assign n132 = ~v & n131;
  assign n133 = ~w & n132;
  assign n134 = p0 & n133;
  assign n135 = e0 & n133;
  assign n136 = ~m & n126;
  assign n137 = o & n136;
  assign n138 = ~p & n137;
  assign n139 = ~u & n138;
  assign n140 = ~v & n139;
  assign n141 = ~w & n140;
  assign n142 = p0 & n141;
  assign n143 = e0 & n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = ~n135 & n144;
  assign b2 = n134 | ~n145;
  assign n147 = v & b0;
  assign n148 = ~v & b0;
  assign n149 = ~m & n148;
  assign c1 = n147 | n149;
  assign n151 = ~m & ~v;
  assign n152 = ~a & n151;
  assign n153 = ~d & n152;
  assign n154 = ~h & n153;
  assign n155 = d0 & n154;
  assign n156 = ~o & n155;
  assign n157 = ~p & n154;
  assign n158 = d0 & n157;
  assign n159 = v & c0;
  assign n160 = ~v & c0;
  assign n161 = ~m & n160;
  assign n162 = ~n159 & ~n161;
  assign n163 = ~n158 & n162;
  assign d1 = n156 | ~n163;
  assign n165 = ~a & g;
  assign n166 = i & n165;
  assign n167 = ~v & n166;
  assign n168 = q0 & n167;
  assign n169 = ~o & n168;
  assign n170 = ~p & n168;
  assign n171 = ~q & n166;
  assign n172 = ~v & n171;
  assign n173 = q0 & n172;
  assign n174 = ~o & n166;
  assign n175 = p0 & n174;
  assign n176 = ~p & n166;
  assign n177 = p0 & n176;
  assign n178 = p0 & n171;
  assign n179 = ~a & i;
  assign n180 = v & n179;
  assign n181 = p0 & n180;
  assign n182 = ~h0 & ~i0;
  assign n183 = ~z & n182;
  assign n184 = ~y & n183;
  assign n185 = ~n181 & n184;
  assign n186 = ~n178 & n185;
  assign n187 = ~n177 & n186;
  assign n188 = ~n175 & n187;
  assign n189 = ~n173 & n188;
  assign n190 = ~n170 & n189;
  assign d2 = n169 | ~n190;
  assign n192 = d & ~m;
  assign n193 = ~o & n192;
  assign n194 = ~u & n193;
  assign n195 = d0 & n194;
  assign n196 = ~e & n195;
  assign n197 = ~w & n196;
  assign n198 = d & g;
  assign n199 = ~m & n198;
  assign n200 = ~o & n199;
  assign n201 = d0 & n200;
  assign n202 = e & n201;
  assign n203 = u & n200;
  assign n204 = d0 & n203;
  assign n205 = o0 & u0;
  assign n206 = ~m & ~o;
  assign n207 = ~a & n206;
  assign n208 = ~h & n207;
  assign n209 = e0 & n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~n204 & n210;
  assign n212 = ~n202 & n211;
  assign e1 = n197 | ~n212;
  assign n214 = ~y & ~z;
  assign n215 = ~h0 & n214;
  assign n216 = ~i0 & n215;
  assign n217 = ~p0 & n216;
  assign n218 = o & n217;
  assign n219 = p & n218;
  assign n220 = q & n219;
  assign n221 = ~v & n216;
  assign n222 = o & n221;
  assign n223 = p & n222;
  assign n224 = q & n223;
  assign n225 = ~q0 & n217;
  assign n226 = v & n216;
  assign n227 = ~p0 & n226;
  assign n228 = ~g & n216;
  assign n229 = ~p0 & n228;
  assign n230 = ~v & n228;
  assign n231 = ~i & n216;
  assign n232 = a & ~y;
  assign n233 = ~z & n232;
  assign n234 = ~h0 & n233;
  assign n235 = ~i0 & n234;
  assign n236 = ~n231 & ~n235;
  assign n237 = ~n230 & n236;
  assign n238 = ~n229 & n237;
  assign n239 = ~n227 & n238;
  assign n240 = ~n225 & n239;
  assign n241 = ~n224 & n240;
  assign e2 = n220 | ~n241;
  assign n243 = ~a & o;
  assign n244 = ~h & n243;
  assign n245 = ~m & n244;
  assign n246 = p & n245;
  assign n247 = e0 & n246;
  assign n248 = ~q & q0;
  assign n249 = ~i & n248;
  assign n250 = ~o & q0;
  assign n251 = ~i & n250;
  assign n252 = ~g & q0;
  assign n253 = ~q & n252;
  assign n254 = ~g & ~o;
  assign n255 = q0 & n254;
  assign n256 = ~n253 & ~n255;
  assign n257 = ~n251 & n256;
  assign n258 = ~n249 & n257;
  assign f1 = n247 | ~n258;
  assign n260 = ~f0 & ~m0;
  assign n261 = ~p0 & n260;
  assign n262 = ~r0 & n261;
  assign n263 = ~s0 & n262;
  assign n264 = ~x0 & n263;
  assign n265 = d & n264;
  assign n266 = ~e0 & n265;
  assign n267 = ~t & n266;
  assign n268 = b & n267;
  assign n269 = ~j & n268;
  assign n270 = l & n269;
  assign n271 = ~m & n270;
  assign n272 = r & n271;
  assign n273 = ~d0 & ~f0;
  assign n274 = ~m0 & n273;
  assign n275 = ~p0 & n274;
  assign n276 = ~r0 & n275;
  assign n277 = ~s0 & n276;
  assign n278 = ~x0 & n277;
  assign n279 = ~e0 & n278;
  assign n280 = ~t & n279;
  assign n281 = b & n280;
  assign n282 = ~j & n281;
  assign n283 = l & n282;
  assign n284 = ~m & n283;
  assign n285 = r & n284;
  assign n286 = o & ~f0;
  assign n287 = ~m0 & n286;
  assign n288 = ~p0 & n287;
  assign n289 = ~r0 & n288;
  assign n290 = ~s0 & n289;
  assign n291 = ~x0 & n290;
  assign n292 = d & n291;
  assign n293 = ~t & n292;
  assign n294 = b & n293;
  assign n295 = ~j & n294;
  assign n296 = l & n295;
  assign n297 = ~m & n296;
  assign n298 = r & n297;
  assign n299 = o & ~d0;
  assign n300 = ~f0 & n299;
  assign n301 = ~m0 & n300;
  assign n302 = ~p0 & n301;
  assign n303 = ~r0 & n302;
  assign n304 = ~s0 & n303;
  assign n305 = ~x0 & n304;
  assign n306 = ~t & n305;
  assign n307 = b & n306;
  assign n308 = ~j & n307;
  assign n309 = l & n308;
  assign n310 = ~m & n309;
  assign n311 = r & n310;
  assign n312 = ~f0 & ~i0;
  assign n313 = ~m0 & n312;
  assign n314 = ~p0 & n313;
  assign n315 = ~r0 & n314;
  assign n316 = ~s0 & n315;
  assign n317 = ~x0 & n316;
  assign n318 = d & n317;
  assign n319 = ~e0 & n318;
  assign n320 = b & n319;
  assign n321 = ~j & n320;
  assign n322 = l & n321;
  assign n323 = ~m & n322;
  assign n324 = r & n323;
  assign n325 = ~i0 & n273;
  assign n326 = ~m0 & n325;
  assign n327 = ~p0 & n326;
  assign n328 = ~r0 & n327;
  assign n329 = ~s0 & n328;
  assign n330 = ~x0 & n329;
  assign n331 = ~e0 & n330;
  assign n332 = b & n331;
  assign n333 = ~j & n332;
  assign n334 = l & n333;
  assign n335 = ~m & n334;
  assign n336 = r & n335;
  assign n337 = ~i0 & n286;
  assign n338 = ~m0 & n337;
  assign n339 = ~p0 & n338;
  assign n340 = ~r0 & n339;
  assign n341 = ~s0 & n340;
  assign n342 = ~x0 & n341;
  assign n343 = d & n342;
  assign n344 = b & n343;
  assign n345 = ~j & n344;
  assign n346 = l & n345;
  assign n347 = ~m & n346;
  assign n348 = r & n347;
  assign n349 = ~i0 & n300;
  assign n350 = ~m0 & n349;
  assign n351 = ~p0 & n350;
  assign n352 = ~r0 & n351;
  assign n353 = ~s0 & n352;
  assign n354 = ~x0 & n353;
  assign n355 = b & n354;
  assign n356 = ~j & n355;
  assign n357 = l & n356;
  assign n358 = ~m & n357;
  assign n359 = r & n358;
  assign n360 = l & n268;
  assign n361 = z0 & n360;
  assign n362 = l & n281;
  assign n363 = z0 & n362;
  assign n364 = l & n294;
  assign n365 = z0 & n364;
  assign n366 = l & n307;
  assign n367 = z0 & n366;
  assign n368 = l & n320;
  assign n369 = z0 & n368;
  assign n370 = l & n332;
  assign n371 = z0 & n370;
  assign n372 = l & n344;
  assign n373 = z0 & n372;
  assign n374 = l & n355;
  assign n375 = z0 & n374;
  assign n376 = ~r0 & n260;
  assign n377 = ~x0 & n376;
  assign n378 = ~h & n377;
  assign n379 = b & n378;
  assign n380 = ~j & n379;
  assign n381 = l & n380;
  assign n382 = ~m & n381;
  assign n383 = r & n382;
  assign n384 = ~a0 & ~f0;
  assign n385 = ~m0 & n384;
  assign n386 = ~p0 & n385;
  assign n387 = ~r0 & n386;
  assign n388 = ~s0 & n387;
  assign n389 = ~x0 & n388;
  assign n390 = d & n389;
  assign n391 = ~e0 & n390;
  assign n392 = ~t & n391;
  assign n393 = ~a0 & ~d0;
  assign n394 = ~f0 & n393;
  assign n395 = ~m0 & n394;
  assign n396 = ~p0 & n395;
  assign n397 = ~r0 & n396;
  assign n398 = ~s0 & n397;
  assign n399 = ~x0 & n398;
  assign n400 = ~e0 & n399;
  assign n401 = ~t & n400;
  assign n402 = o & ~a0;
  assign n403 = ~f0 & n402;
  assign n404 = ~m0 & n403;
  assign n405 = ~p0 & n404;
  assign n406 = ~r0 & n405;
  assign n407 = ~s0 & n406;
  assign n408 = ~x0 & n407;
  assign n409 = d & n408;
  assign n410 = ~t & n409;
  assign n411 = ~d0 & n402;
  assign n412 = ~f0 & n411;
  assign n413 = ~m0 & n412;
  assign n414 = ~p0 & n413;
  assign n415 = ~r0 & n414;
  assign n416 = ~s0 & n415;
  assign n417 = ~x0 & n416;
  assign n418 = ~t & n417;
  assign n419 = ~i0 & n384;
  assign n420 = ~m0 & n419;
  assign n421 = ~p0 & n420;
  assign n422 = ~r0 & n421;
  assign n423 = ~s0 & n422;
  assign n424 = ~x0 & n423;
  assign n425 = d & n424;
  assign n426 = ~e0 & n425;
  assign n427 = ~i0 & n394;
  assign n428 = ~m0 & n427;
  assign n429 = ~p0 & n428;
  assign n430 = ~r0 & n429;
  assign n431 = ~s0 & n430;
  assign n432 = ~x0 & n431;
  assign n433 = ~e0 & n432;
  assign n434 = ~i0 & n403;
  assign n435 = ~m0 & n434;
  assign n436 = ~p0 & n435;
  assign n437 = ~r0 & n436;
  assign n438 = ~s0 & n437;
  assign n439 = ~x0 & n438;
  assign n440 = d & n439;
  assign n441 = ~i0 & n412;
  assign n442 = ~m0 & n441;
  assign n443 = ~p0 & n442;
  assign n444 = ~r0 & n443;
  assign n445 = ~s0 & n444;
  assign n446 = ~x0 & n445;
  assign n447 = l & n379;
  assign n448 = z0 & n447;
  assign n449 = ~r0 & n385;
  assign n450 = ~x0 & n449;
  assign n451 = ~h & n450;
  assign n452 = ~n448 & ~n451;
  assign n453 = ~n446 & n452;
  assign n454 = ~n440 & n453;
  assign n455 = ~n433 & n454;
  assign n456 = ~n426 & n455;
  assign n457 = ~n418 & n456;
  assign n458 = ~n410 & n457;
  assign n459 = ~n401 & n458;
  assign n460 = ~n392 & n459;
  assign n461 = ~n383 & n460;
  assign n462 = ~n375 & n461;
  assign n463 = ~n373 & n462;
  assign n464 = ~n371 & n463;
  assign n465 = ~n369 & n464;
  assign n466 = ~n367 & n465;
  assign n467 = ~n365 & n466;
  assign n468 = ~n363 & n467;
  assign n469 = ~n361 & n468;
  assign n470 = ~n359 & n469;
  assign n471 = ~n348 & n470;
  assign n472 = ~n336 & n471;
  assign n473 = ~n324 & n472;
  assign n474 = ~n311 & n473;
  assign n475 = ~n298 & n474;
  assign n476 = ~n285 & n475;
  assign f2 = n272 | ~n476;
  assign n478 = ~g & n152;
  assign n479 = ~h & n478;
  assign n480 = ~q & n479;
  assign n481 = p0 & n480;
  assign n482 = ~d & n481;
  assign n483 = ~s & n482;
  assign n484 = ~m & ~p;
  assign n485 = ~v & n484;
  assign n486 = ~a & n485;
  assign n487 = ~g & n486;
  assign n488 = ~h & n487;
  assign n489 = p0 & n488;
  assign n490 = ~d & n489;
  assign n491 = ~s & n490;
  assign n492 = ~v & n206;
  assign n493 = ~a & n492;
  assign n494 = ~g & n493;
  assign n495 = ~h & n494;
  assign n496 = p0 & n495;
  assign n497 = ~d & n496;
  assign n498 = ~s & n497;
  assign n499 = ~c & n152;
  assign n500 = ~g & n499;
  assign n501 = ~h & n500;
  assign n502 = ~q & n501;
  assign n503 = p0 & n502;
  assign n504 = ~s & n503;
  assign n505 = ~c & n486;
  assign n506 = ~g & n505;
  assign n507 = ~h & n506;
  assign n508 = p0 & n507;
  assign n509 = ~s & n508;
  assign n510 = ~c & n493;
  assign n511 = ~g & n510;
  assign n512 = ~h & n511;
  assign n513 = p0 & n512;
  assign n514 = ~s & n513;
  assign n515 = ~r & n480;
  assign n516 = p0 & n515;
  assign n517 = ~d & n516;
  assign n518 = ~r & n488;
  assign n519 = p0 & n518;
  assign n520 = ~d & n519;
  assign n521 = ~r & n495;
  assign n522 = p0 & n521;
  assign n523 = ~d & n522;
  assign n524 = ~r & n502;
  assign n525 = p0 & n524;
  assign n526 = ~r & n507;
  assign n527 = p0 & n526;
  assign n528 = ~r & n512;
  assign n529 = p0 & n528;
  assign n530 = ~h & n165;
  assign n531 = ~q & n530;
  assign n532 = p0 & n531;
  assign n533 = ~i & n532;
  assign n534 = ~s & n533;
  assign n535 = ~a & v;
  assign n536 = ~h & n535;
  assign n537 = ~q & n536;
  assign n538 = p0 & n537;
  assign n539 = ~i & n538;
  assign n540 = ~s & n539;
  assign n541 = ~a & ~p;
  assign n542 = g & n541;
  assign n543 = ~h & n542;
  assign n544 = p0 & n543;
  assign n545 = ~i & n544;
  assign n546 = ~s & n545;
  assign n547 = ~a & ~o;
  assign n548 = g & n547;
  assign n549 = ~h & n548;
  assign n550 = p0 & n549;
  assign n551 = ~i & n550;
  assign n552 = ~s & n551;
  assign n553 = ~p & v;
  assign n554 = ~a & n553;
  assign n555 = ~h & n554;
  assign n556 = p0 & n555;
  assign n557 = ~i & n556;
  assign n558 = ~s & n557;
  assign n559 = ~o & v;
  assign n560 = ~a & n559;
  assign n561 = ~h & n560;
  assign n562 = p0 & n561;
  assign n563 = ~i & n562;
  assign n564 = ~s & n563;
  assign n565 = ~r & n531;
  assign n566 = p0 & n565;
  assign n567 = ~i & n566;
  assign n568 = ~r & n537;
  assign n569 = p0 & n568;
  assign n570 = ~i & n569;
  assign n571 = ~r & n543;
  assign n572 = p0 & n571;
  assign n573 = ~i & n572;
  assign n574 = ~r & n549;
  assign n575 = p0 & n574;
  assign n576 = ~i & n575;
  assign n577 = ~r & n555;
  assign n578 = p0 & n577;
  assign n579 = ~i & n578;
  assign n580 = ~r & n561;
  assign n581 = p0 & n580;
  assign n582 = ~i & n581;
  assign n583 = ~m & o;
  assign n584 = p & n583;
  assign n585 = u & n584;
  assign n586 = ~v & n585;
  assign n587 = d0 & n586;
  assign n588 = g & n587;
  assign n589 = e & ~m;
  assign n590 = o & n589;
  assign n591 = p & n590;
  assign n592 = ~v & n591;
  assign n593 = d0 & n592;
  assign n594 = g & n593;
  assign n595 = ~e & ~m;
  assign n596 = o & n595;
  assign n597 = p & n596;
  assign n598 = ~u & n597;
  assign n599 = ~v & n598;
  assign n600 = d0 & n599;
  assign n601 = o0 & v0;
  assign n602 = v & d0;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n600 & n603;
  assign n605 = ~n594 & n604;
  assign n606 = ~n588 & n605;
  assign n607 = ~n582 & n606;
  assign n608 = ~n579 & n607;
  assign n609 = ~n576 & n608;
  assign n610 = ~n573 & n609;
  assign n611 = ~n570 & n610;
  assign n612 = ~n567 & n611;
  assign n613 = ~n564 & n612;
  assign n614 = ~n558 & n613;
  assign n615 = ~n552 & n614;
  assign n616 = ~n546 & n615;
  assign n617 = ~n540 & n616;
  assign n618 = ~n534 & n617;
  assign n619 = ~n529 & n618;
  assign n620 = ~n527 & n619;
  assign n621 = ~n525 & n620;
  assign n622 = ~n523 & n621;
  assign n623 = ~n520 & n622;
  assign n624 = ~n517 & n623;
  assign n625 = ~n514 & n624;
  assign n626 = ~n509 & n625;
  assign n627 = ~n504 & n626;
  assign n628 = ~n498 & n627;
  assign n629 = ~n491 & n628;
  assign g1 = n483 | ~n629;
  assign n631 = b & a0;
  assign n632 = ~z0 & n631;
  assign n633 = j & n632;
  assign n634 = m & n632;
  assign n635 = ~r & n631;
  assign n636 = ~z0 & n635;
  assign n637 = ~d & h;
  assign n638 = d0 & n637;
  assign n639 = h & ~o;
  assign n640 = e0 & n639;
  assign n641 = h & t;
  assign s1 = i0 & n641;
  assign n643 = b & ~l;
  assign n644 = a0 & n643;
  assign n645 = h & s0;
  assign n646 = h & p0;
  assign n647 = ~x0 & ~a2;
  assign n648 = ~m0 & n647;
  assign n649 = ~n92 & n648;
  assign n650 = ~n646 & n649;
  assign n651 = ~n645 & n650;
  assign n652 = ~n644 & n651;
  assign n653 = ~s1 & n652;
  assign n654 = ~n640 & n653;
  assign n655 = ~n638 & n654;
  assign n656 = ~n636 & n655;
  assign n657 = ~n634 & n656;
  assign g2 = n633 | ~n657;
  assign n659 = h & n126;
  assign n660 = ~u & n659;
  assign n661 = ~w & n660;
  assign n662 = ~o & n661;
  assign n663 = e0 & n662;
  assign n664 = ~d & n661;
  assign n665 = d0 & n664;
  assign n666 = p0 & n661;
  assign n667 = s0 & n661;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~n665 & n668;
  assign h1 = n663 | ~n669;
  assign n671 = ~y & n637;
  assign n672 = ~z & n671;
  assign n673 = ~b0 & n672;
  assign n674 = ~c0 & n673;
  assign n675 = ~h0 & n674;
  assign n676 = ~i0 & n675;
  assign n677 = ~a0 & n676;
  assign n678 = ~g0 & n677;
  assign n679 = ~k0 & n678;
  assign n680 = ~i & n637;
  assign n681 = ~y & n680;
  assign n682 = ~z & n681;
  assign n683 = ~b0 & n682;
  assign n684 = ~c0 & n683;
  assign n685 = ~h0 & n684;
  assign n686 = ~a0 & n685;
  assign n687 = ~g0 & n686;
  assign n688 = ~k0 & n687;
  assign n689 = ~c & n675;
  assign n690 = ~i0 & n689;
  assign n691 = ~a0 & n690;
  assign n692 = ~k0 & n691;
  assign n693 = ~j & n637;
  assign n694 = ~y & n693;
  assign n695 = ~z & n694;
  assign n696 = ~b0 & n695;
  assign n697 = ~c0 & n696;
  assign n698 = ~h0 & n697;
  assign n699 = ~i0 & n698;
  assign n700 = ~a0 & n699;
  assign n701 = ~k0 & n700;
  assign n702 = ~c & n685;
  assign n703 = ~a0 & n702;
  assign n704 = ~k0 & n703;
  assign n705 = ~j & n680;
  assign n706 = ~y & n705;
  assign n707 = ~z & n706;
  assign n708 = ~b0 & n707;
  assign n709 = ~c0 & n708;
  assign n710 = ~h0 & n709;
  assign n711 = ~a0 & n710;
  assign n712 = ~k0 & n711;
  assign n713 = ~v & n678;
  assign n714 = ~v & n687;
  assign n715 = ~v & n691;
  assign n716 = ~v & n703;
  assign n717 = j & n637;
  assign n718 = ~y & n717;
  assign n719 = ~z & n718;
  assign n720 = ~b0 & n719;
  assign n721 = ~c0 & n720;
  assign n722 = ~h0 & n721;
  assign n723 = ~i0 & n722;
  assign n724 = ~a0 & n723;
  assign n725 = ~g0 & n724;
  assign n726 = j & n680;
  assign n727 = ~y & n726;
  assign n728 = ~z & n727;
  assign n729 = ~b0 & n728;
  assign n730 = ~c0 & n729;
  assign n731 = ~h0 & n730;
  assign n732 = ~a0 & n731;
  assign n733 = ~g0 & n732;
  assign n734 = ~c & n722;
  assign n735 = ~i0 & n734;
  assign n736 = ~a0 & n735;
  assign n737 = ~c & n731;
  assign n738 = ~a0 & n737;
  assign n739 = ~b0 & n214;
  assign n740 = ~c0 & n739;
  assign n741 = ~h0 & n740;
  assign n742 = ~d0 & n741;
  assign n743 = ~i0 & n742;
  assign n744 = ~a0 & n743;
  assign n745 = ~g0 & n744;
  assign n746 = ~k0 & n745;
  assign n747 = ~i & ~y;
  assign n748 = ~z & n747;
  assign n749 = ~b0 & n748;
  assign n750 = ~c0 & n749;
  assign n751 = ~h0 & n750;
  assign n752 = ~d0 & n751;
  assign n753 = ~a0 & n752;
  assign n754 = ~g0 & n753;
  assign n755 = ~k0 & n754;
  assign n756 = ~c & n741;
  assign n757 = ~d0 & n756;
  assign n758 = ~i0 & n757;
  assign n759 = ~a0 & n758;
  assign n760 = ~k0 & n759;
  assign n761 = ~j & ~y;
  assign n762 = ~z & n761;
  assign n763 = ~b0 & n762;
  assign n764 = ~c0 & n763;
  assign n765 = ~h0 & n764;
  assign n766 = ~d0 & n765;
  assign n767 = ~i0 & n766;
  assign n768 = ~a0 & n767;
  assign n769 = ~k0 & n768;
  assign n770 = ~c & n751;
  assign n771 = ~d0 & n770;
  assign n772 = ~a0 & n771;
  assign n773 = ~k0 & n772;
  assign n774 = ~i & ~j;
  assign n775 = ~y & n774;
  assign n776 = ~z & n775;
  assign n777 = ~b0 & n776;
  assign n778 = ~c0 & n777;
  assign n779 = ~h0 & n778;
  assign n780 = ~d0 & n779;
  assign n781 = ~a0 & n780;
  assign n782 = ~k0 & n781;
  assign n783 = ~g0 & n676;
  assign n784 = n & n783;
  assign n785 = ~g0 & n685;
  assign n786 = n & n785;
  assign n787 = n & n690;
  assign n788 = n & n699;
  assign n789 = n & n702;
  assign n790 = n & n710;
  assign n791 = m & n783;
  assign n792 = m & n785;
  assign n793 = m & n690;
  assign n794 = m & n699;
  assign n795 = m & n702;
  assign n796 = m & n710;
  assign n797 = a & n783;
  assign n798 = a & n785;
  assign n799 = a & n690;
  assign n800 = a & n699;
  assign n801 = a & n702;
  assign n802 = a & n710;
  assign n803 = ~v & n745;
  assign n804 = ~v & n754;
  assign n805 = ~v & n759;
  assign n806 = ~v & n772;
  assign n807 = ~v & n699;
  assign n808 = ~v & n710;
  assign n809 = j & ~y;
  assign n810 = ~z & n809;
  assign n811 = ~b0 & n810;
  assign n812 = ~c0 & n811;
  assign n813 = ~h0 & n812;
  assign n814 = ~d0 & n813;
  assign n815 = ~i0 & n814;
  assign n816 = ~a0 & n815;
  assign n817 = ~g0 & n816;
  assign n818 = ~i & j;
  assign n819 = ~y & n818;
  assign n820 = ~z & n819;
  assign n821 = ~b0 & n820;
  assign n822 = ~c0 & n821;
  assign n823 = ~h0 & n822;
  assign n824 = ~d0 & n823;
  assign n825 = ~a0 & n824;
  assign n826 = ~g0 & n825;
  assign n827 = ~b & n675;
  assign n828 = ~i0 & n827;
  assign n829 = ~g0 & n828;
  assign n830 = ~l & n637;
  assign n831 = ~y & n830;
  assign n832 = ~z & n831;
  assign n833 = ~b0 & n832;
  assign n834 = ~c0 & n833;
  assign n835 = ~h0 & n834;
  assign n836 = ~i0 & n835;
  assign n837 = ~g0 & n836;
  assign n838 = ~b & n685;
  assign n839 = ~g0 & n838;
  assign n840 = ~l & n680;
  assign n841 = ~y & n840;
  assign n842 = ~z & n841;
  assign n843 = ~b0 & n842;
  assign n844 = ~c0 & n843;
  assign n845 = ~h0 & n844;
  assign n846 = ~g0 & n845;
  assign n847 = ~c & n813;
  assign n848 = ~d0 & n847;
  assign n849 = ~i0 & n848;
  assign n850 = ~a0 & n849;
  assign n851 = ~c & n823;
  assign n852 = ~d0 & n851;
  assign n853 = ~a0 & n852;
  assign n854 = ~c & n827;
  assign n855 = ~i0 & n854;
  assign n856 = ~c & n835;
  assign n857 = ~i0 & n856;
  assign n858 = ~b & n698;
  assign n859 = ~i0 & n858;
  assign n860 = ~l & n693;
  assign n861 = ~y & n860;
  assign n862 = ~z & n861;
  assign n863 = ~b0 & n862;
  assign n864 = ~c0 & n863;
  assign n865 = ~h0 & n864;
  assign n866 = ~i0 & n865;
  assign n867 = ~c & n838;
  assign n868 = ~c & n845;
  assign n869 = ~b & n710;
  assign n870 = ~l & n705;
  assign n871 = ~y & n870;
  assign n872 = ~z & n871;
  assign n873 = ~b0 & n872;
  assign n874 = ~c0 & n873;
  assign n875 = ~h0 & n874;
  assign n876 = ~g0 & n743;
  assign n877 = n & n876;
  assign n878 = ~g0 & n752;
  assign n879 = n & n878;
  assign n880 = n & n758;
  assign n881 = n & n767;
  assign n882 = n & n771;
  assign n883 = n & n780;
  assign n884 = m & n876;
  assign n885 = m & n878;
  assign n886 = m & n758;
  assign n887 = m & n767;
  assign n888 = m & n771;
  assign n889 = m & n780;
  assign n890 = a & n876;
  assign n891 = a & n878;
  assign n892 = a & n758;
  assign n893 = a & n767;
  assign n894 = a & n771;
  assign n895 = a & n780;
  assign n896 = ~v & n767;
  assign n897 = ~v & n780;
  assign n898 = ~b & n741;
  assign n899 = ~d0 & n898;
  assign n900 = ~i0 & n899;
  assign n901 = ~g0 & n900;
  assign n902 = ~l & ~y;
  assign n903 = ~z & n902;
  assign n904 = ~b0 & n903;
  assign n905 = ~c0 & n904;
  assign n906 = ~h0 & n905;
  assign n907 = ~d0 & n906;
  assign n908 = ~i0 & n907;
  assign n909 = ~g0 & n908;
  assign n910 = ~b & n751;
  assign n911 = ~d0 & n910;
  assign n912 = ~g0 & n911;
  assign n913 = ~i & ~l;
  assign n914 = ~y & n913;
  assign n915 = ~z & n914;
  assign n916 = ~b0 & n915;
  assign n917 = ~c0 & n916;
  assign n918 = ~h0 & n917;
  assign n919 = ~d0 & n918;
  assign n920 = ~g0 & n919;
  assign n921 = ~c & n898;
  assign n922 = ~d0 & n921;
  assign n923 = ~i0 & n922;
  assign n924 = ~c & n906;
  assign n925 = ~d0 & n924;
  assign n926 = ~i0 & n925;
  assign n927 = ~b & n765;
  assign n928 = ~d0 & n927;
  assign n929 = ~i0 & n928;
  assign n930 = ~j & ~l;
  assign n931 = ~y & n930;
  assign n932 = ~z & n931;
  assign n933 = ~b0 & n932;
  assign n934 = ~c0 & n933;
  assign n935 = ~h0 & n934;
  assign n936 = ~d0 & n935;
  assign n937 = ~i0 & n936;
  assign n938 = ~c & n910;
  assign n939 = ~d0 & n938;
  assign n940 = ~c & n918;
  assign n941 = ~d0 & n940;
  assign n942 = ~b & n779;
  assign n943 = ~d0 & n942;
  assign n944 = ~l & n774;
  assign n945 = ~y & n944;
  assign n946 = ~z & n945;
  assign n947 = ~b0 & n946;
  assign n948 = ~c0 & n947;
  assign n949 = ~h0 & n948;
  assign n950 = ~d0 & n949;
  assign n951 = ~n943 & ~n950;
  assign n952 = ~n941 & n951;
  assign n953 = ~n939 & n952;
  assign n954 = ~n937 & n953;
  assign n955 = ~n929 & n954;
  assign n956 = ~n926 & n955;
  assign n957 = ~n923 & n956;
  assign n958 = ~n920 & n957;
  assign n959 = ~n912 & n958;
  assign n960 = ~n909 & n959;
  assign n961 = ~n901 & n960;
  assign n962 = ~n897 & n961;
  assign n963 = ~n896 & n962;
  assign n964 = ~n895 & n963;
  assign n965 = ~n894 & n964;
  assign n966 = ~n893 & n965;
  assign n967 = ~n892 & n966;
  assign n968 = ~n891 & n967;
  assign n969 = ~n890 & n968;
  assign n970 = ~n889 & n969;
  assign n971 = ~n888 & n970;
  assign n972 = ~n887 & n971;
  assign n973 = ~n886 & n972;
  assign n974 = ~n885 & n973;
  assign n975 = ~n884 & n974;
  assign n976 = ~n883 & n975;
  assign n977 = ~n882 & n976;
  assign n978 = ~n881 & n977;
  assign n979 = ~n880 & n978;
  assign n980 = ~n879 & n979;
  assign n981 = ~n877 & n980;
  assign n982 = ~n875 & n981;
  assign n983 = ~n869 & n982;
  assign n984 = ~n868 & n983;
  assign n985 = ~n867 & n984;
  assign n986 = ~n866 & n985;
  assign n987 = ~n859 & n986;
  assign n988 = ~n857 & n987;
  assign n989 = ~n855 & n988;
  assign n990 = ~n853 & n989;
  assign n991 = ~n850 & n990;
  assign n992 = ~n846 & n991;
  assign n993 = ~n839 & n992;
  assign n994 = ~n837 & n993;
  assign n995 = ~n829 & n994;
  assign n996 = ~n826 & n995;
  assign n997 = ~n817 & n996;
  assign n998 = ~n808 & n997;
  assign n999 = ~n807 & n998;
  assign n1000 = ~n806 & n999;
  assign n1001 = ~n805 & n1000;
  assign n1002 = ~n804 & n1001;
  assign n1003 = ~n803 & n1002;
  assign n1004 = ~n802 & n1003;
  assign n1005 = ~n801 & n1004;
  assign n1006 = ~n800 & n1005;
  assign n1007 = ~n799 & n1006;
  assign n1008 = ~n798 & n1007;
  assign n1009 = ~n797 & n1008;
  assign n1010 = ~n796 & n1009;
  assign n1011 = ~n795 & n1010;
  assign n1012 = ~n794 & n1011;
  assign n1013 = ~n793 & n1012;
  assign n1014 = ~n792 & n1013;
  assign n1015 = ~n791 & n1014;
  assign n1016 = ~n790 & n1015;
  assign n1017 = ~n789 & n1016;
  assign n1018 = ~n788 & n1017;
  assign n1019 = ~n787 & n1018;
  assign n1020 = ~n786 & n1019;
  assign n1021 = ~n784 & n1020;
  assign n1022 = ~n782 & n1021;
  assign n1023 = ~n773 & n1022;
  assign n1024 = ~n769 & n1023;
  assign n1025 = ~n760 & n1024;
  assign n1026 = ~n755 & n1025;
  assign n1027 = ~n746 & n1026;
  assign n1028 = ~n738 & n1027;
  assign n1029 = ~n736 & n1028;
  assign n1030 = ~n733 & n1029;
  assign n1031 = ~n725 & n1030;
  assign n1032 = ~n716 & n1031;
  assign n1033 = ~n715 & n1032;
  assign n1034 = ~n714 & n1033;
  assign n1035 = ~n713 & n1034;
  assign n1036 = ~n712 & n1035;
  assign n1037 = ~n704 & n1036;
  assign n1038 = ~n701 & n1037;
  assign n1039 = ~n692 & n1038;
  assign n1040 = ~n688 & n1039;
  assign h2 = n679 | ~n1040;
  assign n1042 = c & g0;
  assign n1043 = ~a & n1042;
  assign n1044 = b & n1043;
  assign n1045 = l & n1044;
  assign n1046 = ~m & n1045;
  assign n1047 = ~n & n1046;
  assign n1048 = v & n1047;
  assign n1049 = k0 & n1048;
  assign n1050 = ~a & ~j;
  assign n1051 = b & n1050;
  assign n1052 = l & n1051;
  assign n1053 = ~m & n1052;
  assign n1054 = ~n & n1053;
  assign n1055 = v & n1054;
  assign n1056 = k0 & n1055;
  assign n1057 = l & n103;
  assign n1058 = ~m & n1057;
  assign n1059 = ~n & n1058;
  assign n1060 = v & n1059;
  assign n1061 = a0 & n1060;
  assign n1062 = ~a & j;
  assign n1063 = b & n1062;
  assign n1064 = l & n1063;
  assign n1065 = ~m & n1064;
  assign n1066 = ~n & n1065;
  assign n1067 = a0 & n1066;
  assign n1068 = g0 & n118;
  assign n1069 = d & d0;
  assign n1070 = ~h & d0;
  assign n1071 = i & i0;
  assign n1072 = ~z & ~h0;
  assign n1073 = ~c0 & n1072;
  assign n1074 = ~b0 & n1073;
  assign n1075 = ~y & n1074;
  assign n1076 = ~n1071 & n1075;
  assign n1077 = ~n1070 & n1076;
  assign n1078 = ~n1069 & n1077;
  assign n1079 = ~n1068 & n1078;
  assign n1080 = ~n1067 & n1079;
  assign n1081 = ~n1061 & n1080;
  assign n1082 = ~n1056 & n1081;
  assign i2 = n1049 | ~n1082;
  assign n1084 = d & ~v;
  assign n1085 = w & n1084;
  assign n1086 = d0 & n1085;
  assign n1087 = a & g0;
  assign n1088 = ~j & n1087;
  assign n1089 = a & t;
  assign n1090 = i0 & n1089;
  assign n1091 = r & s;
  assign n1092 = l0 & n1091;
  assign n1093 = r & p0;
  assign n1094 = s & n1093;
  assign n1095 = m & ~v;
  assign n1096 = b0 & n1095;
  assign n1097 = c0 & n1095;
  assign n1098 = p0 & n1095;
  assign n1099 = d0 & n1095;
  assign n1100 = a & j0;
  assign n1101 = a & a0;
  assign n1102 = a & s0;
  assign n1103 = a & q0;
  assign n1104 = a & k0;
  assign n1105 = a & p0;
  assign n1106 = a & d0;
  assign n1107 = a & h0;
  assign n1108 = a & e0;
  assign n1109 = m & s0;
  assign n1110 = m & q0;
  assign n1111 = m & k0;
  assign n1112 = b & r0;
  assign n1113 = m & h0;
  assign n1114 = m & g0;
  assign n1115 = m & e0;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~n1113 & n1116;
  assign n1118 = ~n1112 & n1117;
  assign n1119 = ~n1111 & n1118;
  assign n1120 = ~n1110 & n1119;
  assign n1121 = ~n1109 & n1120;
  assign n1122 = ~n1108 & n1121;
  assign n1123 = ~n1107 & n1122;
  assign n1124 = ~n1106 & n1123;
  assign n1125 = ~n1105 & n1124;
  assign n1126 = ~n1104 & n1125;
  assign n1127 = ~n1103 & n1126;
  assign n1128 = ~n1102 & n1127;
  assign n1129 = ~n1101 & n1128;
  assign n1130 = ~n1100 & n1129;
  assign n1131 = ~n1099 & n1130;
  assign n1132 = ~n1098 & n1131;
  assign n1133 = ~n1097 & n1132;
  assign n1134 = ~n1096 & n1133;
  assign n1135 = ~n1094 & n1134;
  assign n1136 = ~n1092 & n1135;
  assign n1137 = ~n1090 & n1136;
  assign n1138 = ~n1088 & n1137;
  assign k1 = n1086 | ~n1138;
  assign n1140 = e & n1070;
  assign n1141 = ~a & n1140;
  assign n1142 = ~d & n1141;
  assign n1143 = ~g & n1142;
  assign n1144 = o & n1143;
  assign n1145 = p & n1144;
  assign n1146 = ~v & n1145;
  assign n1147 = ~h & u;
  assign n1148 = d0 & n1147;
  assign n1149 = ~a & n1148;
  assign n1150 = ~d & n1149;
  assign n1151 = ~g & n1150;
  assign n1152 = o & n1151;
  assign n1153 = p & n1152;
  assign n1154 = ~v & n1153;
  assign n1155 = d & n1141;
  assign n1156 = o & n1155;
  assign n1157 = ~p & n1156;
  assign n1158 = ~v & n1157;
  assign n1159 = d & n1149;
  assign n1160 = o & n1159;
  assign n1161 = ~p & n1160;
  assign n1162 = ~v & n1161;
  assign n1163 = e & ~h;
  assign n1164 = ~a & n1163;
  assign n1165 = o & n1164;
  assign n1166 = ~p & n1165;
  assign n1167 = ~v & n1166;
  assign n1168 = e0 & n1167;
  assign n1169 = ~a & n1147;
  assign n1170 = o & n1169;
  assign n1171 = ~p & n1170;
  assign n1172 = ~v & n1171;
  assign n1173 = e0 & n1172;
  assign n1174 = ~g & n1155;
  assign n1175 = ~v & n1174;
  assign n1176 = ~g & n1159;
  assign n1177 = ~v & n1176;
  assign n1178 = ~g & n1164;
  assign n1179 = ~v & n1178;
  assign n1180 = e0 & n1179;
  assign n1181 = ~g & n1169;
  assign n1182 = ~v & n1181;
  assign n1183 = e0 & n1182;
  assign n1184 = o & p;
  assign n1185 = q & n1184;
  assign n1186 = q0 & n1185;
  assign n1187 = p0 & n1185;
  assign n1188 = b & k;
  assign n1189 = a0 & n1188;
  assign n1190 = e & h;
  assign n1191 = e0 & n1190;
  assign n1192 = h & u;
  assign n1193 = e0 & n1192;
  assign n1194 = h & d0;
  assign n1195 = e & n1194;
  assign n1196 = d0 & n1192;
  assign n1197 = b & f0;
  assign n1198 = w & h0;
  assign n1199 = e & h0;
  assign n1200 = u & h0;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = ~n1198 & n1201;
  assign n1203 = ~n1197 & n1202;
  assign n1204 = ~n1196 & n1203;
  assign n1205 = ~n1195 & n1204;
  assign n1206 = ~n1193 & n1205;
  assign n1207 = ~n1191 & n1206;
  assign n1208 = ~n1189 & n1207;
  assign n1209 = ~n1187 & n1208;
  assign n1210 = ~n1186 & n1209;
  assign n1211 = ~n1183 & n1210;
  assign n1212 = ~n1180 & n1211;
  assign n1213 = ~n1177 & n1212;
  assign n1214 = ~n1175 & n1213;
  assign n1215 = ~n1173 & n1214;
  assign n1216 = ~n1168 & n1215;
  assign n1217 = ~n1162 & n1216;
  assign n1218 = ~n1158 & n1217;
  assign n1219 = ~n1154 & n1218;
  assign l1 = n1146 | ~n1219;
  assign n1221 = j & h0;
  assign n1222 = ~a & d;
  assign n1223 = ~e & n1222;
  assign n1224 = ~m & n1223;
  assign n1225 = o & n1224;
  assign n1226 = ~p & n1225;
  assign n1227 = ~u & n1226;
  assign n1228 = ~v & n1227;
  assign n1229 = ~w & n1228;
  assign n1230 = d0 & n1229;
  assign m1 = n1221 | n1230;
  assign n1232 = ~a & ~v;
  assign n1233 = c & n1232;
  assign n1234 = ~m & n1233;
  assign n1235 = ~e & n1234;
  assign n1236 = ~u & n1235;
  assign n1237 = ~w & n1236;
  assign n1238 = ~g & n1237;
  assign n1239 = d & n1238;
  assign n1240 = p0 & n1239;
  assign n1241 = ~a & ~m;
  assign n1242 = ~e & n1241;
  assign n1243 = o & n1242;
  assign n1244 = p & n1243;
  assign n1245 = ~u & n1244;
  assign n1246 = ~w & n1245;
  assign n1247 = ~g & n1246;
  assign n1248 = ~q & n1247;
  assign n1249 = q0 & n1248;
  assign n1250 = ~p & n1243;
  assign n1251 = ~u & n1250;
  assign n1252 = ~w & n1251;
  assign n1253 = e0 & n1252;
  assign n1254 = ~u & n1242;
  assign n1255 = ~w & n1254;
  assign n1256 = o0 & n1255;
  assign n1257 = w0 & n1256;
  assign n1258 = ~a & ~h;
  assign n1259 = ~m & n1258;
  assign n1260 = ~e & n1259;
  assign n1261 = ~u & n1260;
  assign n1262 = ~w & n1261;
  assign n1263 = s0 & n1262;
  assign n1264 = ~m & n1050;
  assign n1265 = ~e & n1264;
  assign n1266 = ~u & n1265;
  assign n1267 = ~w & n1266;
  assign n1268 = h0 & n1267;
  assign n1269 = g0 & n1062;
  assign n1270 = ~c & n1269;
  assign n1271 = ~h & n1270;
  assign n1272 = ~m & n1271;
  assign n1273 = ~a & f;
  assign n1274 = ~j & n1273;
  assign n1275 = v & n1274;
  assign n1276 = g0 & n1275;
  assign n1277 = ~n1272 & ~n1276;
  assign n1278 = ~n1268 & n1277;
  assign n1279 = ~n1263 & n1278;
  assign n1280 = ~n1257 & n1279;
  assign n1281 = ~n1253 & n1280;
  assign n1282 = ~n1249 & n1281;
  assign n1 = n1240 | ~n1282;
  assign n1284 = ~v & n179;
  assign n1285 = g & n1284;
  assign n1286 = q0 & n1285;
  assign n1287 = ~o & n1286;
  assign n1288 = p0 & n1284;
  assign n1289 = g & n1288;
  assign n1290 = ~o & n1289;
  assign n1291 = ~p & n1286;
  assign n1292 = ~p & n1289;
  assign n1293 = ~q & n1285;
  assign n1294 = q0 & n1293;
  assign n1295 = ~q & n1289;
  assign n1296 = i & n1258;
  assign n1297 = i0 & n1296;
  assign n1298 = ~n181 & ~n1297;
  assign n1299 = ~n1295 & n1298;
  assign n1300 = ~n1294 & n1299;
  assign n1301 = ~n1292 & n1300;
  assign n1302 = ~n1291 & n1301;
  assign n1303 = ~n1290 & n1302;
  assign o1 = n1287 | ~n1303;
  assign n1305 = r & n105;
  assign n1306 = ~s & n1305;
  assign n1307 = ~v & n1306;
  assign n1308 = ~k & n1307;
  assign n1309 = l & n1308;
  assign n1310 = a0 & n1309;
  assign n1311 = k0 & n1307;
  assign n1312 = a & ~h;
  assign n1313 = ~i & n1312;
  assign n1314 = i0 & n1313;
  assign n1315 = ~t & n1314;
  assign n1316 = ~i & n1258;
  assign n1317 = i0 & n1316;
  assign n1318 = ~a & j0;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~n1315 & n1319;
  assign n1321 = ~n1311 & n1320;
  assign r1 = n1310 | ~n1321;
  assign n1323 = v & n1264;
  assign n1324 = g0 & n1323;
  assign n1325 = ~f & n1324;
  assign n1326 = ~v & n1264;
  assign n1327 = k0 & n1326;
  assign n1328 = ~r & n1327;
  assign n1329 = n & n1264;
  assign n1330 = v & n1329;
  assign n1331 = k0 & n1330;
  assign n1332 = g0 & n1326;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1328 & n1333;
  assign v1 = n1325 | ~n1334;
  assign n1336 = k0 & n1091;
  assign n1337 = a0 & n1091;
  assign w1 = n1336 | n1337;
  assign n1339 = ~j & r0;
  assign n1340 = ~j & f0;
  assign n1341 = ~j & g0;
  assign n1342 = n1072 & ~n1341;
  assign n1343 = ~n1340 & n1342;
  assign x1 = n1339 | ~n1343;
  assign n1345 = j & ~z;
  assign n1346 = ~h0 & n1345;
  assign n1347 = ~f0 & n1072;
  assign n1348 = ~g0 & n1347;
  assign n1349 = ~r0 & n1348;
  assign y1 = n1346 | n1349;
  assign z1 = c0 | d0;
  assign c2 = h0;
  assign i1 = m0;
  assign j1 = n0;
  assign p1 = y;
  assign q1 = z;
  assign t1 = x0;
  assign u1 = y0;
endmodule


