// Benchmark "apex6" written by ABC on Tue May 16 16:07:44 2017

module apex6 ( 
    A, B, C, STW_N, QPR0, QPR1, QPR2, QPR3, QPR4, ENWIN, INZZZE, XZFR0,
    XZFR1, VZZZE, RXZ0, RXZ1, INFIN, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, XZ161, XZ162, XZ163, I2ZZZ0, I2ZZZ1,
    I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, XZ160_N, I2ZZZ7, TXMESS_N,
    PZZZE, RYZ, AXZ0, AXZ1, COMPPAR, MMERR, V1ZZZ0, PSRW, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3,
    I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, RPTEN, XZ320, XZ321, XZ322, XZ323,
    XZ324, CBT0, CBT1, CBT2, ESRSUM, SLAD0, SLAD1, SLAD2, SLAD3, XZFS,
    RPTWIN, PFIN, PSYNC, OFS1, OFS2, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3,
    P2ZZZ4, TXWRD0, P2ZZZ5, TXWRD1, P2ZZZ6, TXWRD2, P2ZZZ7, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, INYBB0, INYBB1, INYBB2, INYBB3,
    INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, VYBB0, VYBB1, TXWRD10, TXWRD11,
    TXWRD12, TXWRD13, TXWRD14, TXWRD15, PYBB0, PYBB1, PYBB2, PYBB3, PYBB4,
    PYBB5, PYBB6, PYBB7, PYBB8, ICLR, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3,
    P1ZZZ4, P1ZZZ5, P1ZZZ6, P1ZZZ7, VFIN,
    V2ZZZ2_P, QPR3_P, XZ323_P, P1ZZZ4_P, I1ZZZ3_P, TXWRD5_P, STW_F,
    TXWRD13_P, V1ZZZ4_P, P2ZZZ1_P, I2ZZZ2_P, TXWRD0_P, A_P, V2ZZZ1_P,
    TXWRD8_P, QPR4_P, XZ324_P, P1ZZZ3_P, I1ZZZ4_P, V1ZZZ3_P, COMPPAR_P,
    XZFS_P, P2ZZZ4_P, I2ZZZ3_P, XZ160_F, B_P, TXMESS_F, TXWRD7_P, P1ZZZ6_P,
    V2ZZZ4_P, I1ZZZ5_P, TXWRD15_P, V1ZZZ6_P, XZ161_P, RPTWIN_P, P2ZZZ3_P,
    AXZ0_P, I2ZZZ4_P, TXWRD2_P, C_P, P1ZZZ5_P, V2ZZZ3_P, I1ZZZ6_P, FSESR_P,
    V1ZZZ5_P, XZ162_P, TXWRD10_P, P1ZZZ0_P, OFS1_P, P2ZZZ6_P, AXZ1_P,
    I2ZZZ5_P, TXWRD1_P, I1ZZZ7_P, TXWRD9_P, ENWIN_P, V1ZZZ0_P, V2ZZZ6_P,
    XZ163_P, OFS2_P, P2ZZZ5_P, I1ZZZ0_P, I2ZZZ6_P, QPR0_P, XZ320_P,
    P1ZZZ7_P, TXWRD4_P, RXZ0_P, V2ZZZ5_P, SBUFF, V1ZZZ7_P, P2ZZZ0_P,
    TXWRD12_P, I2ZZZ7_P, P1ZZZ2_P, V2ZZZ0_P, I1ZZZ1_P, QPR1_P, XZ321_P,
    TXWRD3_P, RXZ1_P, V1ZZZ2_P, XZFR0_P, TD_P, I2ZZZ0_P, P2ZZZ7_P,
    TXWRD11_P, P1ZZZ1_P, I1ZZZ2_P, RYZ_P, QPR2_P, XZ322_P, V2ZZZ7_P,
    TXWRD6_P, V1ZZZ1_P, XZFR1_P, TXWRD14_P, P2ZZZ2_P, I2ZZZ1_P  );
  input  A, B, C, STW_N, QPR0, QPR1, QPR2, QPR3, QPR4, ENWIN, INZZZE,
    XZFR0, XZFR1, VZZZE, RXZ0, RXZ1, INFIN, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, XZ161, XZ162, XZ163, I2ZZZ0, I2ZZZ1,
    I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, XZ160_N, I2ZZZ7, TXMESS_N,
    PZZZE, RYZ, AXZ0, AXZ1, COMPPAR, MMERR, V1ZZZ0, PSRW, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3,
    I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, RPTEN, XZ320, XZ321, XZ322, XZ323,
    XZ324, CBT0, CBT1, CBT2, ESRSUM, SLAD0, SLAD1, SLAD2, SLAD3, XZFS,
    RPTWIN, PFIN, PSYNC, OFS1, OFS2, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3,
    P2ZZZ4, TXWRD0, P2ZZZ5, TXWRD1, P2ZZZ6, TXWRD2, P2ZZZ7, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, INYBB0, INYBB1, INYBB2, INYBB3,
    INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, VYBB0, VYBB1, TXWRD10, TXWRD11,
    TXWRD12, TXWRD13, TXWRD14, TXWRD15, PYBB0, PYBB1, PYBB2, PYBB3, PYBB4,
    PYBB5, PYBB6, PYBB7, PYBB8, ICLR, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3,
    P1ZZZ4, P1ZZZ5, P1ZZZ6, P1ZZZ7, VFIN;
  output V2ZZZ2_P, QPR3_P, XZ323_P, P1ZZZ4_P, I1ZZZ3_P, TXWRD5_P, STW_F,
    TXWRD13_P, V1ZZZ4_P, P2ZZZ1_P, I2ZZZ2_P, TXWRD0_P, A_P, V2ZZZ1_P,
    TXWRD8_P, QPR4_P, XZ324_P, P1ZZZ3_P, I1ZZZ4_P, V1ZZZ3_P, COMPPAR_P,
    XZFS_P, P2ZZZ4_P, I2ZZZ3_P, XZ160_F, B_P, TXMESS_F, TXWRD7_P, P1ZZZ6_P,
    V2ZZZ4_P, I1ZZZ5_P, TXWRD15_P, V1ZZZ6_P, XZ161_P, RPTWIN_P, P2ZZZ3_P,
    AXZ0_P, I2ZZZ4_P, TXWRD2_P, C_P, P1ZZZ5_P, V2ZZZ3_P, I1ZZZ6_P, FSESR_P,
    V1ZZZ5_P, XZ162_P, TXWRD10_P, P1ZZZ0_P, OFS1_P, P2ZZZ6_P, AXZ1_P,
    I2ZZZ5_P, TXWRD1_P, I1ZZZ7_P, TXWRD9_P, ENWIN_P, V1ZZZ0_P, V2ZZZ6_P,
    XZ163_P, OFS2_P, P2ZZZ5_P, I1ZZZ0_P, I2ZZZ6_P, QPR0_P, XZ320_P,
    P1ZZZ7_P, TXWRD4_P, RXZ0_P, V2ZZZ5_P, SBUFF, V1ZZZ7_P, P2ZZZ0_P,
    TXWRD12_P, I2ZZZ7_P, P1ZZZ2_P, V2ZZZ0_P, I1ZZZ1_P, QPR1_P, XZ321_P,
    TXWRD3_P, RXZ1_P, V1ZZZ2_P, XZFR0_P, TD_P, I2ZZZ0_P, P2ZZZ7_P,
    TXWRD11_P, P1ZZZ1_P, I1ZZZ2_P, RYZ_P, QPR2_P, XZ322_P, V2ZZZ7_P,
    TXWRD6_P, V1ZZZ1_P, XZFR1_P, TXWRD14_P, P2ZZZ2_P, I2ZZZ1_P;
  wire n235, n236, n237, n238, n239, n241, n242, n243, n244, n245, n247,
    n248, n249, n251, n252, n253, n254, n255, n256, n258, n259, n260, n261,
    n262, n263, n264, n266, n267, n268, n269, n270, n271, n273, n274, n276,
    n277, n278, n279, n280, n281, n283, n284, n285, n286, n287, n288, n289,
    n291, n292, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303,
    n304, n305, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n326, n327, n328, n329,
    n330, n331, n332, n333, n335, n336, n337, n338, n339, n340, n341, n342,
    n344, n345, n346, n347, n349, n350, n352, n353, n355, n356, n357, n358,
    n359, n360, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n380, n381, n383, n384, n385,
    n386, n387, n388, n389, n390, n392, n393, n394, n395, n396, n397, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n410, n411, n413,
    n414, n416, n417, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n477, n478, n479, n481, n482, n483, n485, n486, n488, n489, n491, n492,
    n493, n494, n495, n496, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n518,
    n519, n520, n521, n522, n523, n524, n525, n527, n528, n530, n531, n533,
    n534, n536, n537, n538, n539, n540, n541, n543, n544, n546, n547, n548,
    n549, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n602, n603, n605, n606, n607, n608, n610, n611, n613,
    n614, n615, n616, n617, n618, n619, n620, n622, n623, n624, n625, n627,
    n628, n630, n631, n633, n634, n637, n638, n640, n641, n643, n644, n645,
    n646, n647, n648, n649, n651, n652, n653, n654, n655, n656, n657, n658,
    n660, n661, n663, n664, n666, n667, n668, n669, n670, n672, n673, n675,
    n676, n677, n678, n679, n680, n681, n682, n684, n685, n687, n688, n689,
    n690, n691, n692, n693, n694, n696, n697, n698, n699, n701, n702, n704,
    n705, n707, n708, n709, n710, n711, n712, n713, n715, n716, n718, n719,
    n721, n722, n724, n725, n727, n728, n729, n730, n731, n732, n733, n734,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n752, n753, n756, n757, n759, n760, n762, n763, n764,
    n765, n766, n767, n768, n769, n771, n772, n774, n775, n777, n778, n780,
    n781, n783, n784, n786, n787, n788, n789, n790, n791, n792, n793, n795,
    n796, n797, n798, n799, n800, n802, n803, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n837, n838, n840, n841, n843, n844, n845, n846, n847, n848, n849,
    n850, n852, n853, n855, n856, n858, n859, n860, n862, n863, n865, n866,
    n867, n868, n869, n870, n871, n872, n874, n875, n877, n878, n879, n880,
    n881, n882, n883, n885, n886, n887, n888, n889, n890, n891, n892, n894,
    n895, n897, n898;
  assign n235 = VZZZE & VYBB0;
  assign n236 = ~RYZ & n235;
  assign n237 = ~RYZ & ~n236;
  assign n238 = V2ZZZ3 & n236;
  assign n239 = V2ZZZ2 & n237;
  assign V2ZZZ2_P = n238 | n239;
  assign n241 = ~QPR3 & ~RYZ;
  assign n242 = ~INFIN & ~PFIN;
  assign n243 = ~RYZ & n242;
  assign n244 = TXMESS_N & ~VFIN;
  assign n245 = n243 & n244;
  assign TXMESS_F = RYZ | n245;
  assign n247 = ~QPR0 & ~TXMESS_F;
  assign n248 = QPR0 & TXMESS_F;
  assign n249 = n243 & n248;
  assign QPR0_P = n247 | n249;
  assign n251 = QPR1 & TXMESS_F;
  assign n252 = n243 & n251;
  assign n253 = QPR1 & QPR0_P;
  assign n254 = ~QPR1 & ~TXMESS_F;
  assign n255 = ~QPR0_P & n254;
  assign n256 = ~n253 & ~n255;
  assign QPR1_P = n252 | ~n256;
  assign n258 = ~QPR1 & QPR2;
  assign n259 = QPR1 & ~QPR2;
  assign n260 = ~TXMESS_F & n259;
  assign n261 = ~QPR1_P & n260;
  assign n262 = ~RYZ & n258;
  assign n263 = QPR2 & QPR1_P;
  assign n264 = ~n262 & ~n263;
  assign QPR2_P = n261 | ~n264;
  assign n266 = ~QPR2 & ~RYZ;
  assign n267 = ~n241 & n266;
  assign n268 = ~n241 & QPR2_P;
  assign n269 = QPR2 & ~QPR2_P;
  assign n270 = n241 & n269;
  assign n271 = ~n268 & ~n270;
  assign QPR3_P = n267 | ~n271;
  assign n273 = ~PSYNC & ~ICLR;
  assign n274 = XZ320 & n273;
  assign XZ320_P = ~XZ320 & n273;
  assign n276 = XZ321 & ~XZ322;
  assign n277 = n274 & n276;
  assign n278 = ~XZ321 & XZ322;
  assign n279 = n273 & n278;
  assign n280 = XZ322 & XZ320_P;
  assign n281 = ~n279 & ~n280;
  assign XZ322_P = n277 | ~n281;
  assign n283 = XZ322 & ~XZ323;
  assign n284 = ~XZ322_P & n283;
  assign n285 = n273 & n284;
  assign n286 = XZ323 & XZ322_P;
  assign n287 = ~XZ322 & XZ323;
  assign n288 = n273 & n287;
  assign n289 = ~n286 & ~n288;
  assign XZ323_P = n285 | ~n289;
  assign n291 = PZZZE & PYBB0;
  assign n292 = ~RYZ & n291;
  assign n293 = ~RYZ & ~n292;
  assign n294 = PYBB0 & n293;
  assign n295 = ~RYZ & ~n294;
  assign n296 = PYBB5 & n294;
  assign n297 = P1ZZZ4 & n295;
  assign P1ZZZ4_P = n296 | n297;
  assign n299 = INZZZE & INYBB0;
  assign n300 = ~RYZ & n299;
  assign n301 = ~RYZ & ~n300;
  assign n302 = INYBB0 & n301;
  assign n303 = ~RYZ & ~n302;
  assign n304 = INYBB4 & n302;
  assign n305 = I1ZZZ3 & n303;
  assign I1ZZZ3_P = n304 | n305;
  assign n307 = ~B & ~C;
  assign n308 = ~TXMESS_N & ~VFIN;
  assign n309 = ~n307 & n308;
  assign n310 = n243 & n309;
  assign n311 = VFIN & n243;
  assign n312 = ~VFIN & n243;
  assign n313 = ~n309 & n312;
  assign n314 = ~INFIN & PFIN;
  assign n315 = ~RYZ & n314;
  assign n316 = INFIN & ~RYZ;
  assign n317 = TXWRD6 & n310;
  assign n318 = V1ZZZ5 & n311;
  assign n319 = TXWRD5 & n313;
  assign n320 = P1ZZZ5 & n315;
  assign n321 = I1ZZZ5 & n316;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n319 & n322;
  assign n324 = ~n318 & n323;
  assign TXWRD5_P = n317 | ~n324;
  assign n326 = A & ~VFIN;
  assign n327 = AXZ0 & n326;
  assign n328 = AXZ1 & n327;
  assign n329 = ~TXMESS_F & n328;
  assign n330 = n243 & n329;
  assign n331 = STW_N & ~VFIN;
  assign n332 = n243 & n331;
  assign n333 = ~RYZ & ~n332;
  assign STW_F = n330 | ~n333;
  assign n335 = TXWRD14 & n310;
  assign n336 = V2ZZZ5 & n311;
  assign n337 = TXWRD13 & n313;
  assign n338 = P2ZZZ5 & n315;
  assign n339 = I2ZZZ5 & n316;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~n337 & n340;
  assign n342 = ~n336 & n341;
  assign TXWRD13_P = n335 | ~n342;
  assign n344 = VYBB0 & n237;
  assign n345 = ~RYZ & ~n344;
  assign n346 = V1ZZZ5 & n344;
  assign n347 = V1ZZZ4 & n345;
  assign V1ZZZ4_P = n346 | n347;
  assign n349 = PYBB2 & n292;
  assign n350 = P2ZZZ1 & n293;
  assign P2ZZZ1_P = n349 | n350;
  assign n352 = INYBB3 & n300;
  assign n353 = I2ZZZ2 & n301;
  assign I2ZZZ2_P = n352 | n353;
  assign n355 = TXWRD1 & n310;
  assign n356 = V1ZZZ0 & n311;
  assign n357 = TXWRD0 & n313;
  assign n358 = P1ZZZ0 & n315;
  assign n359 = I1ZZZ0 & n316;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~n356 & n361;
  assign TXWRD0_P = n355 | ~n362;
  assign n364 = QPR0 & n258;
  assign n365 = ~A & CBT2;
  assign n366 = ~QPR3 & n365;
  assign n367 = ~QPR4 & n366;
  assign n368 = ~A & QPR3;
  assign n369 = QPR4 & n368;
  assign n370 = ~A & ~B;
  assign n371 = QPR3 & n370;
  assign n372 = ~A & ~n364;
  assign n373 = ~TXMESS_N & ~n372;
  assign n374 = ~n371 & n373;
  assign n375 = ~n369 & n374;
  assign n376 = ~n367 & n375;
  assign n377 = A & ~RYZ;
  assign n378 = ~RYZ & n376;
  assign A_P = n377 | n378;
  assign n380 = V2ZZZ2 & n236;
  assign n381 = V2ZZZ1 & n237;
  assign V2ZZZ1_P = n380 | n381;
  assign n383 = TXWRD9 & n310;
  assign n384 = V2ZZZ0 & n311;
  assign n385 = TXWRD8 & n313;
  assign n386 = P2ZZZ0 & n315;
  assign n387 = I2ZZZ0 & n316;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~n385 & n388;
  assign n390 = ~n384 & n389;
  assign TXWRD8_P = n383 | ~n390;
  assign n392 = QPR3 & ~QPR4;
  assign n393 = ~TXMESS_F & n392;
  assign n394 = ~QPR3_P & n393;
  assign n395 = QPR4 & n241;
  assign n396 = QPR4 & QPR3_P;
  assign n397 = ~n395 & ~n396;
  assign QPR4_P = n394 | ~n397;
  assign n399 = XZ321 & XZ322;
  assign n400 = XZ323 & n399;
  assign n401 = XZ324 & n400;
  assign n402 = XZ323 & ~XZ323_P;
  assign n403 = n273 & n402;
  assign n404 = ~n401 & n403;
  assign n405 = XZ324 & n273;
  assign n406 = ~n401 & n405;
  assign n407 = XZ323_P & n401;
  assign n408 = ~n406 & ~n407;
  assign XZ324_P = n404 | ~n408;
  assign n410 = PYBB4 & n294;
  assign n411 = P1ZZZ3 & n295;
  assign P1ZZZ3_P = n410 | n411;
  assign n413 = INYBB5 & n302;
  assign n414 = I1ZZZ4 & n303;
  assign I1ZZZ4_P = n413 | n414;
  assign n416 = V1ZZZ4 & n344;
  assign n417 = V1ZZZ3 & n345;
  assign V1ZZZ3_P = n416 | n417;
  assign n419 = ~QPR0 & SLAD3;
  assign n420 = QPR1 & n419;
  assign n421 = ~QPR2 & n420;
  assign n422 = QPR0 & SLAD2;
  assign n423 = QPR1 & n422;
  assign n424 = ~QPR2 & n423;
  assign n425 = SLAD1 & ~n364;
  assign n426 = n258 & n425;
  assign n427 = SLAD0 & n364;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n424 & n428;
  assign n430 = ~n421 & n429;
  assign n431 = ~QPR3 & ~QPR4;
  assign n432 = ~n430 & n431;
  assign n433 = n307 & n432;
  assign n434 = TXWRD0 & ~n307;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~TXMESS_N & ~RYZ;
  assign n437 = ~COMPPAR & n436;
  assign n438 = ~AXZ0 & n437;
  assign n439 = ~AXZ1 & n438;
  assign n440 = ~n435 & n439;
  assign n441 = ~TXMESS_N & ESRSUM;
  assign n442 = ~COMPPAR & n441;
  assign n443 = AXZ1 & n442;
  assign n444 = n377 & n443;
  assign n445 = ~TXMESS_N & ~MMERR;
  assign n446 = ~COMPPAR & n445;
  assign n447 = AXZ0 & n446;
  assign n448 = n377 & n447;
  assign n449 = ~RYZ & COMPPAR;
  assign n450 = ~AXZ0 & n449;
  assign n451 = ~AXZ1 & n450;
  assign n452 = n435 & n451;
  assign n453 = ~A & n437;
  assign n454 = ~n435 & n453;
  assign n455 = ~TXMESS_N & AXZ0;
  assign n456 = AXZ1 & n455;
  assign n457 = n377 & n456;
  assign n458 = COMPPAR & ~ESRSUM;
  assign n459 = AXZ1 & n458;
  assign n460 = n377 & n459;
  assign n461 = COMPPAR & MMERR;
  assign n462 = AXZ0 & n461;
  assign n463 = n377 & n462;
  assign n464 = ~A & n449;
  assign n465 = n435 & n464;
  assign n466 = TXMESS_N & ~RYZ;
  assign n467 = COMPPAR & n466;
  assign n468 = ~n465 & ~n467;
  assign n469 = ~n463 & n468;
  assign n470 = ~n460 & n469;
  assign n471 = ~n457 & n470;
  assign n472 = ~n454 & n471;
  assign n473 = ~n452 & n472;
  assign n474 = ~n448 & n473;
  assign n475 = ~n444 & n474;
  assign COMPPAR_P = n440 | ~n475;
  assign n477 = PSRW & ~OFS1;
  assign n478 = PSRW & ~OFS2;
  assign n479 = ~n477 & ~n478;
  assign OFS1_P = PSYNC & ~ICLR;
  assign n481 = XZFS & ~ICLR;
  assign n482 = ~n479 & n481;
  assign n483 = ~n479 & OFS1_P;
  assign XZFS_P = n482 | n483;
  assign n485 = PYBB5 & n292;
  assign n486 = P2ZZZ4 & n293;
  assign P2ZZZ4_P = n485 | n486;
  assign n488 = INYBB4 & n300;
  assign n489 = I2ZZZ3 & n301;
  assign I2ZZZ3_P = n488 | n489;
  assign n491 = ~XZ160_N & n401;
  assign n492 = n274 & n491;
  assign n493 = XZ160_N & n273;
  assign n494 = ~n401 & n493;
  assign n495 = XZ160_N & XZ320_P;
  assign n496 = ~n494 & ~n495;
  assign XZ160_F = n492 | ~n496;
  assign n498 = ~TXMESS_N & n364;
  assign n499 = ~QPR4 & ~CBT2;
  assign n500 = ~QPR4 & CBT1;
  assign n501 = ~QPR4 & CBT0;
  assign n502 = ~QPR3 & n498;
  assign n503 = ~n501 & n502;
  assign n504 = ~n500 & n503;
  assign n505 = ~n499 & n504;
  assign n506 = n498 & ~n505;
  assign n507 = ~B & CBT2;
  assign n508 = n506 & n507;
  assign n509 = n241 & n508;
  assign n510 = B & ~CBT2;
  assign n511 = n241 & n510;
  assign n512 = B & ~RYZ;
  assign n513 = ~n506 & n512;
  assign n514 = QPR4 & n512;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n511 & n515;
  assign B_P = n509 | ~n516;
  assign n518 = TXWRD8 & n310;
  assign n519 = V1ZZZ7 & n311;
  assign n520 = TXWRD7 & n313;
  assign n521 = P1ZZZ7 & n315;
  assign n522 = I1ZZZ7 & n316;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n520 & n523;
  assign n525 = ~n519 & n524;
  assign TXWRD7_P = n518 | ~n525;
  assign n527 = PYBB7 & n294;
  assign n528 = P1ZZZ6 & n295;
  assign P1ZZZ6_P = n527 | n528;
  assign n530 = V2ZZZ5 & n236;
  assign n531 = V2ZZZ4 & n237;
  assign V2ZZZ4_P = n530 | n531;
  assign n533 = INYBB6 & n302;
  assign n534 = I1ZZZ5 & n303;
  assign I1ZZZ5_P = n533 | n534;
  assign n536 = V2ZZZ7 & n311;
  assign n537 = TXWRD15 & n313;
  assign n538 = P2ZZZ7 & n315;
  assign n539 = I2ZZZ7 & n316;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~n537 & n540;
  assign TXWRD15_P = n536 | ~n541;
  assign n543 = V1ZZZ7 & n344;
  assign n544 = V1ZZZ6 & n345;
  assign V1ZZZ6_P = n543 | n544;
  assign n546 = ~XZ160_N & XZ160_F;
  assign n547 = XZ161 & n273;
  assign n548 = ~n546 & n547;
  assign n549 = ~XZ161 & n546;
  assign XZ161_P = n548 | n549;
  assign n551 = ~SLAD0 & ~SLAD1;
  assign n552 = ~SLAD2 & ~SLAD3;
  assign n553 = XZFS & PSYNC;
  assign n554 = n552 & n553;
  assign n555 = ENWIN & n401;
  assign n556 = ~XZ162 & n552;
  assign n557 = ~XZ163 & n556;
  assign n558 = SLAD2 & ~SLAD3;
  assign n559 = XZ162 & n558;
  assign n560 = ~XZ163 & n559;
  assign n561 = SLAD2 & SLAD3;
  assign n562 = XZ162 & n561;
  assign n563 = XZ163 & n562;
  assign n564 = ~SLAD2 & SLAD3;
  assign n565 = ~XZ162 & n564;
  assign n566 = XZ163 & n565;
  assign n567 = ~n563 & ~n566;
  assign n568 = ~n560 & n567;
  assign n569 = ~n557 & n568;
  assign n570 = n555 & ~n569;
  assign n571 = SLAD0 & ~SLAD1;
  assign n572 = XZ320 & n571;
  assign n573 = ~XZ160_N & n572;
  assign n574 = ~XZ161 & n573;
  assign n575 = n570 & n574;
  assign n576 = SLAD0 & SLAD1;
  assign n577 = XZ320 & n576;
  assign n578 = ~XZ160_N & n577;
  assign n579 = XZ161 & n578;
  assign n580 = n570 & n579;
  assign n581 = ~SLAD0 & SLAD1;
  assign n582 = XZ320 & n581;
  assign n583 = XZ160_N & n582;
  assign n584 = XZ161 & n583;
  assign n585 = n570 & n584;
  assign n586 = XZ160_N & XZ320;
  assign n587 = ~XZ161 & n586;
  assign n588 = n551 & n587;
  assign n589 = n570 & n588;
  assign n590 = ~n585 & ~n589;
  assign n591 = ~n580 & n590;
  assign n592 = ~n575 & n591;
  assign n593 = ~RYZ & n554;
  assign n594 = n551 & n593;
  assign n595 = ~RYZ & RPTWIN;
  assign n596 = ~RXZ1 & n595;
  assign n597 = ~RXZ0 & n595;
  assign n598 = ~RYZ & ~n592;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n596 & n599;
  assign RPTWIN_P = n594 | ~n600;
  assign n602 = PYBB4 & n292;
  assign n603 = P2ZZZ3 & n293;
  assign P2ZZZ3_P = n602 | n603;
  assign n605 = ~RYZ & AXZ0;
  assign n606 = ~n376 & n605;
  assign n607 = ~RYZ & ~AXZ0;
  assign n608 = n376 & n607;
  assign AXZ0_P = n606 | n608;
  assign n610 = INYBB5 & n300;
  assign n611 = I2ZZZ4 & n301;
  assign I2ZZZ4_P = n610 | n611;
  assign n613 = TXWRD3 & n310;
  assign n614 = V1ZZZ2 & n311;
  assign n615 = TXWRD2 & n313;
  assign n616 = P1ZZZ2 & n315;
  assign n617 = I1ZZZ2 & n316;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n615 & n618;
  assign n620 = ~n614 & n619;
  assign TXWRD2_P = n613 | ~n620;
  assign n622 = C & ~RYZ;
  assign n623 = ~n505 & n622;
  assign n624 = ~C & ~RYZ;
  assign n625 = n505 & n624;
  assign C_P = n623 | n625;
  assign n627 = PYBB6 & n294;
  assign n628 = P1ZZZ5 & n295;
  assign P1ZZZ5_P = n627 | n628;
  assign n630 = V2ZZZ4 & n236;
  assign n631 = V2ZZZ3 & n237;
  assign V2ZZZ3_P = n630 | n631;
  assign n633 = INYBB7 & n302;
  assign n634 = I1ZZZ6 & n303;
  assign I1ZZZ6_P = n633 | n634;
  assign OFS2_P = OFS1 & ~ICLR;
  assign n637 = OFS2 & OFS2_P;
  assign n638 = XZFR1 & ~ICLR;
  assign FSESR_P = n637 | n638;
  assign n640 = V1ZZZ6 & n344;
  assign n641 = V1ZZZ5 & n345;
  assign V1ZZZ5_P = n640 | n641;
  assign n643 = XZ161 & ~XZ162;
  assign n644 = XZ160_F & n643;
  assign n645 = ~XZ161_P & n644;
  assign n646 = ~XZ161 & XZ162;
  assign n647 = n273 & n646;
  assign n648 = XZ162 & XZ161_P;
  assign n649 = ~n647 & ~n648;
  assign XZ162_P = n645 | ~n649;
  assign n651 = TXWRD11 & n310;
  assign n652 = V2ZZZ2 & n311;
  assign n653 = TXWRD10 & n313;
  assign n654 = P2ZZZ2 & n315;
  assign n655 = I2ZZZ2 & n316;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n653 & n656;
  assign n658 = ~n652 & n657;
  assign TXWRD10_P = n651 | ~n658;
  assign n660 = PYBB1 & n294;
  assign n661 = P1ZZZ0 & n295;
  assign P1ZZZ0_P = n660 | n661;
  assign n663 = PYBB7 & n292;
  assign n664 = P2ZZZ6 & n293;
  assign P2ZZZ6_P = n663 | n664;
  assign n666 = AXZ0 & n376;
  assign n667 = ~RYZ & AXZ1;
  assign n668 = ~n666 & n667;
  assign n669 = ~RYZ & ~AXZ1;
  assign n670 = n666 & n669;
  assign AXZ1_P = n668 | n670;
  assign n672 = INYBB6 & n300;
  assign n673 = I2ZZZ5 & n301;
  assign I2ZZZ5_P = n672 | n673;
  assign n675 = TXWRD2 & n310;
  assign n676 = V1ZZZ1 & n311;
  assign n677 = TXWRD1 & n313;
  assign n678 = P1ZZZ1 & n315;
  assign n679 = I1ZZZ1 & n316;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~n677 & n680;
  assign n682 = ~n676 & n681;
  assign TXWRD1_P = n675 | ~n682;
  assign n684 = INYBB8 & n302;
  assign n685 = I1ZZZ7 & n303;
  assign I1ZZZ7_P = n684 | n685;
  assign n687 = TXWRD10 & n310;
  assign n688 = V2ZZZ1 & n311;
  assign n689 = TXWRD9 & n313;
  assign n690 = P2ZZZ1 & n315;
  assign n691 = I2ZZZ1 & n316;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n689 & n692;
  assign n694 = ~n688 & n693;
  assign TXWRD9_P = n687 | ~n694;
  assign n696 = XZFS & OFS1_P;
  assign n697 = ~n479 & n696;
  assign n698 = ENWIN & ~ICLR;
  assign n699 = ~n479 & n698;
  assign ENWIN_P = n697 | n699;
  assign n701 = V1ZZZ1 & n344;
  assign n702 = V1ZZZ0 & n345;
  assign V1ZZZ0_P = n701 | n702;
  assign n704 = V2ZZZ7 & n236;
  assign n705 = V2ZZZ6 & n237;
  assign V2ZZZ6_P = n704 | n705;
  assign n707 = XZ162 & ~XZ163;
  assign n708 = XZ160_F & n707;
  assign n709 = ~XZ162_P & n708;
  assign n710 = ~XZ162 & XZ163;
  assign n711 = n273 & n710;
  assign n712 = XZ163 & XZ162_P;
  assign n713 = ~n711 & ~n712;
  assign XZ163_P = n709 | ~n713;
  assign n715 = PYBB6 & n292;
  assign n716 = P2ZZZ5 & n293;
  assign P2ZZZ5_P = n715 | n716;
  assign n718 = INYBB1 & n302;
  assign n719 = I1ZZZ0 & n303;
  assign I1ZZZ0_P = n718 | n719;
  assign n721 = INYBB7 & n300;
  assign n722 = I2ZZZ6 & n301;
  assign I2ZZZ6_P = n721 | n722;
  assign n724 = PYBB8 & n294;
  assign n725 = P1ZZZ7 & n295;
  assign P1ZZZ7_P = n724 | n725;
  assign n727 = TXWRD5 & n310;
  assign n728 = V1ZZZ4 & n311;
  assign n729 = TXWRD4 & n313;
  assign n730 = P1ZZZ4 & n315;
  assign n731 = I1ZZZ4 & n316;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n729 & n732;
  assign n734 = ~n728 & n733;
  assign TXWRD4_P = n727 | ~n734;
  assign n736 = XZFS & n551;
  assign n737 = n552 & n736;
  assign n738 = ~ICLR & ~n554;
  assign n739 = n592 & n738;
  assign n740 = ~ICLR & n592;
  assign n741 = ~n737 & n740;
  assign n742 = ~n739 & ~n741;
  assign n743 = OFS1_P & n737;
  assign n744 = ~ICLR & ~n592;
  assign n745 = RPTWIN & ~ICLR;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~n743 & n746;
  assign n748 = RXZ0 & ~RPTWIN;
  assign n749 = ~n742 & n748;
  assign n750 = ~RXZ0 & ~n747;
  assign RXZ0_P = n749 | n750;
  assign n752 = V2ZZZ6 & n236;
  assign n753 = V2ZZZ5 & n237;
  assign V2ZZZ5_P = n752 | n753;
  assign SBUFF = ~TXMESS_N | RPTWIN;
  assign n756 = VYBB1 & n344;
  assign n757 = V1ZZZ7 & n345;
  assign V1ZZZ7_P = n756 | n757;
  assign n759 = PYBB1 & n292;
  assign n760 = P2ZZZ0 & n293;
  assign P2ZZZ0_P = n759 | n760;
  assign n762 = TXWRD13 & n310;
  assign n763 = V2ZZZ4 & n311;
  assign n764 = TXWRD12 & n313;
  assign n765 = P2ZZZ4 & n315;
  assign n766 = I2ZZZ4 & n316;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n764 & n767;
  assign n769 = ~n763 & n768;
  assign TXWRD12_P = n762 | ~n769;
  assign n771 = INYBB8 & n300;
  assign n772 = I2ZZZ7 & n301;
  assign I2ZZZ7_P = n771 | n772;
  assign n774 = PYBB3 & n294;
  assign n775 = P1ZZZ2 & n295;
  assign P1ZZZ2_P = n774 | n775;
  assign n777 = V2ZZZ1 & n236;
  assign n778 = V2ZZZ0 & n237;
  assign V2ZZZ0_P = n777 | n778;
  assign n780 = INYBB2 & n302;
  assign n781 = I1ZZZ1 & n303;
  assign I1ZZZ1_P = n780 | n781;
  assign n783 = ~XZ321 & n274;
  assign n784 = XZ321 & XZ320_P;
  assign XZ321_P = n783 | n784;
  assign n786 = TXWRD4 & n310;
  assign n787 = V1ZZZ3 & n311;
  assign n788 = TXWRD3 & n313;
  assign n789 = P1ZZZ3 & n315;
  assign n790 = I1ZZZ3 & n316;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n788 & n791;
  assign n793 = ~n787 & n792;
  assign TXWRD3_P = n786 | ~n793;
  assign n795 = RXZ1 & n747;
  assign n796 = ~n742 & n795;
  assign n797 = RXZ1 & RXZ0_P;
  assign n798 = ~RXZ1 & ~RXZ0_P;
  assign n799 = ~n747 & n798;
  assign n800 = ~n797 & ~n799;
  assign RXZ1_P = n796 | ~n800;
  assign n802 = V1ZZZ3 & n344;
  assign n803 = V1ZZZ2 & n345;
  assign V1ZZZ2_P = n802 | n803;
  assign n805 = ~XZ161 & XZ160_N;
  assign n806 = ~XZ162 & n805;
  assign n807 = ~XZ163 & n806;
  assign n808 = n401 & n807;
  assign n809 = ~XZFR0 & n808;
  assign n810 = n274 & n809;
  assign n811 = XZFR0 & XZ320_P;
  assign n812 = XZFR0 & ~n808;
  assign n813 = n273 & n812;
  assign n814 = ~n811 & ~n813;
  assign XZFR0_P = n810 | ~n814;
  assign n816 = RPTEN & ~ESRSUM;
  assign n817 = ~RYZ & n816;
  assign n818 = RPTWIN & n817;
  assign n819 = RXZ0 & n818;
  assign n820 = ~RXZ1 & n819;
  assign n821 = RPTEN & ESRSUM;
  assign n822 = ~RYZ & n821;
  assign n823 = RPTWIN & n822;
  assign n824 = ~RXZ0 & n823;
  assign n825 = RXZ1 & n824;
  assign n826 = ~QPR4 & ~SBUFF;
  assign n827 = ~n430 & n826;
  assign n828 = n241 & n827;
  assign n829 = ~RPTWIN & n449;
  assign n830 = ~COMPPAR_P & n829;
  assign n831 = ~COMPPAR & ~RPTWIN;
  assign n832 = COMPPAR_P & n831;
  assign n833 = ~n830 & ~n832;
  assign n834 = ~n828 & n833;
  assign n835 = ~n825 & n834;
  assign TD_P = n820 | ~n835;
  assign n837 = INYBB1 & n300;
  assign n838 = I2ZZZ0 & n301;
  assign I2ZZZ0_P = n837 | n838;
  assign n840 = PYBB8 & n292;
  assign n841 = P2ZZZ7 & n293;
  assign P2ZZZ7_P = n840 | n841;
  assign n843 = TXWRD12 & n310;
  assign n844 = V2ZZZ3 & n311;
  assign n845 = TXWRD11 & n313;
  assign n846 = P2ZZZ3 & n315;
  assign n847 = I2ZZZ3 & n316;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n845 & n848;
  assign n850 = ~n844 & n849;
  assign TXWRD11_P = n843 | ~n850;
  assign n852 = PYBB2 & n294;
  assign n853 = P1ZZZ1 & n295;
  assign P1ZZZ1_P = n852 | n853;
  assign n855 = INYBB3 & n302;
  assign n856 = I1ZZZ2 & n303;
  assign I1ZZZ2_P = n855 | n856;
  assign n858 = A & ~TXMESS_N;
  assign n859 = AXZ0 & n858;
  assign n860 = AXZ1 & n859;
  assign RYZ_P = ICLR | n860;
  assign n862 = VYBB1 & n236;
  assign n863 = V2ZZZ7 & n237;
  assign V2ZZZ7_P = n862 | n863;
  assign n865 = TXWRD7 & n310;
  assign n866 = V1ZZZ6 & n311;
  assign n867 = TXWRD6 & n313;
  assign n868 = P1ZZZ6 & n315;
  assign n869 = I1ZZZ6 & n316;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n867 & n870;
  assign n872 = ~n866 & n871;
  assign TXWRD6_P = n865 | ~n872;
  assign n874 = V1ZZZ2 & n344;
  assign n875 = V1ZZZ1 & n345;
  assign V1ZZZ1_P = n874 | n875;
  assign n877 = XZFR0 & ~XZFR1;
  assign n878 = ~XZFR0_P & n877;
  assign n879 = n273 & n878;
  assign n880 = XZFR1 & XZFR0_P;
  assign n881 = ~XZFR0 & XZFR1;
  assign n882 = n273 & n881;
  assign n883 = ~n880 & ~n882;
  assign XZFR1_P = n879 | ~n883;
  assign n885 = TXWRD15 & n310;
  assign n886 = V2ZZZ6 & n311;
  assign n887 = TXWRD14 & n313;
  assign n888 = P2ZZZ6 & n315;
  assign n889 = I2ZZZ6 & n316;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~n887 & n890;
  assign n892 = ~n886 & n891;
  assign TXWRD14_P = n885 | ~n892;
  assign n894 = PYBB3 & n292;
  assign n895 = P2ZZZ2 & n293;
  assign P2ZZZ2_P = n894 | n895;
  assign n897 = INYBB2 & n300;
  assign n898 = I2ZZZ1 & n301;
  assign I2ZZZ1_P = n897 | n898;
endmodule


