// Benchmark "rca_128" written by ABC on Sat Apr 23 20:18:06 2016

module rca_128 ( 
    a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7, a8, b8,
    a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15, b15,
    a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22, b22,
    a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29, b29,
    a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36, b36,
    a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43, b43,
    a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50, b50,
    a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57, b57,
    a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64, b64,
    a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71, b71,
    a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78, b78,
    a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85, b85,
    a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92, b92,
    a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99, b99,
    a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105, b105,
    a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111, b111,
    a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117, b117,
    a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123, b123,
    a124, b124, a125, b125, a126, b126, a127, b127,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128  );
  input  a0, b0, a1, b1, a2, b2, a3, b3, a4, b4, a5, b5, a6, b6, a7, b7,
    a8, b8, a9, b9, a10, b10, a11, b11, a12, b12, a13, b13, a14, b14, a15,
    b15, a16, b16, a17, b17, a18, b18, a19, b19, a20, b20, a21, b21, a22,
    b22, a23, b23, a24, b24, a25, b25, a26, b26, a27, b27, a28, b28, a29,
    b29, a30, b30, a31, b31, a32, b32, a33, b33, a34, b34, a35, b35, a36,
    b36, a37, b37, a38, b38, a39, b39, a40, b40, a41, b41, a42, b42, a43,
    b43, a44, b44, a45, b45, a46, b46, a47, b47, a48, b48, a49, b49, a50,
    b50, a51, b51, a52, b52, a53, b53, a54, b54, a55, b55, a56, b56, a57,
    b57, a58, b58, a59, b59, a60, b60, a61, b61, a62, b62, a63, b63, a64,
    b64, a65, b65, a66, b66, a67, b67, a68, b68, a69, b69, a70, b70, a71,
    b71, a72, b72, a73, b73, a74, b74, a75, b75, a76, b76, a77, b77, a78,
    b78, a79, b79, a80, b80, a81, b81, a82, b82, a83, b83, a84, b84, a85,
    b85, a86, b86, a87, b87, a88, b88, a89, b89, a90, b90, a91, b91, a92,
    b92, a93, b93, a94, b94, a95, b95, a96, b96, a97, b97, a98, b98, a99,
    b99, a100, b100, a101, b101, a102, b102, a103, b103, a104, b104, a105,
    b105, a106, b106, a107, b107, a108, b108, a109, b109, a110, b110, a111,
    b111, a112, b112, a113, b113, a114, b114, a115, b115, a116, b116, a117,
    b117, a118, b118, a119, b119, a120, b120, a121, b121, a122, b122, a123,
    b123, a124, b124, a125, b125, a126, b126, a127, b127;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29,
    s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43,
    s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57,
    s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71,
    s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85,
    s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99,
    s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111,
    s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123,
    s124, s125, s126, s127, s128;
  wire n386, n387, n389, n390, n391, n392, n393, n395, n396, n397, n398,
    n399, n400, n402, n403, n404, n405, n406, n407, n409, n410, n411, n412,
    n413, n414, n416, n417, n418, n419, n420, n421, n423, n424, n425, n426,
    n427, n428, n430, n431, n432, n433, n434, n435, n437, n438, n439, n440,
    n441, n442, n444, n445, n446, n447, n448, n449, n451, n452, n453, n454,
    n455, n456, n458, n459, n460, n461, n462, n463, n465, n466, n467, n468,
    n469, n470, n472, n473, n474, n475, n476, n477, n479, n480, n481, n482,
    n483, n484, n486, n487, n488, n489, n490, n491, n493, n494, n495, n496,
    n497, n498, n500, n501, n502, n503, n504, n505, n507, n508, n509, n510,
    n511, n512, n514, n515, n516, n517, n518, n519, n521, n522, n523, n524,
    n525, n526, n528, n529, n530, n531, n532, n533, n535, n536, n537, n538,
    n539, n540, n542, n543, n544, n545, n546, n547, n549, n550, n551, n552,
    n553, n554, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566,
    n567, n568, n570, n571, n572, n573, n574, n575, n577, n578, n579, n580,
    n581, n582, n584, n585, n586, n587, n588, n589, n591, n592, n593, n594,
    n595, n596, n598, n599, n600, n601, n602, n603, n605, n606, n607, n608,
    n609, n610, n612, n613, n614, n615, n616, n617, n619, n620, n621, n622,
    n623, n624, n626, n627, n628, n629, n630, n631, n633, n634, n635, n636,
    n637, n638, n640, n641, n642, n643, n644, n645, n647, n648, n649, n650,
    n651, n652, n654, n655, n656, n657, n658, n659, n661, n662, n663, n664,
    n665, n666, n668, n669, n670, n671, n672, n673, n675, n676, n677, n678,
    n679, n680, n682, n683, n684, n685, n686, n687, n689, n690, n691, n692,
    n693, n694, n696, n697, n698, n699, n700, n701, n703, n704, n705, n706,
    n707, n708, n710, n711, n712, n713, n714, n715, n717, n718, n719, n720,
    n721, n722, n724, n725, n726, n727, n728, n729, n731, n732, n733, n734,
    n735, n736, n738, n739, n740, n741, n742, n743, n745, n746, n747, n748,
    n749, n750, n752, n753, n754, n755, n756, n757, n759, n760, n761, n762,
    n763, n764, n766, n767, n768, n769, n770, n771, n773, n774, n775, n776,
    n777, n778, n780, n781, n782, n783, n784, n785, n787, n788, n789, n790,
    n791, n792, n794, n795, n796, n797, n798, n799, n801, n802, n803, n804,
    n805, n806, n808, n809, n810, n811, n812, n813, n815, n816, n817, n818,
    n819, n820, n822, n823, n824, n825, n826, n827, n829, n830, n831, n832,
    n833, n834, n836, n837, n838, n839, n840, n841, n843, n844, n845, n846,
    n847, n848, n850, n851, n852, n853, n854, n855, n857, n858, n859, n860,
    n861, n862, n864, n865, n866, n867, n868, n869, n871, n872, n873, n874,
    n875, n876, n878, n879, n880, n881, n882, n883, n885, n886, n887, n888,
    n889, n890, n892, n893, n894, n895, n896, n897, n899, n900, n901, n902,
    n903, n904, n906, n907, n908, n909, n910, n911, n913, n914, n915, n916,
    n917, n918, n920, n921, n922, n923, n924, n925, n927, n928, n929, n930,
    n931, n932, n934, n935, n936, n937, n938, n939, n941, n942, n943, n944,
    n945, n946, n948, n949, n950, n951, n952, n953, n955, n956, n957, n958,
    n959, n960, n962, n963, n964, n965, n966, n967, n969, n970, n971, n972,
    n973, n974, n976, n977, n978, n979, n980, n981, n983, n984, n985, n986,
    n987, n988, n990, n991, n992, n993, n994, n995, n997, n998, n999,
    n1000, n1001, n1002, n1004, n1005, n1006, n1007, n1008, n1009, n1011,
    n1012, n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021, n1022,
    n1023, n1025, n1026, n1027, n1028, n1029, n1030, n1032, n1033, n1034,
    n1035, n1036, n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1046,
    n1047, n1048, n1049, n1050, n1051, n1053, n1054, n1055, n1056, n1057,
    n1058, n1060, n1061, n1062, n1063, n1064, n1065, n1067, n1068, n1069,
    n1070, n1071, n1072, n1074, n1075, n1076, n1077, n1078, n1079, n1081,
    n1082, n1083, n1084, n1085, n1086, n1088, n1089, n1090, n1091, n1092,
    n1093, n1095, n1096, n1097, n1098, n1099, n1100, n1102, n1103, n1104,
    n1105, n1106, n1107, n1109, n1110, n1111, n1112, n1113, n1114, n1116,
    n1117, n1118, n1119, n1120, n1121, n1123, n1124, n1125, n1126, n1127,
    n1128, n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139,
    n1140, n1141, n1142, n1144, n1145, n1146, n1147, n1148, n1149, n1151,
    n1152, n1153, n1154, n1155, n1156, n1158, n1159, n1160, n1161, n1162,
    n1163, n1165, n1166, n1167, n1168, n1169, n1170, n1172, n1173, n1174,
    n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1186,
    n1187, n1188, n1189, n1190, n1191, n1193, n1194, n1195, n1196, n1197,
    n1198, n1200, n1201, n1202, n1203, n1204, n1205, n1207, n1208, n1209,
    n1210, n1211, n1212, n1214, n1215, n1216, n1217, n1218, n1219, n1221,
    n1222, n1223, n1224, n1225, n1226, n1228, n1229, n1230, n1231, n1232,
    n1233, n1235, n1236, n1237, n1238, n1239, n1240, n1242, n1243, n1244,
    n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253, n1254, n1256,
    n1257, n1258, n1259, n1260, n1261, n1263, n1264, n1265, n1266, n1267,
    n1268, n1270, n1271, n1272, n1273, n1274, n1275;
  assign n386 = a0 & b0;
  assign n387 = ~a0 & ~b0;
  assign s0 = ~n386 & ~n387;
  assign n389 = a1 & b1;
  assign n390 = ~a1 & ~b1;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & n391;
  assign n393 = ~n386 & ~n391;
  assign s1 = ~n392 & ~n393;
  assign n395 = ~n389 & ~n392;
  assign n396 = a2 & b2;
  assign n397 = ~a2 & ~b2;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n395 & n398;
  assign n400 = n395 & ~n398;
  assign s2 = ~n399 & ~n400;
  assign n402 = ~n396 & ~n399;
  assign n403 = a3 & b3;
  assign n404 = ~a3 & ~b3;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n402 & n405;
  assign n407 = n402 & ~n405;
  assign s3 = ~n406 & ~n407;
  assign n409 = ~n403 & ~n406;
  assign n410 = a4 & b4;
  assign n411 = ~a4 & ~b4;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n409 & n412;
  assign n414 = n409 & ~n412;
  assign s4 = ~n413 & ~n414;
  assign n416 = ~n410 & ~n413;
  assign n417 = a5 & b5;
  assign n418 = ~a5 & ~b5;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~n416 & n419;
  assign n421 = n416 & ~n419;
  assign s5 = ~n420 & ~n421;
  assign n423 = ~n417 & ~n420;
  assign n424 = a6 & b6;
  assign n425 = ~a6 & ~b6;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n423 & n426;
  assign n428 = n423 & ~n426;
  assign s6 = ~n427 & ~n428;
  assign n430 = ~n424 & ~n427;
  assign n431 = a7 & b7;
  assign n432 = ~a7 & ~b7;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n430 & n433;
  assign n435 = n430 & ~n433;
  assign s7 = ~n434 & ~n435;
  assign n437 = ~n431 & ~n434;
  assign n438 = a8 & b8;
  assign n439 = ~a8 & ~b8;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n437 & n440;
  assign n442 = n437 & ~n440;
  assign s8 = ~n441 & ~n442;
  assign n444 = ~n438 & ~n441;
  assign n445 = a9 & b9;
  assign n446 = ~a9 & ~b9;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n444 & n447;
  assign n449 = n444 & ~n447;
  assign s9 = ~n448 & ~n449;
  assign n451 = ~n445 & ~n448;
  assign n452 = a10 & b10;
  assign n453 = ~a10 & ~b10;
  assign n454 = ~n452 & ~n453;
  assign n455 = ~n451 & n454;
  assign n456 = n451 & ~n454;
  assign s10 = ~n455 & ~n456;
  assign n458 = ~n452 & ~n455;
  assign n459 = a11 & b11;
  assign n460 = ~a11 & ~b11;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n458 & n461;
  assign n463 = n458 & ~n461;
  assign s11 = ~n462 & ~n463;
  assign n465 = ~n459 & ~n462;
  assign n466 = a12 & b12;
  assign n467 = ~a12 & ~b12;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n465 & n468;
  assign n470 = n465 & ~n468;
  assign s12 = ~n469 & ~n470;
  assign n472 = ~n466 & ~n469;
  assign n473 = a13 & b13;
  assign n474 = ~a13 & ~b13;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n472 & n475;
  assign n477 = n472 & ~n475;
  assign s13 = ~n476 & ~n477;
  assign n479 = ~n473 & ~n476;
  assign n480 = a14 & b14;
  assign n481 = ~a14 & ~b14;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n479 & n482;
  assign n484 = n479 & ~n482;
  assign s14 = ~n483 & ~n484;
  assign n486 = ~n480 & ~n483;
  assign n487 = a15 & b15;
  assign n488 = ~a15 & ~b15;
  assign n489 = ~n487 & ~n488;
  assign n490 = ~n486 & n489;
  assign n491 = n486 & ~n489;
  assign s15 = ~n490 & ~n491;
  assign n493 = ~n487 & ~n490;
  assign n494 = a16 & b16;
  assign n495 = ~a16 & ~b16;
  assign n496 = ~n494 & ~n495;
  assign n497 = ~n493 & n496;
  assign n498 = n493 & ~n496;
  assign s16 = ~n497 & ~n498;
  assign n500 = ~n494 & ~n497;
  assign n501 = a17 & b17;
  assign n502 = ~a17 & ~b17;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n500 & n503;
  assign n505 = n500 & ~n503;
  assign s17 = ~n504 & ~n505;
  assign n507 = ~n501 & ~n504;
  assign n508 = a18 & b18;
  assign n509 = ~a18 & ~b18;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n507 & n510;
  assign n512 = n507 & ~n510;
  assign s18 = ~n511 & ~n512;
  assign n514 = ~n508 & ~n511;
  assign n515 = a19 & b19;
  assign n516 = ~a19 & ~b19;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n514 & n517;
  assign n519 = n514 & ~n517;
  assign s19 = ~n518 & ~n519;
  assign n521 = ~n515 & ~n518;
  assign n522 = a20 & b20;
  assign n523 = ~a20 & ~b20;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n521 & n524;
  assign n526 = n521 & ~n524;
  assign s20 = ~n525 & ~n526;
  assign n528 = ~n522 & ~n525;
  assign n529 = a21 & b21;
  assign n530 = ~a21 & ~b21;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n528 & n531;
  assign n533 = n528 & ~n531;
  assign s21 = ~n532 & ~n533;
  assign n535 = ~n529 & ~n532;
  assign n536 = a22 & b22;
  assign n537 = ~a22 & ~b22;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n535 & n538;
  assign n540 = n535 & ~n538;
  assign s22 = ~n539 & ~n540;
  assign n542 = ~n536 & ~n539;
  assign n543 = a23 & b23;
  assign n544 = ~a23 & ~b23;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n542 & n545;
  assign n547 = n542 & ~n545;
  assign s23 = ~n546 & ~n547;
  assign n549 = ~n543 & ~n546;
  assign n550 = a24 & b24;
  assign n551 = ~a24 & ~b24;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n549 & n552;
  assign n554 = n549 & ~n552;
  assign s24 = ~n553 & ~n554;
  assign n556 = ~n550 & ~n553;
  assign n557 = a25 & b25;
  assign n558 = ~a25 & ~b25;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n556 & n559;
  assign n561 = n556 & ~n559;
  assign s25 = ~n560 & ~n561;
  assign n563 = ~n557 & ~n560;
  assign n564 = a26 & b26;
  assign n565 = ~a26 & ~b26;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n563 & n566;
  assign n568 = n563 & ~n566;
  assign s26 = ~n567 & ~n568;
  assign n570 = ~n564 & ~n567;
  assign n571 = a27 & b27;
  assign n572 = ~a27 & ~b27;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n570 & n573;
  assign n575 = n570 & ~n573;
  assign s27 = ~n574 & ~n575;
  assign n577 = ~n571 & ~n574;
  assign n578 = a28 & b28;
  assign n579 = ~a28 & ~b28;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n577 & n580;
  assign n582 = n577 & ~n580;
  assign s28 = ~n581 & ~n582;
  assign n584 = ~n578 & ~n581;
  assign n585 = a29 & b29;
  assign n586 = ~a29 & ~b29;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n584 & n587;
  assign n589 = n584 & ~n587;
  assign s29 = ~n588 & ~n589;
  assign n591 = ~n585 & ~n588;
  assign n592 = a30 & b30;
  assign n593 = ~a30 & ~b30;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n591 & n594;
  assign n596 = n591 & ~n594;
  assign s30 = ~n595 & ~n596;
  assign n598 = ~n592 & ~n595;
  assign n599 = a31 & b31;
  assign n600 = ~a31 & ~b31;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n598 & n601;
  assign n603 = n598 & ~n601;
  assign s31 = ~n602 & ~n603;
  assign n605 = ~n599 & ~n602;
  assign n606 = a32 & b32;
  assign n607 = ~a32 & ~b32;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n605 & n608;
  assign n610 = n605 & ~n608;
  assign s32 = ~n609 & ~n610;
  assign n612 = ~n606 & ~n609;
  assign n613 = a33 & b33;
  assign n614 = ~a33 & ~b33;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n612 & n615;
  assign n617 = n612 & ~n615;
  assign s33 = ~n616 & ~n617;
  assign n619 = ~n613 & ~n616;
  assign n620 = a34 & b34;
  assign n621 = ~a34 & ~b34;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n619 & n622;
  assign n624 = n619 & ~n622;
  assign s34 = ~n623 & ~n624;
  assign n626 = ~n620 & ~n623;
  assign n627 = a35 & b35;
  assign n628 = ~a35 & ~b35;
  assign n629 = ~n627 & ~n628;
  assign n630 = ~n626 & n629;
  assign n631 = n626 & ~n629;
  assign s35 = ~n630 & ~n631;
  assign n633 = ~n627 & ~n630;
  assign n634 = a36 & b36;
  assign n635 = ~a36 & ~b36;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n633 & n636;
  assign n638 = n633 & ~n636;
  assign s36 = ~n637 & ~n638;
  assign n640 = ~n634 & ~n637;
  assign n641 = a37 & b37;
  assign n642 = ~a37 & ~b37;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n640 & n643;
  assign n645 = n640 & ~n643;
  assign s37 = ~n644 & ~n645;
  assign n647 = ~n641 & ~n644;
  assign n648 = a38 & b38;
  assign n649 = ~a38 & ~b38;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n647 & n650;
  assign n652 = n647 & ~n650;
  assign s38 = ~n651 & ~n652;
  assign n654 = ~n648 & ~n651;
  assign n655 = a39 & b39;
  assign n656 = ~a39 & ~b39;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n654 & n657;
  assign n659 = n654 & ~n657;
  assign s39 = ~n658 & ~n659;
  assign n661 = ~n655 & ~n658;
  assign n662 = a40 & b40;
  assign n663 = ~a40 & ~b40;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n661 & n664;
  assign n666 = n661 & ~n664;
  assign s40 = ~n665 & ~n666;
  assign n668 = ~n662 & ~n665;
  assign n669 = a41 & b41;
  assign n670 = ~a41 & ~b41;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n668 & n671;
  assign n673 = n668 & ~n671;
  assign s41 = ~n672 & ~n673;
  assign n675 = ~n669 & ~n672;
  assign n676 = a42 & b42;
  assign n677 = ~a42 & ~b42;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n675 & n678;
  assign n680 = n675 & ~n678;
  assign s42 = ~n679 & ~n680;
  assign n682 = ~n676 & ~n679;
  assign n683 = a43 & b43;
  assign n684 = ~a43 & ~b43;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n682 & n685;
  assign n687 = n682 & ~n685;
  assign s43 = ~n686 & ~n687;
  assign n689 = ~n683 & ~n686;
  assign n690 = a44 & b44;
  assign n691 = ~a44 & ~b44;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n689 & n692;
  assign n694 = n689 & ~n692;
  assign s44 = ~n693 & ~n694;
  assign n696 = ~n690 & ~n693;
  assign n697 = a45 & b45;
  assign n698 = ~a45 & ~b45;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n696 & n699;
  assign n701 = n696 & ~n699;
  assign s45 = ~n700 & ~n701;
  assign n703 = ~n697 & ~n700;
  assign n704 = a46 & b46;
  assign n705 = ~a46 & ~b46;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n703 & n706;
  assign n708 = n703 & ~n706;
  assign s46 = ~n707 & ~n708;
  assign n710 = ~n704 & ~n707;
  assign n711 = a47 & b47;
  assign n712 = ~a47 & ~b47;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n710 & n713;
  assign n715 = n710 & ~n713;
  assign s47 = ~n714 & ~n715;
  assign n717 = ~n711 & ~n714;
  assign n718 = a48 & b48;
  assign n719 = ~a48 & ~b48;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~n717 & n720;
  assign n722 = n717 & ~n720;
  assign s48 = ~n721 & ~n722;
  assign n724 = ~n718 & ~n721;
  assign n725 = a49 & b49;
  assign n726 = ~a49 & ~b49;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n724 & n727;
  assign n729 = n724 & ~n727;
  assign s49 = ~n728 & ~n729;
  assign n731 = ~n725 & ~n728;
  assign n732 = a50 & b50;
  assign n733 = ~a50 & ~b50;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n731 & n734;
  assign n736 = n731 & ~n734;
  assign s50 = ~n735 & ~n736;
  assign n738 = ~n732 & ~n735;
  assign n739 = a51 & b51;
  assign n740 = ~a51 & ~b51;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n738 & n741;
  assign n743 = n738 & ~n741;
  assign s51 = ~n742 & ~n743;
  assign n745 = ~n739 & ~n742;
  assign n746 = a52 & b52;
  assign n747 = ~a52 & ~b52;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n745 & n748;
  assign n750 = n745 & ~n748;
  assign s52 = ~n749 & ~n750;
  assign n752 = ~n746 & ~n749;
  assign n753 = a53 & b53;
  assign n754 = ~a53 & ~b53;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n752 & n755;
  assign n757 = n752 & ~n755;
  assign s53 = ~n756 & ~n757;
  assign n759 = ~n753 & ~n756;
  assign n760 = a54 & b54;
  assign n761 = ~a54 & ~b54;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n759 & n762;
  assign n764 = n759 & ~n762;
  assign s54 = ~n763 & ~n764;
  assign n766 = ~n760 & ~n763;
  assign n767 = a55 & b55;
  assign n768 = ~a55 & ~b55;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n766 & n769;
  assign n771 = n766 & ~n769;
  assign s55 = ~n770 & ~n771;
  assign n773 = ~n767 & ~n770;
  assign n774 = a56 & b56;
  assign n775 = ~a56 & ~b56;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n773 & n776;
  assign n778 = n773 & ~n776;
  assign s56 = ~n777 & ~n778;
  assign n780 = ~n774 & ~n777;
  assign n781 = a57 & b57;
  assign n782 = ~a57 & ~b57;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n780 & n783;
  assign n785 = n780 & ~n783;
  assign s57 = ~n784 & ~n785;
  assign n787 = ~n781 & ~n784;
  assign n788 = a58 & b58;
  assign n789 = ~a58 & ~b58;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n787 & n790;
  assign n792 = n787 & ~n790;
  assign s58 = ~n791 & ~n792;
  assign n794 = ~n788 & ~n791;
  assign n795 = a59 & b59;
  assign n796 = ~a59 & ~b59;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n794 & n797;
  assign n799 = n794 & ~n797;
  assign s59 = ~n798 & ~n799;
  assign n801 = ~n795 & ~n798;
  assign n802 = a60 & b60;
  assign n803 = ~a60 & ~b60;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n801 & n804;
  assign n806 = n801 & ~n804;
  assign s60 = ~n805 & ~n806;
  assign n808 = ~n802 & ~n805;
  assign n809 = a61 & b61;
  assign n810 = ~a61 & ~b61;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n808 & n811;
  assign n813 = n808 & ~n811;
  assign s61 = ~n812 & ~n813;
  assign n815 = ~n809 & ~n812;
  assign n816 = a62 & b62;
  assign n817 = ~a62 & ~b62;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n815 & n818;
  assign n820 = n815 & ~n818;
  assign s62 = ~n819 & ~n820;
  assign n822 = ~n816 & ~n819;
  assign n823 = a63 & b63;
  assign n824 = ~a63 & ~b63;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n822 & n825;
  assign n827 = n822 & ~n825;
  assign s63 = ~n826 & ~n827;
  assign n829 = ~n823 & ~n826;
  assign n830 = a64 & b64;
  assign n831 = ~a64 & ~b64;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n829 & n832;
  assign n834 = n829 & ~n832;
  assign s64 = ~n833 & ~n834;
  assign n836 = ~n830 & ~n833;
  assign n837 = a65 & b65;
  assign n838 = ~a65 & ~b65;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n836 & n839;
  assign n841 = n836 & ~n839;
  assign s65 = ~n840 & ~n841;
  assign n843 = ~n837 & ~n840;
  assign n844 = a66 & b66;
  assign n845 = ~a66 & ~b66;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~n843 & n846;
  assign n848 = n843 & ~n846;
  assign s66 = ~n847 & ~n848;
  assign n850 = ~n844 & ~n847;
  assign n851 = a67 & b67;
  assign n852 = ~a67 & ~b67;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n850 & n853;
  assign n855 = n850 & ~n853;
  assign s67 = ~n854 & ~n855;
  assign n857 = ~n851 & ~n854;
  assign n858 = a68 & b68;
  assign n859 = ~a68 & ~b68;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n857 & n860;
  assign n862 = n857 & ~n860;
  assign s68 = ~n861 & ~n862;
  assign n864 = ~n858 & ~n861;
  assign n865 = a69 & b69;
  assign n866 = ~a69 & ~b69;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n864 & n867;
  assign n869 = n864 & ~n867;
  assign s69 = ~n868 & ~n869;
  assign n871 = ~n865 & ~n868;
  assign n872 = a70 & b70;
  assign n873 = ~a70 & ~b70;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n871 & n874;
  assign n876 = n871 & ~n874;
  assign s70 = ~n875 & ~n876;
  assign n878 = ~n872 & ~n875;
  assign n879 = a71 & b71;
  assign n880 = ~a71 & ~b71;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n878 & n881;
  assign n883 = n878 & ~n881;
  assign s71 = ~n882 & ~n883;
  assign n885 = ~n879 & ~n882;
  assign n886 = a72 & b72;
  assign n887 = ~a72 & ~b72;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n885 & n888;
  assign n890 = n885 & ~n888;
  assign s72 = ~n889 & ~n890;
  assign n892 = ~n886 & ~n889;
  assign n893 = a73 & b73;
  assign n894 = ~a73 & ~b73;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n892 & n895;
  assign n897 = n892 & ~n895;
  assign s73 = ~n896 & ~n897;
  assign n899 = ~n893 & ~n896;
  assign n900 = a74 & b74;
  assign n901 = ~a74 & ~b74;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n899 & n902;
  assign n904 = n899 & ~n902;
  assign s74 = ~n903 & ~n904;
  assign n906 = ~n900 & ~n903;
  assign n907 = a75 & b75;
  assign n908 = ~a75 & ~b75;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n906 & n909;
  assign n911 = n906 & ~n909;
  assign s75 = ~n910 & ~n911;
  assign n913 = ~n907 & ~n910;
  assign n914 = a76 & b76;
  assign n915 = ~a76 & ~b76;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~n913 & n916;
  assign n918 = n913 & ~n916;
  assign s76 = ~n917 & ~n918;
  assign n920 = ~n914 & ~n917;
  assign n921 = a77 & b77;
  assign n922 = ~a77 & ~b77;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n920 & n923;
  assign n925 = n920 & ~n923;
  assign s77 = ~n924 & ~n925;
  assign n927 = ~n921 & ~n924;
  assign n928 = a78 & b78;
  assign n929 = ~a78 & ~b78;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n927 & n930;
  assign n932 = n927 & ~n930;
  assign s78 = ~n931 & ~n932;
  assign n934 = ~n928 & ~n931;
  assign n935 = a79 & b79;
  assign n936 = ~a79 & ~b79;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n934 & n937;
  assign n939 = n934 & ~n937;
  assign s79 = ~n938 & ~n939;
  assign n941 = ~n935 & ~n938;
  assign n942 = a80 & b80;
  assign n943 = ~a80 & ~b80;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n941 & n944;
  assign n946 = n941 & ~n944;
  assign s80 = ~n945 & ~n946;
  assign n948 = ~n942 & ~n945;
  assign n949 = a81 & b81;
  assign n950 = ~a81 & ~b81;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n948 & n951;
  assign n953 = n948 & ~n951;
  assign s81 = ~n952 & ~n953;
  assign n955 = ~n949 & ~n952;
  assign n956 = a82 & b82;
  assign n957 = ~a82 & ~b82;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~n955 & n958;
  assign n960 = n955 & ~n958;
  assign s82 = ~n959 & ~n960;
  assign n962 = ~n956 & ~n959;
  assign n963 = a83 & b83;
  assign n964 = ~a83 & ~b83;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n962 & n965;
  assign n967 = n962 & ~n965;
  assign s83 = ~n966 & ~n967;
  assign n969 = ~n963 & ~n966;
  assign n970 = a84 & b84;
  assign n971 = ~a84 & ~b84;
  assign n972 = ~n970 & ~n971;
  assign n973 = ~n969 & n972;
  assign n974 = n969 & ~n972;
  assign s84 = ~n973 & ~n974;
  assign n976 = ~n970 & ~n973;
  assign n977 = a85 & b85;
  assign n978 = ~a85 & ~b85;
  assign n979 = ~n977 & ~n978;
  assign n980 = ~n976 & n979;
  assign n981 = n976 & ~n979;
  assign s85 = ~n980 & ~n981;
  assign n983 = ~n977 & ~n980;
  assign n984 = a86 & b86;
  assign n985 = ~a86 & ~b86;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n983 & n986;
  assign n988 = n983 & ~n986;
  assign s86 = ~n987 & ~n988;
  assign n990 = ~n984 & ~n987;
  assign n991 = a87 & b87;
  assign n992 = ~a87 & ~b87;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n990 & n993;
  assign n995 = n990 & ~n993;
  assign s87 = ~n994 & ~n995;
  assign n997 = ~n991 & ~n994;
  assign n998 = a88 & b88;
  assign n999 = ~a88 & ~b88;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = ~n997 & n1000;
  assign n1002 = n997 & ~n1000;
  assign s88 = ~n1001 & ~n1002;
  assign n1004 = ~n998 & ~n1001;
  assign n1005 = a89 & b89;
  assign n1006 = ~a89 & ~b89;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1004 & n1007;
  assign n1009 = n1004 & ~n1007;
  assign s89 = ~n1008 & ~n1009;
  assign n1011 = ~n1005 & ~n1008;
  assign n1012 = a90 & b90;
  assign n1013 = ~a90 & ~b90;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = ~n1011 & n1014;
  assign n1016 = n1011 & ~n1014;
  assign s90 = ~n1015 & ~n1016;
  assign n1018 = ~n1012 & ~n1015;
  assign n1019 = a91 & b91;
  assign n1020 = ~a91 & ~b91;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = ~n1018 & n1021;
  assign n1023 = n1018 & ~n1021;
  assign s91 = ~n1022 & ~n1023;
  assign n1025 = ~n1019 & ~n1022;
  assign n1026 = a92 & b92;
  assign n1027 = ~a92 & ~b92;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1025 & n1028;
  assign n1030 = n1025 & ~n1028;
  assign s92 = ~n1029 & ~n1030;
  assign n1032 = ~n1026 & ~n1029;
  assign n1033 = a93 & b93;
  assign n1034 = ~a93 & ~b93;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = ~n1032 & n1035;
  assign n1037 = n1032 & ~n1035;
  assign s93 = ~n1036 & ~n1037;
  assign n1039 = ~n1033 & ~n1036;
  assign n1040 = a94 & b94;
  assign n1041 = ~a94 & ~b94;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n1039 & n1042;
  assign n1044 = n1039 & ~n1042;
  assign s94 = ~n1043 & ~n1044;
  assign n1046 = ~n1040 & ~n1043;
  assign n1047 = a95 & b95;
  assign n1048 = ~a95 & ~b95;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = ~n1046 & n1049;
  assign n1051 = n1046 & ~n1049;
  assign s95 = ~n1050 & ~n1051;
  assign n1053 = ~n1047 & ~n1050;
  assign n1054 = a96 & b96;
  assign n1055 = ~a96 & ~b96;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1053 & n1056;
  assign n1058 = n1053 & ~n1056;
  assign s96 = ~n1057 & ~n1058;
  assign n1060 = ~n1054 & ~n1057;
  assign n1061 = a97 & b97;
  assign n1062 = ~a97 & ~b97;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1060 & n1063;
  assign n1065 = n1060 & ~n1063;
  assign s97 = ~n1064 & ~n1065;
  assign n1067 = ~n1061 & ~n1064;
  assign n1068 = a98 & b98;
  assign n1069 = ~a98 & ~b98;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1067 & n1070;
  assign n1072 = n1067 & ~n1070;
  assign s98 = ~n1071 & ~n1072;
  assign n1074 = ~n1068 & ~n1071;
  assign n1075 = a99 & b99;
  assign n1076 = ~a99 & ~b99;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1074 & n1077;
  assign n1079 = n1074 & ~n1077;
  assign s99 = ~n1078 & ~n1079;
  assign n1081 = ~n1075 & ~n1078;
  assign n1082 = a100 & b100;
  assign n1083 = ~a100 & ~b100;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = ~n1081 & n1084;
  assign n1086 = n1081 & ~n1084;
  assign s100 = ~n1085 & ~n1086;
  assign n1088 = ~n1082 & ~n1085;
  assign n1089 = a101 & b101;
  assign n1090 = ~a101 & ~b101;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n1088 & n1091;
  assign n1093 = n1088 & ~n1091;
  assign s101 = ~n1092 & ~n1093;
  assign n1095 = ~n1089 & ~n1092;
  assign n1096 = a102 & b102;
  assign n1097 = ~a102 & ~b102;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1095 & n1098;
  assign n1100 = n1095 & ~n1098;
  assign s102 = ~n1099 & ~n1100;
  assign n1102 = ~n1096 & ~n1099;
  assign n1103 = a103 & b103;
  assign n1104 = ~a103 & ~b103;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~n1102 & n1105;
  assign n1107 = n1102 & ~n1105;
  assign s103 = ~n1106 & ~n1107;
  assign n1109 = ~n1103 & ~n1106;
  assign n1110 = a104 & b104;
  assign n1111 = ~a104 & ~b104;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n1109 & n1112;
  assign n1114 = n1109 & ~n1112;
  assign s104 = ~n1113 & ~n1114;
  assign n1116 = ~n1110 & ~n1113;
  assign n1117 = a105 & b105;
  assign n1118 = ~a105 & ~b105;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1116 & n1119;
  assign n1121 = n1116 & ~n1119;
  assign s105 = ~n1120 & ~n1121;
  assign n1123 = ~n1117 & ~n1120;
  assign n1124 = a106 & b106;
  assign n1125 = ~a106 & ~b106;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n1123 & n1126;
  assign n1128 = n1123 & ~n1126;
  assign s106 = ~n1127 & ~n1128;
  assign n1130 = ~n1124 & ~n1127;
  assign n1131 = a107 & b107;
  assign n1132 = ~a107 & ~b107;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1130 & n1133;
  assign n1135 = n1130 & ~n1133;
  assign s107 = ~n1134 & ~n1135;
  assign n1137 = ~n1131 & ~n1134;
  assign n1138 = a108 & b108;
  assign n1139 = ~a108 & ~b108;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1137 & n1140;
  assign n1142 = n1137 & ~n1140;
  assign s108 = ~n1141 & ~n1142;
  assign n1144 = ~n1138 & ~n1141;
  assign n1145 = a109 & b109;
  assign n1146 = ~a109 & ~b109;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = ~n1144 & n1147;
  assign n1149 = n1144 & ~n1147;
  assign s109 = ~n1148 & ~n1149;
  assign n1151 = ~n1145 & ~n1148;
  assign n1152 = a110 & b110;
  assign n1153 = ~a110 & ~b110;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = ~n1151 & n1154;
  assign n1156 = n1151 & ~n1154;
  assign s110 = ~n1155 & ~n1156;
  assign n1158 = ~n1152 & ~n1155;
  assign n1159 = a111 & b111;
  assign n1160 = ~a111 & ~b111;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = ~n1158 & n1161;
  assign n1163 = n1158 & ~n1161;
  assign s111 = ~n1162 & ~n1163;
  assign n1165 = ~n1159 & ~n1162;
  assign n1166 = a112 & b112;
  assign n1167 = ~a112 & ~b112;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n1165 & n1168;
  assign n1170 = n1165 & ~n1168;
  assign s112 = ~n1169 & ~n1170;
  assign n1172 = ~n1166 & ~n1169;
  assign n1173 = a113 & b113;
  assign n1174 = ~a113 & ~b113;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1172 & n1175;
  assign n1177 = n1172 & ~n1175;
  assign s113 = ~n1176 & ~n1177;
  assign n1179 = ~n1173 & ~n1176;
  assign n1180 = a114 & b114;
  assign n1181 = ~a114 & ~b114;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~n1179 & n1182;
  assign n1184 = n1179 & ~n1182;
  assign s114 = ~n1183 & ~n1184;
  assign n1186 = ~n1180 & ~n1183;
  assign n1187 = a115 & b115;
  assign n1188 = ~a115 & ~b115;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1186 & n1189;
  assign n1191 = n1186 & ~n1189;
  assign s115 = ~n1190 & ~n1191;
  assign n1193 = ~n1187 & ~n1190;
  assign n1194 = a116 & b116;
  assign n1195 = ~a116 & ~b116;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1193 & n1196;
  assign n1198 = n1193 & ~n1196;
  assign s116 = ~n1197 & ~n1198;
  assign n1200 = ~n1194 & ~n1197;
  assign n1201 = a117 & b117;
  assign n1202 = ~a117 & ~b117;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n1200 & n1203;
  assign n1205 = n1200 & ~n1203;
  assign s117 = ~n1204 & ~n1205;
  assign n1207 = ~n1201 & ~n1204;
  assign n1208 = a118 & b118;
  assign n1209 = ~a118 & ~b118;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~n1207 & n1210;
  assign n1212 = n1207 & ~n1210;
  assign s118 = ~n1211 & ~n1212;
  assign n1214 = ~n1208 & ~n1211;
  assign n1215 = a119 & b119;
  assign n1216 = ~a119 & ~b119;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~n1214 & n1217;
  assign n1219 = n1214 & ~n1217;
  assign s119 = ~n1218 & ~n1219;
  assign n1221 = ~n1215 & ~n1218;
  assign n1222 = a120 & b120;
  assign n1223 = ~a120 & ~b120;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n1221 & n1224;
  assign n1226 = n1221 & ~n1224;
  assign s120 = ~n1225 & ~n1226;
  assign n1228 = ~n1222 & ~n1225;
  assign n1229 = a121 & b121;
  assign n1230 = ~a121 & ~b121;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = ~n1228 & n1231;
  assign n1233 = n1228 & ~n1231;
  assign s121 = ~n1232 & ~n1233;
  assign n1235 = ~n1229 & ~n1232;
  assign n1236 = a122 & b122;
  assign n1237 = ~a122 & ~b122;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1235 & n1238;
  assign n1240 = n1235 & ~n1238;
  assign s122 = ~n1239 & ~n1240;
  assign n1242 = ~n1236 & ~n1239;
  assign n1243 = a123 & b123;
  assign n1244 = ~a123 & ~b123;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n1242 & n1245;
  assign n1247 = n1242 & ~n1245;
  assign s123 = ~n1246 & ~n1247;
  assign n1249 = ~n1243 & ~n1246;
  assign n1250 = a124 & b124;
  assign n1251 = ~a124 & ~b124;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1249 & n1252;
  assign n1254 = n1249 & ~n1252;
  assign s124 = ~n1253 & ~n1254;
  assign n1256 = ~n1250 & ~n1253;
  assign n1257 = a125 & b125;
  assign n1258 = ~a125 & ~b125;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1256 & n1259;
  assign n1261 = n1256 & ~n1259;
  assign s125 = ~n1260 & ~n1261;
  assign n1263 = ~n1257 & ~n1260;
  assign n1264 = a126 & b126;
  assign n1265 = ~a126 & ~b126;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1263 & n1266;
  assign n1268 = n1263 & ~n1266;
  assign s126 = ~n1267 & ~n1268;
  assign n1270 = ~n1264 & ~n1267;
  assign n1271 = a127 & b127;
  assign n1272 = ~a127 & ~b127;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~n1270 & n1273;
  assign n1275 = n1270 & ~n1273;
  assign s127 = ~n1274 & ~n1275;
  assign s128 = n1271 | n1274;
endmodule


