// Benchmark "i8" written by ABC on Tue May 16 16:07:50 2017

module i8 ( 
    \V47(24) , \V84(31) , \V15(14) , \V84(30) , \V47(21) , \V47(20) ,
    \V15(11) , \V15(10) , \V47(27) , \V47(26) , \V47(29) , \V47(28) ,
    \V47(31) , \V133(10) , \V47(30) , \V116(27) , \V116(26) , \V116(29) ,
    \V116(28) , \V116(3) , \V116(2) , \V116(5) , \V116(4) , \V116(21) ,
    \V116(1) , \V116(20) , \V116(0) , \V47(0) , \V116(23) , \V47(1) ,
    \V116(22) , \V47(2) , \V116(25) , \V121(17) , \V47(3) , \V116(24) ,
    \V121(16) , \V47(4) , \V116(17) , \V116(7) , \V47(5) , \V116(16) ,
    \V116(6) , \V47(6) , \V116(19) , \V48(0) , \V116(9) , \V47(7) ,
    \V116(18) , \V116(8) , \V47(8) , \V47(9) , \V118(1) , \V118(0) ,
    \V49(0) , \V116(11) , \V84(0) , \V116(10) , \V84(1) , \V116(13) ,
    \V84(2) , \V116(12) , \V84(3) , \V116(15) , \V84(4) , \V119(0) ,
    \V116(14) , \V84(5) , \V84(6) , \V84(7) , \V84(8) , \V84(9) ,
    \V84(13) , \V116(31) , \V84(12) , \V116(30) , \V84(15) , \V84(14) ,
    \V84(11) , \V84(10) , \V133(3) , \V133(2) , \V133(5) , \V15(0) ,
    \V133(4) , \V15(1) , \V84(17) , \V50(0) , \V15(2) , \V84(16) ,
    \V15(3) , \V133(1) , \V84(19) , \V15(4) , \V133(0) , \V84(18) ,
    \V15(5) , \V84(23) , \V15(6) , \V84(22) , \V15(7) , \V84(25) ,
    \V15(8) , \V51(0) , \V47(13) , \V84(24) , \V15(9) , \V47(12) ,
    \V133(7) , \V47(15) , \V133(6) , \V47(14) , \V133(9) , \V84(21) ,
    \V133(8) , \V84(20) , \V47(11) , \V52(0) , \V47(10) , \V84(27) ,
    \V84(26) , \V84(29) , \V47(17) , \V84(28) , \V122(0) , \V47(16) ,
    \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V15(13) , \V47(25) ,
    \V15(12) ,
    \V165(11) , \V165(10) , \V165(13) , \V165(12) , \V165(14) , \V197(31) ,
    \V197(30) , \V212(3) , \V212(2) , \V212(5) , \V212(4) , \V212(1) ,
    \V212(0) , \V212(7) , \V212(6) , \V213(0) , \V212(9) , \V212(8) ,
    \V150(0) , \V214(0) , \V165(3) , \V165(2) , \V165(5) , \V165(4) ,
    \V165(1) , \V165(0) , \V212(11) , \V212(10) , \V212(13) , \V165(7) ,
    \V212(12) , \V165(6) , \V165(9) , \V212(14) , \V165(8) , \V142(3) ,
    \V142(2) , \V142(5) , \V142(4) , \V142(1) , \V142(0) , \V143(0) ,
    \V197(27) , \V197(26) , \V197(29) , \V197(28) , \V145(1) , \V145(0) ,
    \V197(21) , \V197(20) , \V197(23) , \V197(22) , \V197(25) , \V197(24) ,
    \V146(0) , \V197(17) , \V197(16) , \V197(19) , \V197(18) , \V134(0) ,
    \V197(3) , \V197(11) , \V197(2) , \V197(10) , \V197(5) , \V197(13) ,
    \V149(2) , \V197(4) , \V197(12) , \V197(15) , \V197(14) , \V197(1) ,
    \V197(0) , \V149(1) , \V149(0) , \V136(1) , \V197(7) , \V136(0) ,
    \V197(6) , \V197(9) , \V197(8)   );
  input  \V47(24) , \V84(31) , \V15(14) , \V84(30) , \V47(21) ,
    \V47(20) , \V15(11) , \V15(10) , \V47(27) , \V47(26) , \V47(29) ,
    \V47(28) , \V47(31) , \V133(10) , \V47(30) , \V116(27) , \V116(26) ,
    \V116(29) , \V116(28) , \V116(3) , \V116(2) , \V116(5) , \V116(4) ,
    \V116(21) , \V116(1) , \V116(20) , \V116(0) , \V47(0) , \V116(23) ,
    \V47(1) , \V116(22) , \V47(2) , \V116(25) , \V121(17) , \V47(3) ,
    \V116(24) , \V121(16) , \V47(4) , \V116(17) , \V116(7) , \V47(5) ,
    \V116(16) , \V116(6) , \V47(6) , \V116(19) , \V48(0) , \V116(9) ,
    \V47(7) , \V116(18) , \V116(8) , \V47(8) , \V47(9) , \V118(1) ,
    \V118(0) , \V49(0) , \V116(11) , \V84(0) , \V116(10) , \V84(1) ,
    \V116(13) , \V84(2) , \V116(12) , \V84(3) , \V116(15) , \V84(4) ,
    \V119(0) , \V116(14) , \V84(5) , \V84(6) , \V84(7) , \V84(8) ,
    \V84(9) , \V84(13) , \V116(31) , \V84(12) , \V116(30) , \V84(15) ,
    \V84(14) , \V84(11) , \V84(10) , \V133(3) , \V133(2) , \V133(5) ,
    \V15(0) , \V133(4) , \V15(1) , \V84(17) , \V50(0) , \V15(2) ,
    \V84(16) , \V15(3) , \V133(1) , \V84(19) , \V15(4) , \V133(0) ,
    \V84(18) , \V15(5) , \V84(23) , \V15(6) , \V84(22) , \V15(7) ,
    \V84(25) , \V15(8) , \V51(0) , \V47(13) , \V84(24) , \V15(9) ,
    \V47(12) , \V133(7) , \V47(15) , \V133(6) , \V47(14) , \V133(9) ,
    \V84(21) , \V133(8) , \V84(20) , \V47(11) , \V52(0) , \V47(10) ,
    \V84(27) , \V84(26) , \V84(29) , \V47(17) , \V84(28) , \V122(0) ,
    \V47(16) , \V47(19) , \V47(18) , \V47(23) , \V47(22) , \V15(13) ,
    \V47(25) , \V15(12) ;
  output \V165(11) , \V165(10) , \V165(13) , \V165(12) , \V165(14) ,
    \V197(31) , \V197(30) , \V212(3) , \V212(2) , \V212(5) , \V212(4) ,
    \V212(1) , \V212(0) , \V212(7) , \V212(6) , \V213(0) , \V212(9) ,
    \V212(8) , \V150(0) , \V214(0) , \V165(3) , \V165(2) , \V165(5) ,
    \V165(4) , \V165(1) , \V165(0) , \V212(11) , \V212(10) , \V212(13) ,
    \V165(7) , \V212(12) , \V165(6) , \V165(9) , \V212(14) , \V165(8) ,
    \V142(3) , \V142(2) , \V142(5) , \V142(4) , \V142(1) , \V142(0) ,
    \V143(0) , \V197(27) , \V197(26) , \V197(29) , \V197(28) , \V145(1) ,
    \V145(0) , \V197(21) , \V197(20) , \V197(23) , \V197(22) , \V197(25) ,
    \V197(24) , \V146(0) , \V197(17) , \V197(16) , \V197(19) , \V197(18) ,
    \V134(0) , \V197(3) , \V197(11) , \V197(2) , \V197(10) , \V197(5) ,
    \V197(13) , \V149(2) , \V197(4) , \V197(12) , \V197(15) , \V197(14) ,
    \V197(1) , \V197(0) , \V149(1) , \V149(0) , \V136(1) , \V197(7) ,
    \V136(0) , \V197(6) , \V197(9) , \V197(8) ;
  wire n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n384, n385, n386, n388, n389, n390,
    n392, n393, n394, n396, n397, n398, n400, n401, n402, n404, n405, n406,
    n408, n409, n410, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n423, n424, n425, n427, n428, n429, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n466, n467, n468, n469, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n543, n544, n545, n547, n548, n549, n551, n552, n553,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n567,
    n568, n569, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n595, n596, n597, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n623, n624, n625, n626, n627, n628, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n640, n641, n642, n643, n644, n645, n647, n648,
    n649, n650, n651, n652, n654, n655, n656, n657, n658, n659, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n736, n737, n738, n739,
    n740, n741, n742, n743, n745, n746, n747, n748, n749, n750, n751, n752,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201;
  assign n215 = ~\V133(10)  & ~\V133(2) ;
  assign n216 = ~\V133(5)  & ~\V133(6) ;
  assign n217 = ~\V133(10)  & \V133(8) ;
  assign n218 = \V133(1)  & n216;
  assign n219 = n215 & n218;
  assign n220 = \V133(1)  & n217;
  assign n221 = ~\V133(0)  & \V133(7) ;
  assign n222 = ~\V133(5)  & ~\V133(0) ;
  assign n223 = ~n221 & ~n222;
  assign n224 = ~n220 & n223;
  assign n225 = ~n219 & n224;
  assign n226 = \V133(2)  & \V133(1) ;
  assign n227 = \V133(3)  & n226;
  assign n228 = ~\V133(10)  & ~n227;
  assign n229 = ~n225 & n228;
  assign n230 = ~\V133(10)  & \V133(9) ;
  assign n231 = ~\V133(10)  & ~\V133(7) ;
  assign n232 = ~\V133(9)  & n231;
  assign n233 = ~\V133(4)  & ~\V133(9) ;
  assign n234 = \V133(3)  & n233;
  assign n235 = ~\V133(6)  & n233;
  assign n236 = ~\V133(2)  & n235;
  assign n237 = ~n230 & ~n232;
  assign n238 = ~n234 & ~n236;
  assign n239 = ~n237 & n238;
  assign n240 = ~\V133(1)  & n233;
  assign n241 = n235 & n240;
  assign n242 = n239 & ~n241;
  assign n243 = n229 & ~n242;
  assign n244 = n225 & n228;
  assign n245 = \V133(2)  & n216;
  assign n246 = \V133(2)  & \V133(8) ;
  assign n247 = ~n226 & ~n246;
  assign n248 = ~n245 & n247;
  assign n249 = n244 & n248;
  assign n250 = ~n242 & n249;
  assign n251 = ~n228 & ~n242;
  assign n252 = n244 & ~n248;
  assign n253 = ~n242 & n252;
  assign n254 = ~\V133(10)  & ~\V133(9) ;
  assign n255 = n226 & n254;
  assign n256 = n228 & n232;
  assign n257 = n233 & n256;
  assign n258 = n255 & n257;
  assign n259 = ~\V133(7)  & n249;
  assign n260 = ~n216 & n259;
  assign n261 = ~n215 & n249;
  assign n262 = \V133(1)  & n249;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n260 & n263;
  assign n265 = ~n242 & ~n264;
  assign n266 = \V47(20)  & n243;
  assign n267 = \V47(13)  & n250;
  assign n268 = \V47(28)  & n251;
  assign n269 = \V47(17)  & n253;
  assign n270 = \V116(28)  & n230;
  assign n271 = \V84(28)  & n258;
  assign n272 = ~n265 & ~n271;
  assign n273 = ~n270 & n272;
  assign n274 = ~n269 & n273;
  assign n275 = ~n268 & n274;
  assign n276 = ~n267 & n275;
  assign \V165(11)  = n266 | ~n276;
  assign n278 = \V47(19)  & n243;
  assign n279 = \V47(12)  & n250;
  assign n280 = \V47(27)  & n251;
  assign n281 = \V47(16)  & n253;
  assign n282 = \V116(27)  & n230;
  assign n283 = \V84(27)  & n258;
  assign n284 = ~n265 & ~n283;
  assign n285 = ~n282 & n284;
  assign n286 = ~n281 & n285;
  assign n287 = ~n280 & n286;
  assign n288 = ~n279 & n287;
  assign \V165(10)  = n278 | ~n288;
  assign n290 = \V47(22)  & n243;
  assign n291 = \V47(15)  & n250;
  assign n292 = \V47(30)  & n251;
  assign n293 = \V47(19)  & n253;
  assign n294 = \V116(30)  & n230;
  assign n295 = \V84(30)  & n258;
  assign n296 = ~n265 & ~n295;
  assign n297 = ~n294 & n296;
  assign n298 = ~n293 & n297;
  assign n299 = ~n292 & n298;
  assign n300 = ~n291 & n299;
  assign \V165(13)  = n290 | ~n300;
  assign n302 = \V47(21)  & n243;
  assign n303 = \V47(14)  & n250;
  assign n304 = \V47(29)  & n251;
  assign n305 = \V47(18)  & n253;
  assign n306 = \V116(29)  & n230;
  assign n307 = \V84(29)  & n258;
  assign n308 = ~n265 & ~n307;
  assign n309 = ~n306 & n308;
  assign n310 = ~n305 & n309;
  assign n311 = ~n304 & n310;
  assign n312 = ~n303 & n311;
  assign \V165(12)  = n302 | ~n312;
  assign n314 = \V47(23)  & n243;
  assign n315 = \V47(16)  & n250;
  assign n316 = \V47(31)  & n251;
  assign n317 = \V47(20)  & n253;
  assign n318 = \V116(31)  & n230;
  assign n319 = \V84(31)  & n258;
  assign n320 = ~n265 & ~n319;
  assign n321 = ~n318 & n320;
  assign n322 = ~n317 & n321;
  assign n323 = ~n316 & n322;
  assign n324 = ~n315 & n323;
  assign \V165(14)  = n314 | ~n324;
  assign n326 = ~n236 & ~n241;
  assign n327 = \V133(7)  & ~\V133(9) ;
  assign n328 = ~\V133(1)  & n327;
  assign n329 = ~\V133(5)  & n241;
  assign n330 = \V133(5)  & ~\V133(1) ;
  assign n331 = ~\V133(9)  & n330;
  assign n332 = ~\V118(0)  & n331;
  assign n333 = ~\V133(1)  & ~\V133(0) ;
  assign n334 = \V133(5)  & n333;
  assign n335 = ~\V133(9)  & n334;
  assign n336 = n234 & n235;
  assign n337 = n326 & n336;
  assign n338 = ~n328 & ~n329;
  assign n339 = ~n337 & n338;
  assign n340 = ~n335 & n339;
  assign n341 = ~n332 & n340;
  assign n342 = ~\V133(10)  & n341;
  assign n343 = \V84(23)  & ~n342;
  assign n344 = n229 & n343;
  assign n345 = \V84(20)  & n252;
  assign n346 = ~n342 & n345;
  assign n347 = \V84(16)  & n249;
  assign n348 = ~n342 & n347;
  assign n349 = \V84(31)  & ~n228;
  assign n350 = ~n342 & n349;
  assign n351 = ~n264 & ~n342;
  assign n352 = ~n318 & ~n351;
  assign n353 = ~n350 & n352;
  assign n354 = ~n348 & n353;
  assign n355 = ~n346 & n354;
  assign \V197(31)  = n344 | ~n355;
  assign n357 = \V84(22)  & ~n342;
  assign n358 = n229 & n357;
  assign n359 = \V84(19)  & n252;
  assign n360 = ~n342 & n359;
  assign n361 = \V84(15)  & n249;
  assign n362 = ~n342 & n361;
  assign n363 = \V84(30)  & ~n228;
  assign n364 = ~n342 & n363;
  assign n365 = ~n294 & ~n351;
  assign n366 = ~n364 & n365;
  assign n367 = ~n362 & n366;
  assign n368 = ~n360 & n367;
  assign \V197(30)  = n358 | ~n368;
  assign n370 = ~\V133(2)  & n328;
  assign n371 = n236 & n329;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~\V133(10)  & n372;
  assign n374 = ~\V133(2)  & n232;
  assign n375 = ~\V133(1)  & n232;
  assign n376 = ~\V118(0)  & \V133(5) ;
  assign n377 = ~\V118(1)  & n376;
  assign n378 = n375 & n377;
  assign n379 = n374 & n378;
  assign n380 = \V116(3)  & n230;
  assign n381 = \V84(20)  & ~n373;
  assign n382 = ~n379 & ~n381;
  assign \V212(3)  = n380 | ~n382;
  assign n384 = \V116(2)  & n230;
  assign n385 = \V84(19)  & ~n373;
  assign n386 = ~n379 & ~n385;
  assign \V212(2)  = n384 | ~n386;
  assign n388 = \V116(5)  & n230;
  assign n389 = \V84(22)  & ~n373;
  assign n390 = ~n379 & ~n389;
  assign \V212(5)  = n388 | ~n390;
  assign n392 = \V116(4)  & n230;
  assign n393 = \V84(21)  & ~n373;
  assign n394 = ~n379 & ~n393;
  assign \V212(4)  = n392 | ~n394;
  assign n396 = \V116(1)  & n230;
  assign n397 = \V84(18)  & ~n373;
  assign n398 = ~n379 & ~n397;
  assign \V212(1)  = n396 | ~n398;
  assign n400 = \V116(0)  & n230;
  assign n401 = \V84(17)  & ~n373;
  assign n402 = ~n379 & ~n401;
  assign \V212(0)  = n400 | ~n402;
  assign n404 = \V116(7)  & n230;
  assign n405 = \V84(24)  & ~n373;
  assign n406 = ~n379 & ~n405;
  assign \V212(7)  = n404 | ~n406;
  assign n408 = \V116(6)  & n230;
  assign n409 = \V84(23)  & ~n373;
  assign n410 = ~n379 & ~n409;
  assign \V212(6)  = n408 | ~n410;
  assign n412 = ~\V133(10)  & n327;
  assign n413 = ~\V133(10)  & ~n327;
  assign n414 = ~n230 & ~n255;
  assign n415 = n217 & n414;
  assign n416 = \V121(16)  & ~\V133(8) ;
  assign n417 = n412 & n416;
  assign n418 = \V133(10)  & \V119(0) ;
  assign n419 = n413 & n414;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~n417 & n420;
  assign \V213(0)  = n415 | ~n421;
  assign n423 = \V116(9)  & n230;
  assign n424 = \V84(26)  & ~n373;
  assign n425 = ~n379 & ~n424;
  assign \V212(9)  = n423 | ~n425;
  assign n427 = \V116(8)  & n230;
  assign n428 = \V84(25)  & ~n373;
  assign n429 = ~n379 & ~n428;
  assign \V212(8)  = n427 | ~n429;
  assign n431 = \V47(8)  & ~\V133(2) ;
  assign n432 = n229 & n431;
  assign n433 = n240 & n432;
  assign n434 = \V47(5)  & ~\V133(2) ;
  assign n435 = n252 & n434;
  assign n436 = n240 & n435;
  assign n437 = \V47(1)  & ~\V133(2) ;
  assign n438 = n249 & n437;
  assign n439 = n240 & n438;
  assign n440 = ~\V133(2)  & \V47(16) ;
  assign n441 = ~n228 & n440;
  assign n442 = n240 & n441;
  assign n443 = ~\V133(2)  & ~n264;
  assign n444 = n240 & n443;
  assign n445 = \V47(8)  & ~n242;
  assign n446 = n229 & n445;
  assign n447 = \V47(5)  & ~n242;
  assign n448 = n252 & n447;
  assign n449 = \V47(1)  & ~n242;
  assign n450 = n249 & n449;
  assign n451 = \V47(16)  & ~n228;
  assign n452 = ~n242 & n451;
  assign n453 = \V116(16)  & n230;
  assign n454 = \V84(16)  & n258;
  assign n455 = ~n265 & ~n454;
  assign n456 = ~n453 & n455;
  assign n457 = ~n452 & n456;
  assign n458 = ~n450 & n457;
  assign n459 = ~n448 & n458;
  assign n460 = ~n446 & n459;
  assign n461 = ~n444 & n460;
  assign n462 = ~n442 & n461;
  assign n463 = ~n439 & n462;
  assign n464 = ~n436 & n463;
  assign \V150(0)  = n433 | ~n464;
  assign n466 = \V121(17)  & n412;
  assign n467 = \V133(10)  & \V122(0) ;
  assign n468 = n255 & ~n412;
  assign n469 = ~n467 & ~n468;
  assign \V214(0)  = n466 | ~n469;
  assign n471 = \V47(12)  & n243;
  assign n472 = \V47(5)  & n250;
  assign n473 = \V47(20)  & n251;
  assign n474 = \V47(9)  & n253;
  assign n475 = \V116(20)  & n230;
  assign n476 = \V84(20)  & n258;
  assign n477 = ~n265 & ~n476;
  assign n478 = ~n475 & n477;
  assign n479 = ~n474 & n478;
  assign n480 = ~n473 & n479;
  assign n481 = ~n472 & n480;
  assign \V165(3)  = n471 | ~n481;
  assign n483 = \V47(11)  & n243;
  assign n484 = \V47(4)  & n250;
  assign n485 = \V47(19)  & n251;
  assign n486 = \V47(8)  & n253;
  assign n487 = \V116(19)  & n230;
  assign n488 = \V84(19)  & n258;
  assign n489 = ~n265 & ~n488;
  assign n490 = ~n487 & n489;
  assign n491 = ~n486 & n490;
  assign n492 = ~n485 & n491;
  assign n493 = ~n484 & n492;
  assign \V165(2)  = n483 | ~n493;
  assign n495 = \V47(14)  & n243;
  assign n496 = \V47(7)  & n250;
  assign n497 = \V47(22)  & n251;
  assign n498 = \V47(11)  & n253;
  assign n499 = \V116(22)  & n230;
  assign n500 = \V84(22)  & n258;
  assign n501 = ~n265 & ~n500;
  assign n502 = ~n499 & n501;
  assign n503 = ~n498 & n502;
  assign n504 = ~n497 & n503;
  assign n505 = ~n496 & n504;
  assign \V165(5)  = n495 | ~n505;
  assign n507 = \V47(13)  & n243;
  assign n508 = \V47(6)  & n250;
  assign n509 = \V47(21)  & n251;
  assign n510 = \V47(10)  & n253;
  assign n511 = \V116(21)  & n230;
  assign n512 = \V84(21)  & n258;
  assign n513 = ~n265 & ~n512;
  assign n514 = ~n511 & n513;
  assign n515 = ~n510 & n514;
  assign n516 = ~n509 & n515;
  assign n517 = ~n508 & n516;
  assign \V165(4)  = n507 | ~n517;
  assign n519 = \V47(10)  & n243;
  assign n520 = \V47(3)  & n250;
  assign n521 = \V47(18)  & n251;
  assign n522 = \V47(7)  & n253;
  assign n523 = \V116(18)  & n230;
  assign n524 = \V84(18)  & n258;
  assign n525 = ~n265 & ~n524;
  assign n526 = ~n523 & n525;
  assign n527 = ~n522 & n526;
  assign n528 = ~n521 & n527;
  assign n529 = ~n520 & n528;
  assign \V165(1)  = n519 | ~n529;
  assign n531 = \V47(9)  & n243;
  assign n532 = \V47(2)  & n250;
  assign n533 = \V47(17)  & n251;
  assign n534 = \V47(6)  & n253;
  assign n535 = \V116(17)  & n230;
  assign n536 = \V84(17)  & n258;
  assign n537 = ~n265 & ~n536;
  assign n538 = ~n535 & n537;
  assign n539 = ~n534 & n538;
  assign n540 = ~n533 & n539;
  assign n541 = ~n532 & n540;
  assign \V165(0)  = n531 | ~n541;
  assign n543 = \V116(11)  & n230;
  assign n544 = \V84(28)  & ~n373;
  assign n545 = ~n379 & ~n544;
  assign \V212(11)  = n543 | ~n545;
  assign n547 = \V116(10)  & n230;
  assign n548 = \V84(27)  & ~n373;
  assign n549 = ~n379 & ~n548;
  assign \V212(10)  = n547 | ~n549;
  assign n551 = \V116(13)  & n230;
  assign n552 = \V84(30)  & ~n373;
  assign n553 = ~n379 & ~n552;
  assign \V212(13)  = n551 | ~n553;
  assign n555 = \V47(16)  & n243;
  assign n556 = \V47(9)  & n250;
  assign n557 = \V47(24)  & n251;
  assign n558 = \V47(13)  & n253;
  assign n559 = \V116(24)  & n230;
  assign n560 = \V84(24)  & n258;
  assign n561 = ~n265 & ~n560;
  assign n562 = ~n559 & n561;
  assign n563 = ~n558 & n562;
  assign n564 = ~n557 & n563;
  assign n565 = ~n556 & n564;
  assign \V165(7)  = n555 | ~n565;
  assign n567 = \V116(12)  & n230;
  assign n568 = \V84(29)  & ~n373;
  assign n569 = ~n379 & ~n568;
  assign \V212(12)  = n567 | ~n569;
  assign n571 = \V47(15)  & n243;
  assign n572 = \V47(8)  & n250;
  assign n573 = \V47(23)  & n251;
  assign n574 = \V47(12)  & n253;
  assign n575 = \V116(23)  & n230;
  assign n576 = \V84(23)  & n258;
  assign n577 = ~n265 & ~n576;
  assign n578 = ~n575 & n577;
  assign n579 = ~n574 & n578;
  assign n580 = ~n573 & n579;
  assign n581 = ~n572 & n580;
  assign \V165(6)  = n571 | ~n581;
  assign n583 = \V47(18)  & n243;
  assign n584 = \V47(11)  & n250;
  assign n585 = \V47(26)  & n251;
  assign n586 = \V47(15)  & n253;
  assign n587 = \V116(26)  & n230;
  assign n588 = \V84(26)  & n258;
  assign n589 = ~n265 & ~n588;
  assign n590 = ~n587 & n589;
  assign n591 = ~n586 & n590;
  assign n592 = ~n585 & n591;
  assign n593 = ~n584 & n592;
  assign \V165(9)  = n583 | ~n593;
  assign n595 = \V116(14)  & n230;
  assign n596 = \V84(31)  & ~n373;
  assign n597 = ~n379 & ~n596;
  assign \V212(14)  = n595 | ~n597;
  assign n599 = \V47(17)  & n243;
  assign n600 = \V47(10)  & n250;
  assign n601 = \V47(25)  & n251;
  assign n602 = \V47(14)  & n253;
  assign n603 = \V116(25)  & n230;
  assign n604 = \V84(25)  & n258;
  assign n605 = ~n265 & ~n604;
  assign n606 = ~n603 & n605;
  assign n607 = ~n602 & n606;
  assign n608 = ~n601 & n607;
  assign n609 = ~n600 & n608;
  assign \V165(8)  = n599 | ~n609;
  assign n611 = ~n235 & n413;
  assign n612 = n249 & ~n611;
  assign n613 = ~n228 & ~n611;
  assign n614 = n252 & ~n611;
  assign n615 = ~n264 & ~n611;
  assign n616 = \V15(5)  & n612;
  assign n617 = \V47(6)  & n613;
  assign n618 = \V84(6)  & n614;
  assign n619 = ~n615 & ~n618;
  assign n620 = ~n617 & n619;
  assign n621 = ~n408 & n620;
  assign \V142(3)  = n616 | ~n621;
  assign n623 = \V15(4)  & n612;
  assign n624 = \V47(5)  & n613;
  assign n625 = \V84(5)  & n614;
  assign n626 = ~n615 & ~n625;
  assign n627 = ~n624 & n626;
  assign n628 = ~n388 & n627;
  assign \V142(2)  = n623 | ~n628;
  assign n630 = n229 & ~n611;
  assign n631 = \V47(0)  & n630;
  assign n632 = \V15(7)  & n612;
  assign n633 = \V47(8)  & n613;
  assign n634 = \V84(8)  & n614;
  assign n635 = ~n615 & ~n634;
  assign n636 = ~n633 & n635;
  assign n637 = ~n427 & n636;
  assign n638 = ~n632 & n637;
  assign \V142(5)  = n631 | ~n638;
  assign n640 = \V15(6)  & n612;
  assign n641 = \V47(7)  & n613;
  assign n642 = \V84(7)  & n614;
  assign n643 = ~n615 & ~n642;
  assign n644 = ~n641 & n643;
  assign n645 = ~n404 & n644;
  assign \V142(4)  = n640 | ~n645;
  assign n647 = \V15(3)  & n612;
  assign n648 = \V47(4)  & n613;
  assign n649 = \V84(4)  & n614;
  assign n650 = ~n615 & ~n649;
  assign n651 = ~n648 & n650;
  assign n652 = ~n392 & n651;
  assign \V142(1)  = n647 | ~n652;
  assign n654 = \V15(2)  & n612;
  assign n655 = \V47(3)  & n613;
  assign n656 = \V84(3)  & n614;
  assign n657 = ~n615 & ~n656;
  assign n658 = ~n655 & n657;
  assign n659 = ~n380 & n658;
  assign \V142(0)  = n654 | ~n659;
  assign n661 = \V84(9)  & n252;
  assign n662 = n264 & ~n661;
  assign n663 = \V47(1)  & ~n413;
  assign n664 = n229 & n663;
  assign n665 = \V47(1)  & n233;
  assign n666 = n229 & n665;
  assign n667 = \V15(8)  & ~n413;
  assign n668 = n249 & n667;
  assign n669 = \V15(8)  & n233;
  assign n670 = n249 & n669;
  assign n671 = \V47(9)  & ~n228;
  assign n672 = ~n413 & n671;
  assign n673 = n233 & n671;
  assign n674 = ~n413 & ~n662;
  assign n675 = n233 & ~n662;
  assign n676 = ~n423 & ~n675;
  assign n677 = ~n674 & n676;
  assign n678 = ~n673 & n677;
  assign n679 = ~n672 & n678;
  assign n680 = ~n670 & n679;
  assign n681 = ~n668 & n680;
  assign n682 = ~n666 & n681;
  assign \V143(0)  = n664 | ~n682;
  assign n684 = \V84(19)  & ~n342;
  assign n685 = n229 & n684;
  assign n686 = \V84(16)  & n252;
  assign n687 = ~n342 & n686;
  assign n688 = \V84(12)  & n249;
  assign n689 = ~n342 & n688;
  assign n690 = \V84(27)  & ~n228;
  assign n691 = ~n342 & n690;
  assign n692 = ~n282 & ~n351;
  assign n693 = ~n691 & n692;
  assign n694 = ~n689 & n693;
  assign n695 = ~n687 & n694;
  assign \V197(27)  = n685 | ~n695;
  assign n697 = \V84(18)  & ~n342;
  assign n698 = n229 & n697;
  assign n699 = \V84(15)  & n252;
  assign n700 = ~n342 & n699;
  assign n701 = \V84(11)  & n249;
  assign n702 = ~n342 & n701;
  assign n703 = \V84(26)  & ~n228;
  assign n704 = ~n342 & n703;
  assign n705 = ~n351 & ~n587;
  assign n706 = ~n704 & n705;
  assign n707 = ~n702 & n706;
  assign n708 = ~n700 & n707;
  assign \V197(26)  = n698 | ~n708;
  assign n710 = \V84(21)  & ~n342;
  assign n711 = n229 & n710;
  assign n712 = \V84(18)  & n252;
  assign n713 = ~n342 & n712;
  assign n714 = \V84(14)  & n249;
  assign n715 = ~n342 & n714;
  assign n716 = \V84(29)  & ~n228;
  assign n717 = ~n342 & n716;
  assign n718 = ~n306 & ~n351;
  assign n719 = ~n717 & n718;
  assign n720 = ~n715 & n719;
  assign n721 = ~n713 & n720;
  assign \V197(29)  = n711 | ~n721;
  assign n723 = \V84(20)  & ~n342;
  assign n724 = n229 & n723;
  assign n725 = \V84(17)  & n252;
  assign n726 = ~n342 & n725;
  assign n727 = \V84(13)  & n249;
  assign n728 = ~n342 & n727;
  assign n729 = \V84(28)  & ~n228;
  assign n730 = ~n342 & n729;
  assign n731 = ~n270 & ~n351;
  assign n732 = ~n730 & n731;
  assign n733 = ~n728 & n732;
  assign n734 = ~n726 & n733;
  assign \V197(28)  = n724 | ~n734;
  assign n736 = \V47(3)  & n630;
  assign n737 = \V15(10)  & n612;
  assign n738 = \V47(11)  & n613;
  assign n739 = \V84(11)  & n614;
  assign n740 = ~n615 & ~n739;
  assign n741 = ~n738 & n740;
  assign n742 = ~n543 & n741;
  assign n743 = ~n737 & n742;
  assign \V145(1)  = n736 | ~n743;
  assign n745 = \V47(2)  & n630;
  assign n746 = \V15(9)  & n612;
  assign n747 = \V47(10)  & n613;
  assign n748 = \V84(10)  & n614;
  assign n749 = ~n615 & ~n748;
  assign n750 = ~n747 & n749;
  assign n751 = ~n547 & n750;
  assign n752 = ~n746 & n751;
  assign \V145(0)  = n745 | ~n752;
  assign n754 = \V84(13)  & ~n342;
  assign n755 = n229 & n754;
  assign n756 = \V84(10)  & n252;
  assign n757 = ~n342 & n756;
  assign n758 = \V84(6)  & n249;
  assign n759 = ~n342 & n758;
  assign n760 = \V84(21)  & ~n228;
  assign n761 = ~n342 & n760;
  assign n762 = ~n351 & ~n511;
  assign n763 = ~n761 & n762;
  assign n764 = ~n759 & n763;
  assign n765 = ~n757 & n764;
  assign \V197(21)  = n755 | ~n765;
  assign n767 = \V84(12)  & ~n342;
  assign n768 = n229 & n767;
  assign n769 = \V84(5)  & n249;
  assign n770 = ~n342 & n769;
  assign n771 = \V84(20)  & ~n228;
  assign n772 = ~n342 & n771;
  assign n773 = ~n342 & ~n662;
  assign n774 = ~n475 & ~n773;
  assign n775 = ~n772 & n774;
  assign n776 = ~n770 & n775;
  assign \V197(20)  = n768 | ~n776;
  assign n778 = \V84(15)  & ~n342;
  assign n779 = n229 & n778;
  assign n780 = \V84(12)  & n252;
  assign n781 = ~n342 & n780;
  assign n782 = \V84(8)  & n249;
  assign n783 = ~n342 & n782;
  assign n784 = \V84(23)  & ~n228;
  assign n785 = ~n342 & n784;
  assign n786 = ~n351 & ~n575;
  assign n787 = ~n785 & n786;
  assign n788 = ~n783 & n787;
  assign n789 = ~n781 & n788;
  assign \V197(23)  = n779 | ~n789;
  assign n791 = \V84(14)  & ~n342;
  assign n792 = n229 & n791;
  assign n793 = \V84(11)  & n252;
  assign n794 = ~n342 & n793;
  assign n795 = \V84(7)  & n249;
  assign n796 = ~n342 & n795;
  assign n797 = \V84(22)  & ~n228;
  assign n798 = ~n342 & n797;
  assign n799 = ~n351 & ~n499;
  assign n800 = ~n798 & n799;
  assign n801 = ~n796 & n800;
  assign n802 = ~n794 & n801;
  assign \V197(22)  = n792 | ~n802;
  assign n804 = \V84(17)  & ~n342;
  assign n805 = n229 & n804;
  assign n806 = \V84(14)  & n252;
  assign n807 = ~n342 & n806;
  assign n808 = \V84(10)  & n249;
  assign n809 = ~n342 & n808;
  assign n810 = \V84(25)  & ~n228;
  assign n811 = ~n342 & n810;
  assign n812 = ~n351 & ~n603;
  assign n813 = ~n811 & n812;
  assign n814 = ~n809 & n813;
  assign n815 = ~n807 & n814;
  assign \V197(25)  = n805 | ~n815;
  assign n817 = \V84(16)  & ~n342;
  assign n818 = n229 & n817;
  assign n819 = \V84(13)  & n252;
  assign n820 = ~n342 & n819;
  assign n821 = \V84(9)  & n249;
  assign n822 = ~n342 & n821;
  assign n823 = \V84(24)  & ~n228;
  assign n824 = ~n342 & n823;
  assign n825 = ~n351 & ~n559;
  assign n826 = ~n824 & n825;
  assign n827 = ~n822 & n826;
  assign n828 = ~n820 & n827;
  assign \V197(24)  = n818 | ~n828;
  assign n830 = \V47(4)  & n229;
  assign n831 = n240 & n830;
  assign n832 = \V47(1)  & n252;
  assign n833 = n240 & n832;
  assign n834 = \V15(11)  & n249;
  assign n835 = n240 & n834;
  assign n836 = \V47(12)  & ~n228;
  assign n837 = n240 & n836;
  assign n838 = \V84(12)  & ~n236;
  assign n839 = n258 & n838;
  assign n840 = \V47(4)  & ~n239;
  assign n841 = n229 & n840;
  assign n842 = \V47(1)  & ~n239;
  assign n843 = n252 & n842;
  assign n844 = \V15(11)  & ~n239;
  assign n845 = n249 & n844;
  assign n846 = ~n239 & n836;
  assign n847 = \V116(12)  & ~n236;
  assign n848 = n230 & n847;
  assign n849 = n240 & ~n264;
  assign n850 = ~n239 & ~n264;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n848 & n851;
  assign n853 = ~n846 & n852;
  assign n854 = ~n845 & n853;
  assign n855 = ~n843 & n854;
  assign n856 = ~n841 & n855;
  assign n857 = ~n839 & n856;
  assign n858 = ~n837 & n857;
  assign n859 = ~n835 & n858;
  assign n860 = ~n833 & n859;
  assign \V146(0)  = n831 | ~n860;
  assign n862 = \V84(9)  & ~n342;
  assign n863 = n229 & n862;
  assign n864 = \V84(6)  & n252;
  assign n865 = ~n342 & n864;
  assign n866 = \V84(2)  & n249;
  assign n867 = ~n342 & n866;
  assign n868 = \V84(17)  & ~n228;
  assign n869 = ~n342 & n868;
  assign n870 = ~n351 & ~n535;
  assign n871 = ~n869 & n870;
  assign n872 = ~n867 & n871;
  assign n873 = ~n865 & n872;
  assign \V197(17)  = n863 | ~n873;
  assign n875 = \V84(8)  & ~n342;
  assign n876 = n229 & n875;
  assign n877 = \V84(5)  & n252;
  assign n878 = ~n342 & n877;
  assign n879 = \V84(1)  & n249;
  assign n880 = ~n342 & n879;
  assign n881 = \V84(16)  & ~n228;
  assign n882 = ~n342 & n881;
  assign n883 = ~n351 & ~n453;
  assign n884 = ~n882 & n883;
  assign n885 = ~n880 & n884;
  assign n886 = ~n878 & n885;
  assign \V197(16)  = n876 | ~n886;
  assign n888 = \V84(11)  & ~n342;
  assign n889 = n229 & n888;
  assign n890 = \V84(8)  & n252;
  assign n891 = ~n342 & n890;
  assign n892 = \V84(4)  & n249;
  assign n893 = ~n342 & n892;
  assign n894 = \V84(19)  & ~n228;
  assign n895 = ~n342 & n894;
  assign n896 = ~n351 & ~n487;
  assign n897 = ~n895 & n896;
  assign n898 = ~n893 & n897;
  assign n899 = ~n891 & n898;
  assign \V197(19)  = n889 | ~n899;
  assign n901 = \V84(10)  & ~n342;
  assign n902 = n229 & n901;
  assign n903 = \V84(7)  & n252;
  assign n904 = ~n342 & n903;
  assign n905 = \V84(3)  & n249;
  assign n906 = ~n342 & n905;
  assign n907 = \V84(18)  & ~n228;
  assign n908 = ~n342 & n907;
  assign n909 = ~n351 & ~n523;
  assign n910 = ~n908 & n909;
  assign n911 = ~n906 & n910;
  assign n912 = ~n904 & n911;
  assign \V197(18)  = n902 | ~n912;
  assign n914 = n328 & n412;
  assign n915 = \V84(0)  & ~n914;
  assign n916 = ~n413 & n915;
  assign n917 = ~n215 & n916;
  assign n918 = ~\V133(10)  & ~n914;
  assign n919 = ~n413 & n918;
  assign n920 = ~n215 & n919;
  assign n921 = ~\V133(10)  & \V48(0) ;
  assign n922 = ~n413 & n921;
  assign n923 = \V49(0)  & n232;
  assign n924 = ~n400 & ~n923;
  assign n925 = ~n922 & n924;
  assign n926 = ~n920 & n925;
  assign \V134(0)  = n917 | ~n926;
  assign n928 = \V47(27)  & ~n342;
  assign n929 = n229 & n928;
  assign n930 = \V47(24)  & n252;
  assign n931 = ~n342 & n930;
  assign n932 = \V47(20)  & n249;
  assign n933 = ~n342 & n932;
  assign n934 = \V84(3)  & ~n228;
  assign n935 = ~n342 & n934;
  assign n936 = ~n351 & ~n380;
  assign n937 = ~n935 & n936;
  assign n938 = ~n933 & n937;
  assign n939 = ~n931 & n938;
  assign \V197(3)  = n929 | ~n939;
  assign n941 = \V84(3)  & ~n342;
  assign n942 = n229 & n941;
  assign n943 = \V84(0)  & n252;
  assign n944 = ~n342 & n943;
  assign n945 = \V47(28)  & n249;
  assign n946 = ~n342 & n945;
  assign n947 = \V84(11)  & ~n228;
  assign n948 = ~n342 & n947;
  assign n949 = ~n351 & ~n543;
  assign n950 = ~n948 & n949;
  assign n951 = ~n946 & n950;
  assign n952 = ~n944 & n951;
  assign \V197(11)  = n942 | ~n952;
  assign n954 = \V47(26)  & ~n342;
  assign n955 = n229 & n954;
  assign n956 = \V47(23)  & n252;
  assign n957 = ~n342 & n956;
  assign n958 = \V47(19)  & n249;
  assign n959 = ~n342 & n958;
  assign n960 = \V84(2)  & ~n228;
  assign n961 = ~n342 & n960;
  assign n962 = ~n351 & ~n384;
  assign n963 = ~n961 & n962;
  assign n964 = ~n959 & n963;
  assign n965 = ~n957 & n964;
  assign \V197(2)  = n955 | ~n965;
  assign n967 = \V84(2)  & ~n342;
  assign n968 = n229 & n967;
  assign n969 = \V47(31)  & n252;
  assign n970 = ~n342 & n969;
  assign n971 = \V47(27)  & n249;
  assign n972 = ~n342 & n971;
  assign n973 = \V84(10)  & ~n228;
  assign n974 = ~n342 & n973;
  assign n975 = ~n351 & ~n547;
  assign n976 = ~n974 & n975;
  assign n977 = ~n972 & n976;
  assign n978 = ~n970 & n977;
  assign \V197(10)  = n968 | ~n978;
  assign n980 = \V47(29)  & ~n342;
  assign n981 = n229 & n980;
  assign n982 = \V47(26)  & n252;
  assign n983 = ~n342 & n982;
  assign n984 = \V47(22)  & n249;
  assign n985 = ~n342 & n984;
  assign n986 = \V84(5)  & ~n228;
  assign n987 = ~n342 & n986;
  assign n988 = ~n351 & ~n388;
  assign n989 = ~n987 & n988;
  assign n990 = ~n985 & n989;
  assign n991 = ~n983 & n990;
  assign \V197(5)  = n981 | ~n991;
  assign n993 = \V84(2)  & n252;
  assign n994 = n264 & ~n993;
  assign n995 = \V84(5)  & ~n342;
  assign n996 = n229 & n995;
  assign n997 = \V47(30)  & n249;
  assign n998 = ~n342 & n997;
  assign n999 = \V84(13)  & ~n228;
  assign n1000 = ~n342 & n999;
  assign n1001 = ~n342 & ~n994;
  assign n1002 = ~n551 & ~n1001;
  assign n1003 = ~n1000 & n1002;
  assign n1004 = ~n998 & n1003;
  assign \V197(13)  = n996 | ~n1004;
  assign n1006 = \V47(7)  & n243;
  assign n1007 = \V15(14)  & n250;
  assign n1008 = \V47(15)  & n251;
  assign n1009 = \V47(4)  & n253;
  assign n1010 = \V116(15)  & n230;
  assign n1011 = \V84(15)  & n258;
  assign n1012 = ~n265 & ~n1011;
  assign n1013 = ~n1010 & n1012;
  assign n1014 = ~n1009 & n1013;
  assign n1015 = ~n1008 & n1014;
  assign n1016 = ~n1007 & n1015;
  assign \V149(2)  = n1006 | ~n1016;
  assign n1018 = \V47(28)  & ~n342;
  assign n1019 = n229 & n1018;
  assign n1020 = \V47(25)  & n252;
  assign n1021 = ~n342 & n1020;
  assign n1022 = \V47(21)  & n249;
  assign n1023 = ~n342 & n1022;
  assign n1024 = \V84(4)  & ~n228;
  assign n1025 = ~n342 & n1024;
  assign n1026 = ~n351 & ~n392;
  assign n1027 = ~n1025 & n1026;
  assign n1028 = ~n1023 & n1027;
  assign n1029 = ~n1021 & n1028;
  assign \V197(4)  = n1019 | ~n1029;
  assign n1031 = \V84(1)  & n252;
  assign n1032 = n264 & ~n1031;
  assign n1033 = \V84(4)  & ~n342;
  assign n1034 = n229 & n1033;
  assign n1035 = \V47(29)  & n249;
  assign n1036 = ~n342 & n1035;
  assign n1037 = \V84(12)  & ~n228;
  assign n1038 = ~n342 & n1037;
  assign n1039 = ~n342 & ~n1032;
  assign n1040 = ~n567 & ~n1039;
  assign n1041 = ~n1038 & n1040;
  assign n1042 = ~n1036 & n1041;
  assign \V197(12)  = n1034 | ~n1042;
  assign n1044 = \V84(7)  & ~n342;
  assign n1045 = n229 & n1044;
  assign n1046 = \V84(4)  & n252;
  assign n1047 = ~n342 & n1046;
  assign n1048 = \V84(0)  & n249;
  assign n1049 = ~n342 & n1048;
  assign n1050 = \V84(15)  & ~n228;
  assign n1051 = ~n342 & n1050;
  assign n1052 = ~n351 & ~n1010;
  assign n1053 = ~n1051 & n1052;
  assign n1054 = ~n1049 & n1053;
  assign n1055 = ~n1047 & n1054;
  assign \V197(15)  = n1045 | ~n1055;
  assign n1057 = \V84(6)  & ~n342;
  assign n1058 = n229 & n1057;
  assign n1059 = \V84(3)  & n252;
  assign n1060 = ~n342 & n1059;
  assign n1061 = \V47(31)  & n249;
  assign n1062 = ~n342 & n1061;
  assign n1063 = \V84(14)  & ~n228;
  assign n1064 = ~n342 & n1063;
  assign n1065 = ~n351 & ~n595;
  assign n1066 = ~n1064 & n1065;
  assign n1067 = ~n1062 & n1066;
  assign n1068 = ~n1060 & n1067;
  assign \V197(14)  = n1058 | ~n1068;
  assign n1070 = \V47(25)  & ~n342;
  assign n1071 = n229 & n1070;
  assign n1072 = \V47(22)  & n252;
  assign n1073 = ~n342 & n1072;
  assign n1074 = \V47(18)  & n249;
  assign n1075 = ~n342 & n1074;
  assign n1076 = \V84(1)  & ~n228;
  assign n1077 = ~n342 & n1076;
  assign n1078 = ~n351 & ~n396;
  assign n1079 = ~n1077 & n1078;
  assign n1080 = ~n1075 & n1079;
  assign n1081 = ~n1073 & n1080;
  assign \V197(1)  = n1071 | ~n1081;
  assign n1083 = \V47(24)  & ~n342;
  assign n1084 = n229 & n1083;
  assign n1085 = \V47(21)  & n252;
  assign n1086 = ~n342 & n1085;
  assign n1087 = \V47(17)  & n249;
  assign n1088 = ~n342 & n1087;
  assign n1089 = \V84(0)  & ~n228;
  assign n1090 = ~n342 & n1089;
  assign n1091 = ~n351 & ~n400;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = ~n1088 & n1092;
  assign n1094 = ~n1086 & n1093;
  assign \V197(0)  = n1084 | ~n1094;
  assign n1096 = \V47(6)  & n243;
  assign n1097 = \V15(13)  & n250;
  assign n1098 = \V47(14)  & n251;
  assign n1099 = \V47(3)  & n253;
  assign n1100 = \V84(14)  & n258;
  assign n1101 = ~n265 & ~n1100;
  assign n1102 = ~n595 & n1101;
  assign n1103 = ~n1099 & n1102;
  assign n1104 = ~n1098 & n1103;
  assign n1105 = ~n1097 & n1104;
  assign \V149(1)  = n1096 | ~n1105;
  assign n1107 = \V47(5)  & n243;
  assign n1108 = \V15(12)  & n250;
  assign n1109 = \V47(13)  & n251;
  assign n1110 = \V47(2)  & n253;
  assign n1111 = \V84(13)  & n258;
  assign n1112 = ~n265 & ~n1111;
  assign n1113 = ~n551 & n1112;
  assign n1114 = ~n1110 & n1113;
  assign n1115 = ~n1109 & n1114;
  assign n1116 = ~n1108 & n1115;
  assign \V149(0)  = n1107 | ~n1116;
  assign n1118 = ~\V133(8)  & n233;
  assign n1119 = n226 & n1118;
  assign n1120 = ~\V133(8)  & n327;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~\V133(10)  & n1121;
  assign n1123 = ~\V133(8)  & n413;
  assign n1124 = ~n230 & ~n1123;
  assign n1125 = ~n374 & ~n375;
  assign n1126 = \V15(1)  & n249;
  assign n1127 = ~n1122 & n1126;
  assign n1128 = \V47(2)  & ~n228;
  assign n1129 = ~n1122 & n1128;
  assign n1130 = \V52(0)  & ~n1125;
  assign n1131 = ~n1124 & n1130;
  assign n1132 = ~n994 & ~n1122;
  assign n1133 = ~n384 & ~n1132;
  assign n1134 = ~n1131 & n1133;
  assign n1135 = ~n1129 & n1134;
  assign \V136(1)  = n1127 | ~n1135;
  assign n1137 = \V47(31)  & ~n342;
  assign n1138 = n229 & n1137;
  assign n1139 = \V47(28)  & n252;
  assign n1140 = ~n342 & n1139;
  assign n1141 = \V47(24)  & n249;
  assign n1142 = ~n342 & n1141;
  assign n1143 = \V84(7)  & ~n228;
  assign n1144 = ~n342 & n1143;
  assign n1145 = ~n351 & ~n404;
  assign n1146 = ~n1144 & n1145;
  assign n1147 = ~n1142 & n1146;
  assign n1148 = ~n1140 & n1147;
  assign \V197(7)  = n1138 | ~n1148;
  assign n1150 = \V50(0)  & ~n230;
  assign n1151 = n217 & n1150;
  assign n1152 = \V15(0)  & n249;
  assign n1153 = ~n1122 & n1152;
  assign n1154 = \V47(1)  & ~n228;
  assign n1155 = ~n1122 & n1154;
  assign n1156 = \V51(0)  & ~n1125;
  assign n1157 = ~n1124 & n1156;
  assign n1158 = ~n1032 & ~n1122;
  assign n1159 = ~n396 & ~n1158;
  assign n1160 = ~n1157 & n1159;
  assign n1161 = ~n1155 & n1160;
  assign n1162 = ~n1153 & n1161;
  assign \V136(0)  = n1151 | ~n1162;
  assign n1164 = \V47(30)  & ~n342;
  assign n1165 = n229 & n1164;
  assign n1166 = \V47(27)  & n252;
  assign n1167 = ~n342 & n1166;
  assign n1168 = \V47(23)  & n249;
  assign n1169 = ~n342 & n1168;
  assign n1170 = \V84(6)  & ~n228;
  assign n1171 = ~n342 & n1170;
  assign n1172 = ~n351 & ~n408;
  assign n1173 = ~n1171 & n1172;
  assign n1174 = ~n1169 & n1173;
  assign n1175 = ~n1167 & n1174;
  assign \V197(6)  = n1165 | ~n1175;
  assign n1177 = \V84(1)  & ~n342;
  assign n1178 = n229 & n1177;
  assign n1179 = \V47(30)  & n252;
  assign n1180 = ~n342 & n1179;
  assign n1181 = \V47(26)  & n249;
  assign n1182 = ~n342 & n1181;
  assign n1183 = \V84(9)  & ~n228;
  assign n1184 = ~n342 & n1183;
  assign n1185 = ~n351 & ~n423;
  assign n1186 = ~n1184 & n1185;
  assign n1187 = ~n1182 & n1186;
  assign n1188 = ~n1180 & n1187;
  assign \V197(9)  = n1178 | ~n1188;
  assign n1190 = \V84(0)  & ~n342;
  assign n1191 = n229 & n1190;
  assign n1192 = \V47(29)  & n252;
  assign n1193 = ~n342 & n1192;
  assign n1194 = \V47(25)  & n249;
  assign n1195 = ~n342 & n1194;
  assign n1196 = \V84(8)  & ~n228;
  assign n1197 = ~n342 & n1196;
  assign n1198 = ~n351 & ~n427;
  assign n1199 = ~n1197 & n1198;
  assign n1200 = ~n1195 & n1199;
  assign n1201 = ~n1193 & n1200;
  assign \V197(8)  = n1191 | ~n1201;
endmodule


