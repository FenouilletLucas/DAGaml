// Benchmark "i10" written by ABC on Tue May 16 16:07:49 2017

module i10 ( 
    \V246(0) , \V229(3) , \V229(2) , \V229(5) , \V229(4) , \V38(0) ,
    \V171(0) , \V229(1) , \V229(0) , \V57(0) , \V248(0) , \V118(3) ,
    \V118(2) , \V118(5) , \V59(0) , \V118(4) , \V288(3) , \V288(2) ,
    \V78(0) , \V288(5) , \V118(1) , \V78(1) , \V302(0) , \V288(4) ,
    \V118(0) , \V78(2) , \V269(0) , \V78(3) , \V78(4) , \V288(1) ,
    \V78(5) , \V288(0) , \V118(7) , \V194(3) , \V118(6) , \V194(2) ,
    \V194(4) , \V288(7) , \V175(0) , \V288(6) , \V194(1) , \V194(0) ,
    \V177(0) , \V40(0) , \V1(0) , \V214(0) , \V42(0) , \V3(0) , \V101(0) ,
    \V271(0) , \V290(0) , \V216(0) , \V44(0) , \V5(0) , \V63(0) ,
    \V292(0) , \V46(0) , \V124(3) , \V7(0) , \V124(2) , \V124(5) ,
    \V65(0) , \V124(4) , \V84(0) , \V124(1) , \V84(1) , \V124(0) ,
    \V84(2) , \V275(0) , \V84(3) , \V84(4) , \V84(5) , \V294(0) ,
    \V239(3) , \V239(2) , \V239(4) , \V48(0) , \V9(0) , \V239(1) ,
    \V239(0) , \V67(0) , \V258(0) , \V277(0) , \V183(3) , \V183(2) ,
    \V183(5) , \V183(4) , \V183(1) , \V183(0) , \V69(0) , \V109(0) ,
    \V88(0) , \V88(1) , \V88(2) , \V279(0) , \V88(3) , \V149(3) ,
    \V149(2) , \V149(5) , \V149(4) , \V149(1) , \V10(0) , \V149(0) ,
    \V149(7) , \V149(6) , \V189(3) , \V12(0) , \V189(2) , \V189(5) ,
    \V203(0) , \V189(4) , \V189(1) , \V50(0) , \V189(0) , \V241(0) ,
    \V260(0) , \V14(0) , \V205(0) , \V33(0) , \V52(0) , \V243(0) ,
    \V71(0) , \V262(0) , \V16(0) , \V207(0) , \V35(0) , \V132(3) ,
    \V132(2) , \V245(0) , \V132(5) , \V132(4) , \V132(1) , \V132(0) ,
    \V132(7) , \V37(0) , \V132(6) , \V56(0) , \V247(0) , \V94(0) ,
    \V134(1) , \V94(1) , \V134(0) , \V39(0) , \V172(0) , \V268(3) ,
    \V268(2) , \V268(5) , \V268(4) , \V249(0) , \V301(0) , \V268(1) ,
    \V268(0) , \V174(0) , \V289(0) , \V213(3) , \V213(2) , \V213(5) ,
    \V213(4) , \V199(3) , \V199(2) , \V100(3) , \V213(1) , \V100(2) ,
    \V213(0) , \V199(4) , \V100(5) , \V41(0) , \V100(4) , \V2(0) ,
    \V199(1) , \V60(0) , \V199(0) , \V100(1) , \V100(0) , \V270(0) ,
    \V234(3) , \V234(2) , \V234(4) , \V215(0) , \V43(0) , \V4(0) ,
    \V234(1) , \V234(0) , \V62(0) , \V102(0) , \V32(11) , \V272(0) ,
    \V32(10) , \V291(0) , \V45(0) , \V6(0) , \V274(0) , \V293(0) ,
    \V257(3) , \V257(2) , \V257(5) , \V8(0) , \V257(4) , \V66(0) ,
    \V257(1) , \V257(0) , \V257(7) , \V257(6) , \V295(0) , \V108(3) ,
    \V108(2) , \V108(5) , \V108(4) , \V68(0) , \V108(1) , \V108(0) ,
    \V259(0) , \V165(3) , \V165(2) , \V278(0) , \V165(5) , \V165(4) ,
    \V165(1) , \V165(0) , \V165(7) , \V165(6) , \V11(0) , \V202(0) ,
    \V169(1) , \V169(0) , \V240(0) , \V223(3) , \V223(2) , \V13(0) ,
    \V223(5) , \V223(4) , \V204(0) , \V32(0) , \V32(1) , \V223(1) ,
    \V32(2) , \V223(0) , \V32(3) , \V51(0) , \V32(4) , \V32(5) , \V242(0) ,
    \V32(6) , \V70(0) , \V32(7) , \V110(0) , \V32(8) , \V261(0) , \V32(9) ,
    \V280(0) , \V15(0) , \V34(0) , \V53(0) , \V244(0) , \V91(0) , \V91(1) ,
    \V55(0) ,
    \V1213(10) , \V1213(11) , \V1440(0) , \V1833(0) , \V1536(0) ,
    \V321(2) , \V585(0) , \V1480(0) , \V1741(0) , \V1760(0) , \V603(0) ,
    \V1781(1) , \V1781(0) , \V1726(0) , V356, V357, \V1745(0) , \V1896(0) ,
    \V1613(1) , V373, V377, \V1613(0) , \V511(0) , \V1467(0) , \V1709(1) ,
    \V1709(0) , \V1709(3) , \V1709(2) , V432, \V1709(4) , \V1898(0) ,
    \V1392(0) , \V1243(7) , \V1243(6) , \V1243(9) , V512, \V1243(8) ,
    \V609(0) , V527, V537, V538, V539, V540, V541, V542, V543, V544, V545,
    V546, V547, V548, \V798(0) , \V1243(1) , V587, \V1243(0) , \V1243(3) ,
    \V1243(2) , \V572(3) , \V1243(5) , \V572(2) , \V1243(4) , \V572(5) ,
    \V572(4) , \V1281(0) , \V572(1) , V620, V621, \V572(0) , V630,
    \V1693(0) , V650, V651, V652, V653, V654, V655, V656, V657, \V591(0) ,
    \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) , \V1992(0) ,
    V707, \V423(0) , V763, V775, V778, V779, V780, V781, V782, V783, V784,
    V787, V789, V801, \V1864(0) , V966, \V597(0) , V986, \V1492(0) ,
    \V500(0) , \V1901(0) , \V1717(0) , \V634(0) , \V1213(7) , \V1439(0) ,
    \V1213(6) , \V1213(9) , \V1213(8) , \V375(0) , \V1213(1) , \V1213(0) ,
    \V1213(3) , \V1213(2) , \V1757(0) , \V1213(5) , \V1960(1) , \V1213(4) ,
    \V1960(0) , \V1512(1) , \V1512(3) , \V410(0) , \V1512(2) , V1256,
    V1257, V1258, V1259, \V1759(0) , V1260, V1261, V1262, V1263, V1264,
    V1265, V1266, V1267, \V1552(1) , \V398(0) , \V1552(0) , V1365, V1370,
    V1371, \V508(0) , V1372, V1373, V1374, V1375, V1378, V1380, V1382,
    V1384, V1386, \V1629(0) , V1387, \V1274(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V826(0) , V1470, \V435(0) , V1537, V1539,
    \V1968(0) , \V1297(1) , \V1481(0) , \V1297(0) , \V1297(3) , \V1297(2) ,
    \V1297(4) , \V640(0) , V1669, V1719, V1736, V1832, \V1897(0) ,
    \V1652(0) , \V1671(0) , \V1899(0) , \V1953(7) , \V1953(6) , \V1953(1) ,
    \V1953(0) , \V1953(3) , \V1953(2) , \V1953(5) , \V1953(4) , \V1451(0) ,
    \V1863(0) , \V1679(0) , \V1829(7) , \V1829(6) , \V1829(9) , \V1829(8) ,
    \V1771(1) , \V1620(0) , \V1771(0) , \V1829(1) , \V1829(0) , \V1829(3) ,
    \V1829(2) , \V1829(5) , \V1829(4) , \V1900(0) , \V1921(1) , \V1495(0) ,
    \V1921(0) , \V1921(3) , \V393(0) , \V1921(2) , \V1921(5) , \V1921(4) ,
    \V1459(0) , \V802(0) , \V821(0) , \V1758(0) , \V1645(0)   );
  input  \V246(0) , \V229(3) , \V229(2) , \V229(5) , \V229(4) , \V38(0) ,
    \V171(0) , \V229(1) , \V229(0) , \V57(0) , \V248(0) , \V118(3) ,
    \V118(2) , \V118(5) , \V59(0) , \V118(4) , \V288(3) , \V288(2) ,
    \V78(0) , \V288(5) , \V118(1) , \V78(1) , \V302(0) , \V288(4) ,
    \V118(0) , \V78(2) , \V269(0) , \V78(3) , \V78(4) , \V288(1) ,
    \V78(5) , \V288(0) , \V118(7) , \V194(3) , \V118(6) , \V194(2) ,
    \V194(4) , \V288(7) , \V175(0) , \V288(6) , \V194(1) , \V194(0) ,
    \V177(0) , \V40(0) , \V1(0) , \V214(0) , \V42(0) , \V3(0) , \V101(0) ,
    \V271(0) , \V290(0) , \V216(0) , \V44(0) , \V5(0) , \V63(0) ,
    \V292(0) , \V46(0) , \V124(3) , \V7(0) , \V124(2) , \V124(5) ,
    \V65(0) , \V124(4) , \V84(0) , \V124(1) , \V84(1) , \V124(0) ,
    \V84(2) , \V275(0) , \V84(3) , \V84(4) , \V84(5) , \V294(0) ,
    \V239(3) , \V239(2) , \V239(4) , \V48(0) , \V9(0) , \V239(1) ,
    \V239(0) , \V67(0) , \V258(0) , \V277(0) , \V183(3) , \V183(2) ,
    \V183(5) , \V183(4) , \V183(1) , \V183(0) , \V69(0) , \V109(0) ,
    \V88(0) , \V88(1) , \V88(2) , \V279(0) , \V88(3) , \V149(3) ,
    \V149(2) , \V149(5) , \V149(4) , \V149(1) , \V10(0) , \V149(0) ,
    \V149(7) , \V149(6) , \V189(3) , \V12(0) , \V189(2) , \V189(5) ,
    \V203(0) , \V189(4) , \V189(1) , \V50(0) , \V189(0) , \V241(0) ,
    \V260(0) , \V14(0) , \V205(0) , \V33(0) , \V52(0) , \V243(0) ,
    \V71(0) , \V262(0) , \V16(0) , \V207(0) , \V35(0) , \V132(3) ,
    \V132(2) , \V245(0) , \V132(5) , \V132(4) , \V132(1) , \V132(0) ,
    \V132(7) , \V37(0) , \V132(6) , \V56(0) , \V247(0) , \V94(0) ,
    \V134(1) , \V94(1) , \V134(0) , \V39(0) , \V172(0) , \V268(3) ,
    \V268(2) , \V268(5) , \V268(4) , \V249(0) , \V301(0) , \V268(1) ,
    \V268(0) , \V174(0) , \V289(0) , \V213(3) , \V213(2) , \V213(5) ,
    \V213(4) , \V199(3) , \V199(2) , \V100(3) , \V213(1) , \V100(2) ,
    \V213(0) , \V199(4) , \V100(5) , \V41(0) , \V100(4) , \V2(0) ,
    \V199(1) , \V60(0) , \V199(0) , \V100(1) , \V100(0) , \V270(0) ,
    \V234(3) , \V234(2) , \V234(4) , \V215(0) , \V43(0) , \V4(0) ,
    \V234(1) , \V234(0) , \V62(0) , \V102(0) , \V32(11) , \V272(0) ,
    \V32(10) , \V291(0) , \V45(0) , \V6(0) , \V274(0) , \V293(0) ,
    \V257(3) , \V257(2) , \V257(5) , \V8(0) , \V257(4) , \V66(0) ,
    \V257(1) , \V257(0) , \V257(7) , \V257(6) , \V295(0) , \V108(3) ,
    \V108(2) , \V108(5) , \V108(4) , \V68(0) , \V108(1) , \V108(0) ,
    \V259(0) , \V165(3) , \V165(2) , \V278(0) , \V165(5) , \V165(4) ,
    \V165(1) , \V165(0) , \V165(7) , \V165(6) , \V11(0) , \V202(0) ,
    \V169(1) , \V169(0) , \V240(0) , \V223(3) , \V223(2) , \V13(0) ,
    \V223(5) , \V223(4) , \V204(0) , \V32(0) , \V32(1) , \V223(1) ,
    \V32(2) , \V223(0) , \V32(3) , \V51(0) , \V32(4) , \V32(5) , \V242(0) ,
    \V32(6) , \V70(0) , \V32(7) , \V110(0) , \V32(8) , \V261(0) , \V32(9) ,
    \V280(0) , \V15(0) , \V34(0) , \V53(0) , \V244(0) , \V91(0) , \V91(1) ,
    \V55(0) ;
  output \V1213(10) , \V1213(11) , \V1440(0) , \V1833(0) , \V1536(0) ,
    \V321(2) , \V585(0) , \V1480(0) , \V1741(0) , \V1760(0) , \V603(0) ,
    \V1781(1) , \V1781(0) , \V1726(0) , V356, V357, \V1745(0) , \V1896(0) ,
    \V1613(1) , V373, V377, \V1613(0) , \V511(0) , \V1467(0) , \V1709(1) ,
    \V1709(0) , \V1709(3) , \V1709(2) , V432, \V1709(4) , \V1898(0) ,
    \V1392(0) , \V1243(7) , \V1243(6) , \V1243(9) , V512, \V1243(8) ,
    \V609(0) , V527, V537, V538, V539, V540, V541, V542, V543, V544, V545,
    V546, V547, V548, \V798(0) , \V1243(1) , V587, \V1243(0) , \V1243(3) ,
    \V1243(2) , \V572(3) , \V1243(5) , \V572(2) , \V1243(4) , \V572(5) ,
    \V572(4) , \V1281(0) , \V572(1) , V620, V621, \V572(0) , V630,
    \V1693(0) , V650, V651, V652, V653, V654, V655, V656, V657, \V591(0) ,
    \V572(7) , \V572(6) , \V572(9) , \V572(8) , \V1992(1) , \V1992(0) ,
    V707, \V423(0) , V763, V775, V778, V779, V780, V781, V782, V783, V784,
    V787, V789, V801, \V1864(0) , V966, \V597(0) , V986, \V1492(0) ,
    \V500(0) , \V1901(0) , \V1717(0) , \V634(0) , \V1213(7) , \V1439(0) ,
    \V1213(6) , \V1213(9) , \V1213(8) , \V375(0) , \V1213(1) , \V1213(0) ,
    \V1213(3) , \V1213(2) , \V1757(0) , \V1213(5) , \V1960(1) , \V1213(4) ,
    \V1960(0) , \V1512(1) , \V1512(3) , \V410(0) , \V1512(2) , V1256,
    V1257, V1258, V1259, \V1759(0) , V1260, V1261, V1262, V1263, V1264,
    V1265, V1266, V1267, \V1552(1) , \V398(0) , \V1552(0) , V1365, V1370,
    V1371, \V508(0) , V1372, V1373, V1374, V1375, V1378, V1380, V1382,
    V1384, V1386, \V1629(0) , V1387, \V1274(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V826(0) , V1470, \V435(0) , V1537, V1539,
    \V1968(0) , \V1297(1) , \V1481(0) , \V1297(0) , \V1297(3) , \V1297(2) ,
    \V1297(4) , \V640(0) , V1669, V1719, V1736, V1832, \V1897(0) ,
    \V1652(0) , \V1671(0) , \V1899(0) , \V1953(7) , \V1953(6) , \V1953(1) ,
    \V1953(0) , \V1953(3) , \V1953(2) , \V1953(5) , \V1953(4) , \V1451(0) ,
    \V1863(0) , \V1679(0) , \V1829(7) , \V1829(6) , \V1829(9) , \V1829(8) ,
    \V1771(1) , \V1620(0) , \V1771(0) , \V1829(1) , \V1829(0) , \V1829(3) ,
    \V1829(2) , \V1829(5) , \V1829(4) , \V1900(0) , \V1921(1) , \V1495(0) ,
    \V1921(0) , \V1921(3) , \V393(0) , \V1921(2) , \V1921(5) , \V1921(4) ,
    \V1459(0) , \V802(0) , \V821(0) , \V1758(0) , \V1645(0) ;
  wire n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n866, n867, n868, n869, n870, n871, n872, n874,
    n876, n877, n878, n879, n880, n881, n882, n884, n885, n886, n887, n888,
    n889, n890, n892, n893, n895, n896, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n912, n913, n914, n915, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n949, n950, n951, n952, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1724, n1725,
    n1726, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1736, n1737,
    n1738, n1739, n1741, n1742, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1759, n1760, n1761,
    n1762, n1763, n1765, n1766, n1768, n1769, n1770, n1771, n1772, n1774,
    n1775, n1776, n1777, n1778, n1780, n1781, n1782, n1783, n1784, n1787,
    n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1801, n1802, n1803, n1804, n1806, n1807, n1808, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1833,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1855, n1856,
    n1857, n1858, n1859, n1861, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1894, n1895, n1897, n1898, n1900, n1901, n1903,
    n1904, n1905, n1906, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2025,
    n2026, n2027, n2028, n2029, n2030, n2032, n2033, n2034, n2035, n2036,
    n2037, n2039, n2040, n2041, n2042, n2043, n2044, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2102, n2103, n2105, n2106, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2149, n2150, n2151, n2152, n2158, n2159, n2160, n2161,
    n2162, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2319, n2320, n2321,
    n2322, n2323, n2324, n2325, n2326, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2345, n2346, n2347, n2348, n2349, n2350, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2398,
    n2399, n2400, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2455, n2456, n2457, n2459, n2460, n2462, n2463, n2465, n2466,
    n2467, n2469, n2470, n2471, n2473, n2474, n2476, n2477, n2478, n2480,
    n2481, n2482, n2483, n2484, n2485, n2487, n2488, n2489, n2490, n2491,
    n2492, n2494, n2495, n2497, n2498, n2499, n2500, n2501, n2502, n2504,
    n2505, n2506, n2507, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2517, n2520, n2523, n2524, n2525, n2526, n2527, n2528, n2535, n2536,
    n2537, n2538, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2586, n2587, n2588, n2590, n2591, n2592, n2593,
    n2594, n2596, n2597, n2598, n2600, n2601, n2607, n2608, n2609, n2610,
    n2611, n2612, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2639, n2641, n2642, n2643, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2663, n2664, n2665, n2674, n2675,
    n2676, n2678, n2679, n2680, n2682, n2683, n2684, n2685, n2686, n2687,
    n2689, n2690, n2691, n2693, n2694, n2696, n2697, n2699, n2700, n2701,
    n2703, n2704, n2705, n2707, n2708, n2709, n2711, n2712, n2715, n2716,
    n2717, n2718, n2719, n2720, n2722, n2723, n2725, n2726, n2727, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2739, n2740, n2741,
    n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2759, n2760, n2763, n2764, n2765, n2766, n2767,
    n2768, n2770, n2774, n2775, n2777, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2805, n2806, n2808, n2809, n2811, n2812, n2814, n2815, n2817, n2818,
    n2820, n2822, n2823, n2824, n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2854, n2855, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2866, n2867, n2869, n2870, n2871, n2872, n2873, n2875, n2876,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2887, n2888,
    n2890, n2891, n2893, n2894, n2896, n2897, n2899, n2900, n2902, n2903,
    n2904, n2905, n2906, n2908, n2909, n2911, n2912, n2914, n2916, n2917,
    n2919, n2920, n2922, n2923, n2925, n2926, n2928, n2930, n2931, n2932,
    n2933, n2935, n2936, n2938, n2939, n2940;
  assign n482 = \V149(2)  & ~\V149(0) ;
  assign n483 = \V149(1)  & n482;
  assign n484 = ~\V149(3)  & ~\V149(4) ;
  assign n485 = n483 & n484;
  assign n486 = \V149(3)  & n483;
  assign n487 = ~\V165(5)  & ~\V165(4) ;
  assign n488 = ~\V165(6)  & \V70(0) ;
  assign n489 = \V165(3)  & n488;
  assign n490 = n487 & n489;
  assign n491 = \V149(5)  & \V149(4) ;
  assign n492 = \V149(1)  & ~\V149(0) ;
  assign n493 = ~\V149(2)  & n492;
  assign n494 = ~\V149(3)  & n493;
  assign n495 = \V149(6)  & n494;
  assign n496 = n491 & n495;
  assign \V802(0)  = \V52(0)  | \V51(0) ;
  assign n498 = ~\V149(3)  & \V149(4) ;
  assign n499 = n483 & n498;
  assign n500 = ~\V149(2)  & ~\V149(1) ;
  assign n501 = ~\V149(0)  & n500;
  assign n502 = ~n499 & ~n501;
  assign n503 = \V169(0)  & ~\V55(0) ;
  assign n504 = ~\V292(0)  & n503;
  assign n505 = ~\V291(0)  & n504;
  assign n506 = ~\V802(0)  & n505;
  assign n507 = n496 & n506;
  assign n508 = ~n490 & n507;
  assign n509 = ~\V292(0)  & \V169(0) ;
  assign n510 = ~\V291(0)  & n509;
  assign n511 = ~n490 & n510;
  assign n512 = ~n502 & n511;
  assign V763 = n508 | n512;
  assign n514 = \V70(0)  & V763;
  assign n515 = \V165(2)  & \V165(0) ;
  assign n516 = \V165(4)  & n515;
  assign n517 = \V165(5)  & n516;
  assign n518 = \V165(6)  & n517;
  assign n519 = \V165(7)  & n518;
  assign n520 = \V165(1)  & n519;
  assign n521 = \V165(3)  & n520;
  assign n522 = \V261(0)  & n521;
  assign n523 = n514 & n522;
  assign n524 = ~\V204(0)  & n521;
  assign n525 = \V261(0)  & n524;
  assign n526 = ~n523 & ~n525;
  assign n527 = ~\V262(0)  & n526;
  assign n528 = \V149(5)  & ~\V149(4) ;
  assign n529 = ~\V174(0)  & n501;
  assign V707 = ~\V149(3)  & n529;
  assign n531 = ~\V149(5)  & ~\V149(4) ;
  assign n532 = \V88(2)  & \V88(3) ;
  assign n533 = V707 & n532;
  assign n534 = n528 & n533;
  assign n535 = ~\V88(2)  & ~\V88(3) ;
  assign n536 = V707 & n535;
  assign n537 = n531 & n536;
  assign n538 = ~n534 & ~n537;
  assign n539 = V707 & n538;
  assign n540 = ~\V149(1)  & n482;
  assign n541 = ~n501 & ~n540;
  assign n542 = \V169(1)  & ~n541;
  assign n543 = n539 & n542;
  assign n544 = ~\V56(0)  & ~\V60(0) ;
  assign n545 = \V149(3)  & n529;
  assign n546 = ~n543 & ~n545;
  assign n547 = ~\V174(0)  & n499;
  assign n548 = \V278(0)  & ~n547;
  assign n549 = ~\V277(0)  & \V278(0) ;
  assign n550 = ~n548 & ~n549;
  assign n551 = \V149(3)  & n540;
  assign n552 = n540 & ~n551;
  assign n553 = ~n491 & n552;
  assign n554 = ~n551 & ~n553;
  assign n555 = n547 & n550;
  assign n556 = n554 & ~n555;
  assign n557 = ~n542 & n545;
  assign n558 = \V149(7)  & n495;
  assign n559 = ~\V149(5)  & \V149(4) ;
  assign n560 = n558 & n559;
  assign n561 = ~\V56(0)  & \V53(0) ;
  assign n562 = n527 & n561;
  assign n563 = ~n486 & n562;
  assign n564 = ~n485 & n563;
  assign n565 = \V57(0)  & ~n543;
  assign n566 = n539 & n565;
  assign n567 = \V53(0)  & ~n543;
  assign n568 = n539 & n567;
  assign n569 = \V56(0)  & ~n543;
  assign n570 = n539 & n569;
  assign n571 = \V57(0)  & ~n546;
  assign n572 = n544 & n571;
  assign n573 = \V53(0)  & ~n546;
  assign n574 = n544 & n573;
  assign n575 = \V57(0)  & ~n556;
  assign n576 = \V53(0)  & ~n556;
  assign n577 = \V56(0)  & ~n556;
  assign n578 = \V57(0)  & n557;
  assign n579 = \V53(0)  & n557;
  assign n580 = \V56(0)  & n557;
  assign n581 = ~n560 & ~n580;
  assign n582 = ~n579 & n581;
  assign n583 = ~n578 & n582;
  assign n584 = ~n577 & n583;
  assign n585 = ~n576 & n584;
  assign n586 = ~n575 & n585;
  assign n587 = ~n574 & n586;
  assign n588 = ~n572 & n587;
  assign n589 = ~n570 & n588;
  assign n590 = ~n568 & n589;
  assign n591 = ~n566 & n590;
  assign n592 = ~n564 & n591;
  assign n593 = V763 & n527;
  assign n594 = n592 & ~n593;
  assign n595 = ~\V59(0)  & n486;
  assign n596 = n550 & n595;
  assign n597 = n594 & ~n596;
  assign n598 = ~n486 & ~n547;
  assign n599 = ~n596 & ~n598;
  assign n600 = \V60(0)  & ~n598;
  assign n601 = ~\V174(0)  & n485;
  assign n602 = ~\V174(0)  & ~n541;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n600 & n603;
  assign n605 = ~n599 & n604;
  assign n606 = ~n527 & n605;
  assign n607 = n597 & n606;
  assign n608 = n592 & n593;
  assign n609 = V763 & ~n544;
  assign n610 = \V59(0)  & V763;
  assign n611 = ~n609 & ~n610;
  assign n612 = n608 & n611;
  assign n613 = n608 & ~n611;
  assign n614 = n527 & ~n605;
  assign n615 = n597 & n614;
  assign n616 = n541 & n615;
  assign n617 = ~n541 & n615;
  assign n618 = \V60(0)  & n547;
  assign n619 = \V60(0)  & n551;
  assign n620 = ~n592 & ~n619;
  assign n621 = ~n618 & n620;
  assign n622 = \V257(5)  & n607;
  assign n623 = \V32(3)  & n612;
  assign n624 = \V32(0)  & n613;
  assign n625 = \V189(4)  & n616;
  assign n626 = \V229(4)  & n617;
  assign n627 = \V32(10)  & n621;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~n625 & n628;
  assign n630 = ~n624 & n629;
  assign n631 = ~n623 & n630;
  assign \V1213(10)  = n622 | ~n631;
  assign n633 = \V257(6)  & n607;
  assign n634 = \V32(4)  & n612;
  assign n635 = \V32(1)  & n613;
  assign n636 = \V189(5)  & n616;
  assign n637 = \V229(5)  & n617;
  assign n638 = \V32(11)  & n621;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n636 & n639;
  assign n641 = ~n635 & n640;
  assign n642 = ~n634 & n641;
  assign \V1213(11)  = n633 | ~n642;
  assign \V1440(0)  = ~\V14(0)  | ~n550;
  assign n645 = \V207(0)  & ~\V172(0) ;
  assign n646 = \V207(0)  & ~\V56(0) ;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~\V149(7)  & n647;
  assign n649 = n540 & ~n648;
  assign n650 = \V56(0)  & ~n598;
  assign n651 = ~n485 & n598;
  assign n652 = ~\V241(0)  & ~n485;
  assign n653 = ~n651 & ~n652;
  assign n654 = \V261(0)  & n653;
  assign n655 = \V149(7)  & ~\V174(0) ;
  assign n656 = n496 & n655;
  assign n657 = ~n542 & ~n656;
  assign n658 = ~\V149(6)  & n494;
  assign n659 = ~\V149(7)  & n658;
  assign n660 = n528 & n659;
  assign n661 = n657 & ~n660;
  assign n662 = \V59(0)  & ~n657;
  assign n663 = ~n661 & ~n662;
  assign n664 = \V67(0)  & \V215(0) ;
  assign n665 = \V172(0)  & n664;
  assign n666 = ~n540 & ~n647;
  assign n667 = ~n663 & n666;
  assign n668 = ~\V214(0)  & ~n665;
  assign n669 = \V62(0)  & ~n647;
  assign n670 = n660 & n669;
  assign n671 = n668 & ~n670;
  assign n672 = ~n667 & n671;
  assign n673 = ~\V275(0)  & \V242(0) ;
  assign n674 = \V134(1)  & n673;
  assign n675 = \V134(0)  & n674;
  assign n676 = \V272(0)  & n675;
  assign n677 = ~\V802(0)  & n676;
  assign n678 = ~n550 & n677;
  assign n679 = \V242(0)  & ~\V802(0) ;
  assign n680 = n550 & n679;
  assign n681 = ~n651 & n680;
  assign n682 = ~n650 & n681;
  assign n683 = ~\V275(0)  & \V272(0) ;
  assign n684 = ~\V802(0)  & n683;
  assign n685 = n654 & n684;
  assign n686 = ~\V802(0)  & n550;
  assign n687 = n654 & n686;
  assign n688 = n672 & ~n687;
  assign n689 = ~n685 & n688;
  assign n690 = ~n682 & n689;
  assign n691 = ~n678 & n690;
  assign n692 = n540 & ~n647;
  assign n693 = ~\V56(0)  & n647;
  assign n694 = n649 & ~n693;
  assign n695 = ~\V149(3)  & n540;
  assign n696 = n491 & n695;
  assign n697 = ~n538 & ~n542;
  assign n698 = ~n696 & ~n697;
  assign n699 = \V56(0)  & ~n698;
  assign n700 = ~\V248(0)  & \V177(0) ;
  assign n701 = ~\V172(0)  & n700;
  assign n702 = n651 & n701;
  assign n703 = n541 & n702;
  assign n704 = n691 & n703;
  assign n705 = ~n649 & n704;
  assign n706 = ~\V248(0)  & ~\V278(0) ;
  assign n707 = \V177(0)  & n706;
  assign n708 = ~\V172(0)  & n707;
  assign n709 = n541 & n708;
  assign n710 = n691 & n709;
  assign n711 = ~n649 & n710;
  assign n712 = ~\V171(0)  & n701;
  assign n713 = n651 & n712;
  assign n714 = n691 & n713;
  assign n715 = ~n649 & n714;
  assign n716 = ~\V171(0)  & n708;
  assign n717 = n691 & n716;
  assign n718 = ~n649 & n717;
  assign n719 = ~\V248(0)  & ~\V56(0) ;
  assign n720 = \V177(0)  & n719;
  assign n721 = n651 & n720;
  assign n722 = n691 & n721;
  assign n723 = ~n692 & n722;
  assign n724 = ~\V278(0)  & n719;
  assign n725 = \V177(0)  & n724;
  assign n726 = n691 & n725;
  assign n727 = ~n692 & n726;
  assign n728 = \V59(0)  & ~n538;
  assign n729 = n542 & n728;
  assign n730 = n691 & n729;
  assign n731 = ~n694 & n730;
  assign n732 = ~\V271(0)  & ~\V274(0) ;
  assign n733 = n691 & n732;
  assign n734 = ~n694 & n733;
  assign n735 = ~\V172(0)  & n691;
  assign n736 = ~n649 & n735;
  assign n737 = n699 & n736;
  assign n738 = ~n734 & ~n737;
  assign n739 = ~n731 & n738;
  assign n740 = ~n727 & n739;
  assign n741 = ~n723 & n740;
  assign n742 = ~n718 & n741;
  assign n743 = ~n715 & n742;
  assign n744 = ~n711 & n743;
  assign \V1536(0)  = ~n705 & n744;
  assign n746 = n527 & n605;
  assign n747 = n596 & n746;
  assign n748 = \V149(4)  & n747;
  assign n749 = \V257(7)  & n607;
  assign n750 = \V32(5)  & n612;
  assign n751 = \V32(2)  & n613;
  assign n752 = \V194(0)  & n616;
  assign n753 = \V234(0)  & n617;
  assign n754 = \V78(4)  & n621;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n752 & n755;
  assign n757 = ~n751 & n756;
  assign n758 = ~n750 & n757;
  assign n759 = ~n749 & n758;
  assign \V321(2)  = ~n748 & n759;
  assign n761 = \V84(4)  & ~\V84(5) ;
  assign n762 = ~\V84(4)  & \V84(5) ;
  assign n763 = ~n761 & ~n762;
  assign n764 = \V84(3)  & ~n763;
  assign n765 = ~\V84(3)  & n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = \V84(2)  & ~n766;
  assign n768 = ~\V84(2)  & n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~\V94(1)  & ~n769;
  assign n771 = \V94(1)  & n769;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~\V88(2)  & \V88(3) ;
  assign n774 = \V88(2)  & ~\V88(3) ;
  assign n775 = ~n773 & ~n774;
  assign n776 = \V88(1)  & ~n775;
  assign n777 = ~\V88(1)  & n775;
  assign n778 = ~n776 & ~n777;
  assign n779 = \V88(0)  & ~n778;
  assign n780 = ~\V88(0)  & n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = \V149(7)  & n658;
  assign n783 = n528 & n782;
  assign n784 = ~\V149(7)  & n495;
  assign n785 = n559 & n784;
  assign n786 = ~\V78(2)  & \V78(3) ;
  assign n787 = \V78(2)  & ~\V78(3) ;
  assign n788 = ~n786 & ~n787;
  assign n789 = \V78(1)  & ~n788;
  assign n790 = ~\V78(1)  & n788;
  assign n791 = ~n789 & ~n790;
  assign n792 = \V78(0)  & ~n791;
  assign n793 = ~\V78(0)  & n791;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~\V94(0)  & ~n794;
  assign n796 = \V94(0)  & n794;
  assign n797 = ~n795 & ~n796;
  assign n798 = \V84(0)  & ~\V84(1) ;
  assign n799 = ~\V84(0)  & \V84(1) ;
  assign n800 = ~n798 & ~n799;
  assign n801 = \V78(5)  & ~n800;
  assign n802 = ~\V78(5)  & n800;
  assign n803 = ~n801 & ~n802;
  assign n804 = \V78(4)  & ~n803;
  assign n805 = ~\V78(4)  & n803;
  assign n806 = ~n804 & ~n805;
  assign n807 = \V802(0)  & n547;
  assign n808 = \V802(0)  & n529;
  assign n809 = \V802(0)  & n540;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n807 & n810;
  assign n812 = \V56(0)  & n560;
  assign n813 = n781 & n812;
  assign n814 = n772 & n813;
  assign n815 = \V56(0)  & n783;
  assign n816 = n781 & n815;
  assign n817 = n772 & n816;
  assign n818 = \V56(0)  & n785;
  assign n819 = n781 & n818;
  assign n820 = n772 & n819;
  assign n821 = ~n781 & n812;
  assign n822 = ~n772 & n821;
  assign n823 = ~n781 & n815;
  assign n824 = ~n772 & n823;
  assign n825 = ~n781 & n818;
  assign n826 = ~n772 & n825;
  assign n827 = n806 & n812;
  assign n828 = n797 & n827;
  assign n829 = n806 & n815;
  assign n830 = n797 & n829;
  assign n831 = n806 & n818;
  assign n832 = n797 & n831;
  assign n833 = ~n806 & n812;
  assign n834 = ~n797 & n833;
  assign n835 = ~n806 & n815;
  assign n836 = ~n797 & n835;
  assign n837 = ~n806 & n818;
  assign n838 = ~n797 & n837;
  assign n839 = n772 & n781;
  assign n840 = ~n811 & n839;
  assign n841 = ~n772 & ~n781;
  assign n842 = ~n811 & n841;
  assign n843 = n797 & n806;
  assign n844 = ~n811 & n843;
  assign n845 = ~n797 & ~n806;
  assign n846 = ~n811 & n845;
  assign n847 = ~n844 & ~n846;
  assign n848 = ~n842 & n847;
  assign n849 = ~n840 & n848;
  assign n850 = ~n838 & n849;
  assign n851 = ~n836 & n850;
  assign n852 = ~n834 & n851;
  assign n853 = ~n832 & n852;
  assign n854 = ~n830 & n853;
  assign n855 = ~n828 & n854;
  assign n856 = ~n826 & n855;
  assign n857 = ~n824 & n856;
  assign n858 = ~n822 & n857;
  assign n859 = ~n820 & n858;
  assign n860 = ~n817 & n859;
  assign n861 = ~n814 & n860;
  assign n862 = \V15(0)  & ~n540;
  assign n863 = \V15(0)  & \V802(0) ;
  assign n864 = n861 & ~n863;
  assign \V1480(0)  = n862 | ~n864;
  assign n866 = ~\V165(2)  & \V165(0) ;
  assign n867 = \V165(1)  & n866;
  assign n868 = ~n647 & ~n867;
  assign n869 = \V290(0)  & n867;
  assign n870 = ~n540 & ~n663;
  assign n871 = n868 & n870;
  assign n872 = ~n670 & ~n869;
  assign \V1741(0)  = n871 | ~n872;
  assign n874 = \V802(0)  & ~n651;
  assign V587 = ~\V243(0)  & ~n874;
  assign n876 = \V243(0)  & \V244(0) ;
  assign n877 = ~\V245(0)  & n876;
  assign n878 = ~n874 & n877;
  assign n879 = \V245(0)  & ~\V244(0) ;
  assign n880 = ~n874 & n879;
  assign n881 = \V245(0)  & V587;
  assign n882 = ~n880 & ~n881;
  assign \V597(0)  = n878 | ~n882;
  assign n884 = ~\V246(0)  & \V245(0) ;
  assign n885 = ~\V597(0)  & n884;
  assign n886 = ~n874 & n885;
  assign n887 = \V246(0)  & \V597(0) ;
  assign n888 = \V246(0)  & ~\V245(0) ;
  assign n889 = ~n874 & n888;
  assign n890 = ~n887 & ~n889;
  assign \V603(0)  = n886 | ~n890;
  assign n892 = ~n560 & ~\V1213(11) ;
  assign n893 = ~\V78(3)  & n560;
  assign \V1781(1)  = n892 | n893;
  assign n895 = ~n560 & ~\V1213(10) ;
  assign n896 = ~\V78(2)  & n560;
  assign \V1781(0)  = n895 | n896;
  assign n898 = \V199(3)  & \V199(4) ;
  assign n899 = \V199(2)  & n898;
  assign n900 = \V199(1)  & \V199(0) ;
  assign n901 = n899 & n900;
  assign n902 = \V194(4)  & n901;
  assign n903 = \V194(3)  & n902;
  assign n904 = \V194(2)  & \V194(1) ;
  assign n905 = n903 & n904;
  assign n906 = \V194(0)  & n905;
  assign n907 = \V14(0)  & \V242(0) ;
  assign n908 = n598 & n907;
  assign n909 = ~n651 & ~\V1536(0) ;
  assign n910 = n906 & n909;
  assign \V1726(0)  = n908 | n910;
  assign n912 = \V183(1)  & n616;
  assign n913 = \V223(1)  & n617;
  assign n914 = \V32(1)  & n621;
  assign n915 = ~n913 & ~n914;
  assign \V1213(1)  = n912 | ~n915;
  assign n917 = ~\V149(7)  & n531;
  assign n918 = \V149(3)  & n493;
  assign n919 = ~\V149(6)  & n918;
  assign n920 = n917 & n919;
  assign n921 = ~\V802(0)  & n920;
  assign n922 = \V1213(1)  & ~n921;
  assign n923 = \V183(3)  & n616;
  assign n924 = \V223(3)  & n617;
  assign n925 = \V32(3)  & n621;
  assign n926 = ~n924 & ~n925;
  assign \V1213(3)  = n923 | ~n926;
  assign n928 = \V288(7)  & ~\V288(6) ;
  assign n929 = \V288(5)  & ~\V288(4) ;
  assign n930 = ~n928 & ~n929;
  assign n931 = n928 & n929;
  assign n932 = ~n930 & ~n931;
  assign n933 = \V288(3)  & ~\V288(2) ;
  assign n934 = ~n932 & ~n933;
  assign n935 = n932 & n933;
  assign n936 = ~n934 & ~n935;
  assign n937 = \V288(1)  & ~\V288(0) ;
  assign n938 = ~n936 & ~n937;
  assign n939 = n936 & n937;
  assign n940 = ~n938 & ~n939;
  assign n941 = \V1213(3)  & n940;
  assign n942 = ~\V1213(3)  & ~n940;
  assign n943 = ~n941 & ~n942;
  assign n944 = \V183(2)  & n616;
  assign n945 = \V223(2)  & n617;
  assign n946 = \V32(2)  & n621;
  assign n947 = ~n945 & ~n946;
  assign \V1213(2)  = n944 | ~n947;
  assign n949 = \V183(0)  & n616;
  assign n950 = \V223(0)  & n617;
  assign n951 = \V32(0)  & n621;
  assign n952 = ~n950 & ~n951;
  assign \V1213(0)  = n949 | ~n952;
  assign n954 = ~\V288(1)  & \V288(0) ;
  assign n955 = ~n936 & n937;
  assign n956 = ~n932 & n933;
  assign n957 = ~\V288(7)  & \V288(6) ;
  assign n958 = ~n928 & ~n957;
  assign n959 = ~\V288(5)  & \V288(4) ;
  assign n960 = ~n958 & n959;
  assign n961 = n958 & ~n959;
  assign n962 = ~n960 & ~n961;
  assign n963 = ~n929 & ~n962;
  assign n964 = n929 & n932;
  assign n965 = n962 & n964;
  assign n966 = ~n963 & ~n965;
  assign n967 = ~\V288(3)  & \V288(2) ;
  assign n968 = ~n966 & ~n967;
  assign n969 = n966 & n967;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n956 & ~n970;
  assign n972 = n956 & n970;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n954 & ~n973;
  assign n975 = n954 & n973;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n955 & ~n976;
  assign n978 = n955 & n976;
  assign n979 = ~n977 & ~n978;
  assign n980 = n954 & ~n979;
  assign n981 = ~n954 & n979;
  assign n982 = ~n980 & ~n981;
  assign n983 = n940 & n982;
  assign n984 = ~n937 & ~n940;
  assign n985 = ~n982 & n984;
  assign n986 = n937 & ~n979;
  assign n987 = ~n983 & ~n986;
  assign n988 = ~n985 & n987;
  assign n989 = n940 & n979;
  assign n990 = ~n940 & ~n979;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n940 & n991;
  assign n993 = \V288(1)  & \V288(0) ;
  assign n994 = \V288(3)  & \V288(2) ;
  assign n995 = ~\V288(7)  & ~\V288(6) ;
  assign n996 = \V288(5)  & \V288(4) ;
  assign n997 = ~n995 & n996;
  assign n998 = n995 & ~n996;
  assign n999 = ~n997 & ~n998;
  assign n1000 = n959 & n962;
  assign n1001 = n929 & ~n962;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~n999 & n1002;
  assign n1004 = n999 & ~n1002;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~n994 & ~n1005;
  assign n1007 = n994 & n1005;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n966 & n973;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = n1008 & n1009;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n993 & ~n1012;
  assign n1014 = n993 & n1012;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = ~n973 & n979;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = n1015 & n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = ~n989 & ~n1019;
  assign n1021 = n989 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = n992 & n1022;
  assign n1024 = ~n954 & ~n1022;
  assign n1025 = ~n992 & n1024;
  assign n1026 = ~n954 & n1023;
  assign n1027 = n954 & ~n1019;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1025 & n1028;
  assign n1030 = n983 & n1029;
  assign n1031 = ~n937 & ~n1029;
  assign n1032 = ~n983 & n1031;
  assign n1033 = ~n937 & n1030;
  assign n1034 = n937 & ~n1019;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = ~n1032 & n1035;
  assign n1037 = n1019 & ~n1022;
  assign n1038 = n995 & ~n1005;
  assign n1039 = n1008 & ~n1038;
  assign n1040 = n994 & n1039;
  assign n1041 = ~n1012 & n1038;
  assign n1042 = n1009 & ~n1038;
  assign n1043 = ~n1008 & n1042;
  assign n1044 = ~n1041 & ~n1043;
  assign n1045 = ~n1040 & n1044;
  assign n1046 = n1015 & n1045;
  assign n1047 = n993 & n1046;
  assign n1048 = n1015 & ~n1045;
  assign n1049 = ~n993 & n1048;
  assign n1050 = ~n1019 & ~n1045;
  assign n1051 = n1016 & n1045;
  assign n1052 = ~n1015 & n1051;
  assign n1053 = ~n1050 & ~n1052;
  assign n1054 = ~n1049 & n1053;
  assign n1055 = ~n1047 & n1054;
  assign n1056 = ~n1037 & ~n1055;
  assign n1057 = ~n1023 & n1056;
  assign n1058 = n954 & ~n1055;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = n937 & ~n1055;
  assign n1061 = ~n937 & ~n1059;
  assign n1062 = ~n1030 & n1061;
  assign n1063 = ~n1060 & ~n1062;
  assign n1064 = ~\V1213(1)  & ~n921;
  assign n1065 = n922 & ~\V1213(0) ;
  assign n1066 = ~\V1213(0)  & n1064;
  assign n1067 = n991 & ~n1022;
  assign n1068 = \V1213(0)  & n1067;
  assign n1069 = ~\V1213(2)  & n1068;
  assign n1070 = n1056 & n1069;
  assign n1071 = ~n943 & n1070;
  assign n1072 = n922 & n1071;
  assign n1073 = n993 & n1072;
  assign n1074 = ~n991 & ~n1022;
  assign n1075 = \V1213(0)  & n1074;
  assign n1076 = \V1213(2)  & n1075;
  assign n1077 = n1056 & n1076;
  assign n1078 = ~n943 & n1077;
  assign n1079 = n922 & n1078;
  assign n1080 = n993 & n1079;
  assign n1081 = n991 & n1022;
  assign n1082 = \V1213(0)  & n1081;
  assign n1083 = ~\V1213(2)  & n1082;
  assign n1084 = n1056 & n1083;
  assign n1085 = ~n943 & n1084;
  assign n1086 = n1064 & n1085;
  assign n1087 = n993 & n1086;
  assign n1088 = ~n991 & n1022;
  assign n1089 = \V1213(0)  & n1088;
  assign n1090 = \V1213(2)  & n1089;
  assign n1091 = n1056 & n1090;
  assign n1092 = ~n943 & n1091;
  assign n1093 = n1064 & n1092;
  assign n1094 = n993 & n1093;
  assign n1095 = ~\V1213(2)  & n1067;
  assign n1096 = ~n1056 & n1095;
  assign n1097 = ~n943 & n1096;
  assign n1098 = n993 & n1097;
  assign n1099 = n1065 & n1098;
  assign n1100 = \V1213(2)  & n1074;
  assign n1101 = ~n1056 & n1100;
  assign n1102 = ~n943 & n1101;
  assign n1103 = n993 & n1102;
  assign n1104 = n1065 & n1103;
  assign n1105 = ~\V1213(2)  & n1081;
  assign n1106 = ~n1056 & n1105;
  assign n1107 = ~n943 & n1106;
  assign n1108 = n993 & n1107;
  assign n1109 = n1066 & n1108;
  assign n1110 = \V1213(2)  & n1088;
  assign n1111 = ~n1056 & n1110;
  assign n1112 = ~n943 & n1111;
  assign n1113 = n993 & n1112;
  assign n1114 = n1066 & n1113;
  assign n1115 = ~n1109 & ~n1114;
  assign n1116 = ~n1104 & n1115;
  assign n1117 = ~n1099 & n1116;
  assign n1118 = ~n1094 & n1117;
  assign n1119 = ~n1087 & n1118;
  assign n1120 = ~n1080 & n1119;
  assign n1121 = ~n1073 & n1120;
  assign n1122 = n937 & n1063;
  assign n1123 = ~n1036 & n1122;
  assign n1124 = n988 & n1123;
  assign n1125 = ~\V1213(0)  & n1124;
  assign n1126 = ~\V1213(2)  & n1125;
  assign n1127 = n943 & n1126;
  assign n1128 = n922 & n1127;
  assign n1129 = n937 & ~n1063;
  assign n1130 = ~n1036 & n1129;
  assign n1131 = n988 & n1130;
  assign n1132 = \V1213(0)  & n1131;
  assign n1133 = ~\V1213(2)  & n1132;
  assign n1134 = n943 & n1133;
  assign n1135 = n922 & n1134;
  assign n1136 = ~n988 & n1123;
  assign n1137 = ~\V1213(0)  & n1136;
  assign n1138 = \V1213(2)  & n1137;
  assign n1139 = n943 & n1138;
  assign n1140 = n922 & n1139;
  assign n1141 = ~n988 & n1130;
  assign n1142 = \V1213(0)  & n1141;
  assign n1143 = \V1213(2)  & n1142;
  assign n1144 = n943 & n1143;
  assign n1145 = n922 & n1144;
  assign n1146 = \V288(0)  & n1063;
  assign n1147 = ~n1036 & n1146;
  assign n1148 = n988 & n1147;
  assign n1149 = ~\V1213(0)  & n1148;
  assign n1150 = ~\V1213(2)  & n1149;
  assign n1151 = ~n943 & n1150;
  assign n1152 = n922 & n1151;
  assign n1153 = \V288(0)  & ~n1063;
  assign n1154 = ~n1036 & n1153;
  assign n1155 = n988 & n1154;
  assign n1156 = \V1213(0)  & n1155;
  assign n1157 = ~\V1213(2)  & n1156;
  assign n1158 = ~n943 & n1157;
  assign n1159 = n922 & n1158;
  assign n1160 = ~n988 & n1147;
  assign n1161 = ~\V1213(0)  & n1160;
  assign n1162 = \V1213(2)  & n1161;
  assign n1163 = ~n943 & n1162;
  assign n1164 = n922 & n1163;
  assign n1165 = ~n988 & n1154;
  assign n1166 = \V1213(0)  & n1165;
  assign n1167 = \V1213(2)  & n1166;
  assign n1168 = ~n943 & n1167;
  assign n1169 = n922 & n1168;
  assign n1170 = n1036 & n1122;
  assign n1171 = n988 & n1170;
  assign n1172 = ~\V1213(0)  & n1171;
  assign n1173 = ~\V1213(2)  & n1172;
  assign n1174 = n943 & n1173;
  assign n1175 = n1064 & n1174;
  assign n1176 = n1036 & n1129;
  assign n1177 = n988 & n1176;
  assign n1178 = \V1213(0)  & n1177;
  assign n1179 = ~\V1213(2)  & n1178;
  assign n1180 = n943 & n1179;
  assign n1181 = n1064 & n1180;
  assign n1182 = ~n988 & n1170;
  assign n1183 = ~\V1213(0)  & n1182;
  assign n1184 = \V1213(2)  & n1183;
  assign n1185 = n943 & n1184;
  assign n1186 = n1064 & n1185;
  assign n1187 = ~n988 & n1176;
  assign n1188 = \V1213(0)  & n1187;
  assign n1189 = \V1213(2)  & n1188;
  assign n1190 = n943 & n1189;
  assign n1191 = n1064 & n1190;
  assign n1192 = n1036 & n1146;
  assign n1193 = n988 & n1192;
  assign n1194 = ~\V1213(0)  & n1193;
  assign n1195 = ~\V1213(2)  & n1194;
  assign n1196 = ~n943 & n1195;
  assign n1197 = n1064 & n1196;
  assign n1198 = n1036 & n1153;
  assign n1199 = n988 & n1198;
  assign n1200 = \V1213(0)  & n1199;
  assign n1201 = ~\V1213(2)  & n1200;
  assign n1202 = ~n943 & n1201;
  assign n1203 = n1064 & n1202;
  assign n1204 = ~n988 & n1192;
  assign n1205 = ~\V1213(0)  & n1204;
  assign n1206 = \V1213(2)  & n1205;
  assign n1207 = ~n943 & n1206;
  assign n1208 = n1064 & n1207;
  assign n1209 = ~n988 & n1198;
  assign n1210 = \V1213(0)  & n1209;
  assign n1211 = \V1213(2)  & n1210;
  assign n1212 = ~n943 & n1211;
  assign n1213 = n1064 & n1212;
  assign n1214 = n1121 & ~n1213;
  assign n1215 = ~n1208 & n1214;
  assign n1216 = ~n1203 & n1215;
  assign n1217 = ~n1197 & n1216;
  assign n1218 = ~n1191 & n1217;
  assign n1219 = ~n1186 & n1218;
  assign n1220 = ~n1181 & n1219;
  assign n1221 = ~n1175 & n1220;
  assign n1222 = ~n1169 & n1221;
  assign n1223 = ~n1164 & n1222;
  assign n1224 = ~n1159 & n1223;
  assign n1225 = ~n1152 & n1224;
  assign n1226 = ~n1145 & n1225;
  assign n1227 = ~n1140 & n1226;
  assign n1228 = ~n1135 & n1227;
  assign n1229 = ~n1128 & n1228;
  assign n1230 = n527 & n1229;
  assign n1231 = \V1213(3)  & n936;
  assign n1232 = ~\V1213(3)  & ~n936;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = n967 & ~n973;
  assign n1235 = ~n967 & n973;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = n936 & n1236;
  assign n1238 = ~n933 & ~n936;
  assign n1239 = ~n1236 & n1238;
  assign n1240 = n933 & ~n973;
  assign n1241 = ~n1237 & ~n1240;
  assign n1242 = ~n1239 & n1241;
  assign n1243 = ~n967 & n1012;
  assign n1244 = ~n1236 & n1243;
  assign n1245 = ~n973 & ~n1012;
  assign n1246 = ~n1012 & n1236;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1244 & n1247;
  assign n1249 = n933 & ~n1012;
  assign n1250 = ~n933 & ~n1248;
  assign n1251 = ~n1237 & n1250;
  assign n1252 = ~n1249 & ~n1251;
  assign n1253 = n936 & n973;
  assign n1254 = ~n1012 & ~n1253;
  assign n1255 = n1012 & n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n936 & n973;
  assign n1258 = n1256 & n1257;
  assign n1259 = ~n1045 & n1256;
  assign n1260 = ~n1258 & n1259;
  assign n1261 = n967 & ~n1045;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~n933 & ~n1262;
  assign n1264 = n933 & ~n1045;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = \V1213(2)  & n973;
  assign n1267 = ~\V1213(2)  & ~n973;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~n936 & \V1213(0) ;
  assign n1270 = ~\V1213(3)  & n1269;
  assign n1271 = ~n1256 & n1270;
  assign n1272 = n1259 & n1271;
  assign n1273 = n1268 & n1272;
  assign n1274 = n922 & n1273;
  assign n1275 = n994 & n1274;
  assign n1276 = n936 & \V1213(0) ;
  assign n1277 = \V1213(3)  & n1276;
  assign n1278 = ~n1256 & n1277;
  assign n1279 = n1259 & n1278;
  assign n1280 = ~n1268 & n1279;
  assign n1281 = n922 & n1280;
  assign n1282 = n994 & n1281;
  assign n1283 = n1256 & n1270;
  assign n1284 = n1259 & n1283;
  assign n1285 = n1268 & n1284;
  assign n1286 = n1064 & n1285;
  assign n1287 = n994 & n1286;
  assign n1288 = n1256 & n1277;
  assign n1289 = n1259 & n1288;
  assign n1290 = ~n1268 & n1289;
  assign n1291 = n1064 & n1290;
  assign n1292 = n994 & n1291;
  assign n1293 = n1232 & ~n1256;
  assign n1294 = ~n1259 & n1293;
  assign n1295 = n1268 & n1294;
  assign n1296 = n994 & n1295;
  assign n1297 = n1065 & n1296;
  assign n1298 = n1231 & ~n1256;
  assign n1299 = ~n1259 & n1298;
  assign n1300 = ~n1268 & n1299;
  assign n1301 = n994 & n1300;
  assign n1302 = n1065 & n1301;
  assign n1303 = n1232 & n1256;
  assign n1304 = ~n1259 & n1303;
  assign n1305 = n1268 & n1304;
  assign n1306 = n994 & n1305;
  assign n1307 = n1066 & n1306;
  assign n1308 = n1231 & n1256;
  assign n1309 = ~n1259 & n1308;
  assign n1310 = ~n1268 & n1309;
  assign n1311 = n994 & n1310;
  assign n1312 = n1066 & n1311;
  assign n1313 = ~n1307 & ~n1312;
  assign n1314 = ~n1302 & n1313;
  assign n1315 = ~n1297 & n1314;
  assign n1316 = ~n1292 & n1315;
  assign n1317 = ~n1287 & n1316;
  assign n1318 = ~n1282 & n1317;
  assign n1319 = ~n1275 & n1318;
  assign n1320 = ~\V1213(2)  & ~\V1213(0) ;
  assign n1321 = n933 & n1320;
  assign n1322 = n1265 & n1321;
  assign n1323 = ~n1252 & n1322;
  assign n1324 = n1242 & n1323;
  assign n1325 = n1233 & n1324;
  assign n1326 = n922 & n1325;
  assign n1327 = ~\V1213(2)  & \V1213(0) ;
  assign n1328 = n933 & n1327;
  assign n1329 = ~n1265 & n1328;
  assign n1330 = ~n1252 & n1329;
  assign n1331 = n1242 & n1330;
  assign n1332 = n1233 & n1331;
  assign n1333 = n922 & n1332;
  assign n1334 = \V1213(2)  & ~\V1213(0) ;
  assign n1335 = n933 & n1334;
  assign n1336 = n1265 & n1335;
  assign n1337 = ~n1252 & n1336;
  assign n1338 = ~n1242 & n1337;
  assign n1339 = n1233 & n1338;
  assign n1340 = n922 & n1339;
  assign n1341 = \V1213(2)  & \V1213(0) ;
  assign n1342 = n933 & n1341;
  assign n1343 = ~n1265 & n1342;
  assign n1344 = ~n1252 & n1343;
  assign n1345 = ~n1242 & n1344;
  assign n1346 = n1233 & n1345;
  assign n1347 = n922 & n1346;
  assign n1348 = \V288(2)  & ~\V1213(0) ;
  assign n1349 = ~\V1213(2)  & n1348;
  assign n1350 = n1265 & n1349;
  assign n1351 = ~n1252 & n1350;
  assign n1352 = n1242 & n1351;
  assign n1353 = ~n1233 & n1352;
  assign n1354 = n922 & n1353;
  assign n1355 = \V288(2)  & \V1213(0) ;
  assign n1356 = ~\V1213(2)  & n1355;
  assign n1357 = ~n1265 & n1356;
  assign n1358 = ~n1252 & n1357;
  assign n1359 = n1242 & n1358;
  assign n1360 = ~n1233 & n1359;
  assign n1361 = n922 & n1360;
  assign n1362 = \V1213(2)  & n1348;
  assign n1363 = n1265 & n1362;
  assign n1364 = ~n1252 & n1363;
  assign n1365 = ~n1242 & n1364;
  assign n1366 = ~n1233 & n1365;
  assign n1367 = n922 & n1366;
  assign n1368 = \V1213(2)  & n1355;
  assign n1369 = ~n1265 & n1368;
  assign n1370 = ~n1252 & n1369;
  assign n1371 = ~n1242 & n1370;
  assign n1372 = ~n1233 & n1371;
  assign n1373 = n922 & n1372;
  assign n1374 = n1252 & n1322;
  assign n1375 = n1242 & n1374;
  assign n1376 = n1233 & n1375;
  assign n1377 = n1064 & n1376;
  assign n1378 = n1252 & n1329;
  assign n1379 = n1242 & n1378;
  assign n1380 = n1233 & n1379;
  assign n1381 = n1064 & n1380;
  assign n1382 = n1252 & n1336;
  assign n1383 = ~n1242 & n1382;
  assign n1384 = n1233 & n1383;
  assign n1385 = n1064 & n1384;
  assign n1386 = n1252 & n1343;
  assign n1387 = ~n1242 & n1386;
  assign n1388 = n1233 & n1387;
  assign n1389 = n1064 & n1388;
  assign n1390 = n1252 & n1350;
  assign n1391 = n1242 & n1390;
  assign n1392 = ~n1233 & n1391;
  assign n1393 = n1064 & n1392;
  assign n1394 = n1252 & n1357;
  assign n1395 = n1242 & n1394;
  assign n1396 = ~n1233 & n1395;
  assign n1397 = n1064 & n1396;
  assign n1398 = n1252 & n1363;
  assign n1399 = ~n1242 & n1398;
  assign n1400 = ~n1233 & n1399;
  assign n1401 = n1064 & n1400;
  assign n1402 = n1252 & n1369;
  assign n1403 = ~n1242 & n1402;
  assign n1404 = ~n1233 & n1403;
  assign n1405 = n1064 & n1404;
  assign n1406 = n1319 & ~n1405;
  assign n1407 = ~n1401 & n1406;
  assign n1408 = ~n1397 & n1407;
  assign n1409 = ~n1393 & n1408;
  assign n1410 = ~n1389 & n1409;
  assign n1411 = ~n1385 & n1410;
  assign n1412 = ~n1381 & n1411;
  assign n1413 = ~n1377 & n1412;
  assign n1414 = ~n1373 & n1413;
  assign n1415 = ~n1367 & n1414;
  assign n1416 = ~n1361 & n1415;
  assign n1417 = ~n1354 & n1416;
  assign n1418 = ~n1347 & n1417;
  assign n1419 = ~n1340 & n1418;
  assign n1420 = ~n1333 & n1419;
  assign n1421 = ~n1326 & n1420;
  assign n1422 = ~\V1213(3)  & ~n932;
  assign n1423 = \V1213(3)  & n932;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n959 & n966;
  assign n1426 = n959 & ~n966;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = n932 & n1427;
  assign n1429 = ~n929 & ~n932;
  assign n1430 = ~n1427 & n1429;
  assign n1431 = ~n1428 & ~n1430;
  assign n1432 = ~n1005 & ~n1425;
  assign n1433 = n1005 & n1425;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n929 & ~n1434;
  assign n1436 = n929 & ~n1005;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = \V1213(2)  & ~n966;
  assign n1439 = ~\V1213(2)  & n966;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n932 & ~n1005;
  assign n1442 = n932 & n1005;
  assign n1443 = ~n1441 & ~n1442;
  assign n1444 = n1422 & n1443;
  assign n1445 = ~n1440 & n1444;
  assign n1446 = n996 & n1445;
  assign n1447 = n1066 & n1446;
  assign n1448 = ~\V1213(3)  & ~n1443;
  assign n1449 = ~n1440 & n1448;
  assign n1450 = n996 & n1449;
  assign n1451 = n1065 & n1450;
  assign n1452 = n1423 & n1440;
  assign n1453 = n996 & n1452;
  assign n1454 = n1066 & n1453;
  assign n1455 = ~n1451 & ~n1454;
  assign n1456 = ~n1447 & n1455;
  assign n1457 = n929 & ~\V1213(2) ;
  assign n1458 = n1437 & n1457;
  assign n1459 = n1431 & n1458;
  assign n1460 = n1424 & n1459;
  assign n1461 = n1066 & n1460;
  assign n1462 = \V288(4)  & ~\V1213(2) ;
  assign n1463 = n1437 & n1462;
  assign n1464 = n1431 & n1463;
  assign n1465 = ~n1424 & n1464;
  assign n1466 = n1066 & n1465;
  assign n1467 = ~n1437 & n1457;
  assign n1468 = n1424 & n1467;
  assign n1469 = n1065 & n1468;
  assign n1470 = ~n1437 & n1462;
  assign n1471 = ~n1424 & n1470;
  assign n1472 = n1065 & n1471;
  assign n1473 = n929 & \V1213(2) ;
  assign n1474 = ~n1431 & n1473;
  assign n1475 = n1424 & n1474;
  assign n1476 = n1066 & n1475;
  assign n1477 = \V288(4)  & \V1213(2) ;
  assign n1478 = ~n1431 & n1477;
  assign n1479 = ~n1424 & n1478;
  assign n1480 = n1066 & n1479;
  assign n1481 = n1456 & ~n1480;
  assign n1482 = ~n1476 & n1481;
  assign n1483 = ~n1472 & n1482;
  assign n1484 = ~n1469 & n1483;
  assign n1485 = ~n1466 & n1484;
  assign n1486 = ~n1461 & n1485;
  assign n1487 = \V288(6)  & n1066;
  assign n1488 = \V288(7)  & \V1213(2) ;
  assign n1489 = n1487 & n1488;
  assign n1490 = ~n921 & \V1213(2) ;
  assign n1491 = ~n1489 & n1490;
  assign n1492 = n1486 & n1491;
  assign n1493 = n1421 & n1492;
  assign n1494 = n1230 & n1493;
  assign n1495 = ~n921 & n1486;
  assign n1496 = n1421 & n1495;
  assign n1497 = n1230 & n1496;
  assign n1498 = n995 & n1497;
  assign n1499 = ~n921 & \V1213(3) ;
  assign n1500 = n1486 & n1499;
  assign n1501 = n1421 & n1500;
  assign n1502 = n1230 & n1501;
  assign n1503 = ~n921 & \V1213(0) ;
  assign n1504 = n1486 & n1503;
  assign n1505 = n1421 & n1504;
  assign n1506 = n1230 & n1505;
  assign n1507 = n922 & n1486;
  assign n1508 = n1421 & n1507;
  assign n1509 = n1230 & n1508;
  assign n1510 = ~n1506 & ~n1509;
  assign n1511 = ~n1502 & n1510;
  assign n1512 = ~n1498 & n1511;
  assign V356 = n1494 | ~n1512;
  assign n1514 = n1012 & n1045;
  assign n1515 = n1233 & n1514;
  assign n1516 = n1268 & n1515;
  assign n1517 = n994 & n1516;
  assign n1518 = n1066 & n1517;
  assign n1519 = ~n1045 & n1233;
  assign n1520 = n1268 & n1519;
  assign n1521 = n1064 & n1520;
  assign n1522 = n994 & n1521;
  assign n1523 = ~n1066 & n1522;
  assign n1524 = ~n1012 & n1233;
  assign n1525 = n1268 & n1524;
  assign n1526 = n994 & n1525;
  assign n1527 = n1065 & n1526;
  assign n1528 = ~n1523 & ~n1527;
  assign n1529 = ~n1518 & n1528;
  assign n1530 = n1262 & n1349;
  assign n1531 = ~n1248 & n1530;
  assign n1532 = n1236 & n1531;
  assign n1533 = n1233 & n1532;
  assign n1534 = n922 & n1533;
  assign n1535 = ~n1262 & n1356;
  assign n1536 = ~n1248 & n1535;
  assign n1537 = n1236 & n1536;
  assign n1538 = n1233 & n1537;
  assign n1539 = n922 & n1538;
  assign n1540 = n1262 & n1362;
  assign n1541 = ~n1248 & n1540;
  assign n1542 = ~n1236 & n1541;
  assign n1543 = n1233 & n1542;
  assign n1544 = n922 & n1543;
  assign n1545 = ~n1262 & n1368;
  assign n1546 = ~n1248 & n1545;
  assign n1547 = ~n1236 & n1546;
  assign n1548 = n1233 & n1547;
  assign n1549 = n922 & n1548;
  assign n1550 = n1248 & n1530;
  assign n1551 = n1236 & n1550;
  assign n1552 = n1233 & n1551;
  assign n1553 = n1064 & n1552;
  assign n1554 = n1248 & n1535;
  assign n1555 = n1236 & n1554;
  assign n1556 = n1233 & n1555;
  assign n1557 = n1064 & n1556;
  assign n1558 = n1248 & n1540;
  assign n1559 = ~n1236 & n1558;
  assign n1560 = n1233 & n1559;
  assign n1561 = n1064 & n1560;
  assign n1562 = n1248 & n1545;
  assign n1563 = ~n1236 & n1562;
  assign n1564 = n1233 & n1563;
  assign n1565 = n1064 & n1564;
  assign n1566 = n1529 & ~n1565;
  assign n1567 = ~n1561 & n1566;
  assign n1568 = ~n1557 & n1567;
  assign n1569 = ~n1553 & n1568;
  assign n1570 = ~n1549 & n1569;
  assign n1571 = ~n1544 & n1570;
  assign n1572 = ~n1539 & n1571;
  assign n1573 = ~n1534 & n1572;
  assign n1574 = ~n1005 & ~n1038;
  assign n1575 = ~n1443 & n1574;
  assign n1576 = ~n1005 & n1424;
  assign n1577 = ~n1440 & n1576;
  assign n1578 = n996 & n1577;
  assign n1579 = n1065 & n1578;
  assign n1580 = n1005 & n1424;
  assign n1581 = ~n1440 & n1580;
  assign n1582 = n996 & n1581;
  assign n1583 = n1066 & n1582;
  assign n1584 = ~n1579 & ~n1583;
  assign n1585 = n1434 & n1462;
  assign n1586 = n1427 & n1585;
  assign n1587 = n1424 & n1586;
  assign n1588 = n1066 & n1587;
  assign n1589 = ~\V1213(2)  & n1575;
  assign n1590 = ~n1434 & n1589;
  assign n1591 = n1424 & n1590;
  assign n1592 = n1065 & n1591;
  assign n1593 = ~n1427 & n1477;
  assign n1594 = n1424 & n1593;
  assign n1595 = n1066 & n1594;
  assign n1596 = n1584 & ~n1595;
  assign n1597 = ~n1592 & n1596;
  assign n1598 = ~n1588 & n1597;
  assign n1599 = ~n1019 & n1055;
  assign n1600 = n979 & n1599;
  assign n1601 = ~\V1213(0)  & n1600;
  assign n1602 = ~\V1213(2)  & n1601;
  assign n1603 = n943 & n1602;
  assign n1604 = n922 & n1603;
  assign n1605 = n993 & n1604;
  assign n1606 = ~n1019 & ~n1055;
  assign n1607 = n979 & n1606;
  assign n1608 = \V1213(0)  & n1607;
  assign n1609 = ~\V1213(2)  & n1608;
  assign n1610 = n943 & n1609;
  assign n1611 = n922 & n1610;
  assign n1612 = n993 & n1611;
  assign n1613 = ~n979 & n1599;
  assign n1614 = ~\V1213(0)  & n1613;
  assign n1615 = \V1213(2)  & n1614;
  assign n1616 = n943 & n1615;
  assign n1617 = n922 & n1616;
  assign n1618 = n993 & n1617;
  assign n1619 = ~n979 & n1606;
  assign n1620 = \V1213(0)  & n1619;
  assign n1621 = \V1213(2)  & n1620;
  assign n1622 = n943 & n1621;
  assign n1623 = n922 & n1622;
  assign n1624 = n993 & n1623;
  assign n1625 = n1019 & n1055;
  assign n1626 = n979 & n1625;
  assign n1627 = ~\V1213(0)  & n1626;
  assign n1628 = ~\V1213(2)  & n1627;
  assign n1629 = n943 & n1628;
  assign n1630 = n1064 & n1629;
  assign n1631 = n993 & n1630;
  assign n1632 = n1019 & ~n1055;
  assign n1633 = n979 & n1632;
  assign n1634 = \V1213(0)  & n1633;
  assign n1635 = ~\V1213(2)  & n1634;
  assign n1636 = n943 & n1635;
  assign n1637 = n1064 & n1636;
  assign n1638 = n993 & n1637;
  assign n1639 = ~n979 & n1625;
  assign n1640 = ~\V1213(0)  & n1639;
  assign n1641 = \V1213(2)  & n1640;
  assign n1642 = n943 & n1641;
  assign n1643 = n1064 & n1642;
  assign n1644 = n993 & n1643;
  assign n1645 = ~n979 & n1632;
  assign n1646 = \V1213(0)  & n1645;
  assign n1647 = \V1213(2)  & n1646;
  assign n1648 = n943 & n1647;
  assign n1649 = n1064 & n1648;
  assign n1650 = n993 & n1649;
  assign n1651 = ~n1644 & ~n1650;
  assign n1652 = ~n1638 & n1651;
  assign n1653 = ~n1631 & n1652;
  assign n1654 = ~n1624 & n1653;
  assign n1655 = ~n1618 & n1654;
  assign n1656 = ~n1612 & n1655;
  assign n1657 = ~n1605 & n1656;
  assign n1658 = \V288(0)  & n1059;
  assign n1659 = ~n1029 & n1658;
  assign n1660 = n982 & n1659;
  assign n1661 = ~\V1213(0)  & n1660;
  assign n1662 = ~\V1213(2)  & n1661;
  assign n1663 = n943 & n1662;
  assign n1664 = n922 & n1663;
  assign n1665 = \V288(0)  & ~n1059;
  assign n1666 = ~n1029 & n1665;
  assign n1667 = n982 & n1666;
  assign n1668 = \V1213(0)  & n1667;
  assign n1669 = ~\V1213(2)  & n1668;
  assign n1670 = n943 & n1669;
  assign n1671 = n922 & n1670;
  assign n1672 = ~n982 & n1659;
  assign n1673 = ~\V1213(0)  & n1672;
  assign n1674 = \V1213(2)  & n1673;
  assign n1675 = n943 & n1674;
  assign n1676 = n922 & n1675;
  assign n1677 = ~n982 & n1666;
  assign n1678 = \V1213(0)  & n1677;
  assign n1679 = \V1213(2)  & n1678;
  assign n1680 = n943 & n1679;
  assign n1681 = n922 & n1680;
  assign n1682 = n1029 & n1658;
  assign n1683 = n982 & n1682;
  assign n1684 = ~\V1213(0)  & n1683;
  assign n1685 = ~\V1213(2)  & n1684;
  assign n1686 = n943 & n1685;
  assign n1687 = n1064 & n1686;
  assign n1688 = n1029 & n1665;
  assign n1689 = n982 & n1688;
  assign n1690 = \V1213(0)  & n1689;
  assign n1691 = ~\V1213(2)  & n1690;
  assign n1692 = n943 & n1691;
  assign n1693 = n1064 & n1692;
  assign n1694 = ~n982 & n1682;
  assign n1695 = ~\V1213(0)  & n1694;
  assign n1696 = \V1213(2)  & n1695;
  assign n1697 = n943 & n1696;
  assign n1698 = n1064 & n1697;
  assign n1699 = ~n982 & n1688;
  assign n1700 = \V1213(0)  & n1699;
  assign n1701 = \V1213(2)  & n1700;
  assign n1702 = n943 & n1701;
  assign n1703 = n1064 & n1702;
  assign n1704 = n1657 & ~n1703;
  assign n1705 = ~n1698 & n1704;
  assign n1706 = ~n1693 & n1705;
  assign n1707 = ~n1687 & n1706;
  assign n1708 = ~n1681 & n1707;
  assign n1709 = ~n1676 & n1708;
  assign n1710 = ~n1671 & n1709;
  assign n1711 = ~n1664 & n1710;
  assign n1712 = \V1213(3)  & n1487;
  assign n1713 = n1488 & n1712;
  assign n1714 = n527 & \V1213(2) ;
  assign n1715 = ~n1713 & n1714;
  assign n1716 = n1711 & n1715;
  assign n1717 = n1598 & n1716;
  assign n1718 = n1573 & n1717;
  assign n1719 = n527 & n1711;
  assign n1720 = ~n1712 & n1719;
  assign n1721 = n1598 & n1720;
  assign n1722 = n1573 & n1721;
  assign V357 = n1718 | n1722;
  assign n1724 = ~\V149(7)  & n496;
  assign n1725 = \V33(0)  & \V289(0) ;
  assign n1726 = ~n499 & n1725;
  assign \V1745(0)  = n1724 | ~n1726;
  assign n1728 = \V149(7)  & ~\V149(6) ;
  assign n1729 = n531 & n1728;
  assign n1730 = n918 & n1729;
  assign n1731 = \V56(0)  & n1730;
  assign n1732 = \V108(0)  & ~n1731;
  assign n1733 = \V16(0)  & \V15(0) ;
  assign n1734 = n861 & ~n1733;
  assign \V1896(0)  = n1732 | ~n1734;
  assign n1736 = n559 & n782;
  assign n1737 = n559 & n659;
  assign n1738 = \V118(4)  & n1736;
  assign n1739 = \V132(6)  & n1737;
  assign \V1953(6)  = n1738 | n1739;
  assign n1741 = \V118(5)  & n1736;
  assign n1742 = \V132(7)  & n1737;
  assign \V1953(7)  = n1741 | n1742;
  assign n1744 = \V1953(6)  & ~\V1953(7) ;
  assign n1745 = ~\V1953(6)  & \V1953(7) ;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = n528 & n784;
  assign n1748 = n528 & n558;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = \V46(0)  & ~n1749;
  assign n1751 = \V118(7)  & n1736;
  assign \V1960(1)  = n1750 | n1751;
  assign n1753 = ~n1746 & \V1960(1) ;
  assign n1754 = n1746 & ~\V1960(1) ;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = \V48(0)  & ~n1749;
  assign n1757 = \V118(6)  & n1736;
  assign \V1960(0)  = n1756 | n1757;
  assign n1759 = ~n1755 & \V1960(0) ;
  assign n1760 = n1755 & ~\V1960(0) ;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = \V118(2)  & n1736;
  assign n1763 = \V132(4)  & n1737;
  assign \V1953(4)  = n1762 | n1763;
  assign n1765 = \V118(3)  & n1736;
  assign n1766 = \V132(5)  & n1737;
  assign \V1953(5)  = n1765 | n1766;
  assign n1768 = \V1953(4)  & ~\V1953(5) ;
  assign n1769 = ~\V1953(4)  & \V1953(5) ;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = \V118(1)  & n1736;
  assign n1772 = \V132(3)  & n1737;
  assign \V1953(3)  = n1771 | n1772;
  assign n1774 = ~n1770 & \V1953(3) ;
  assign n1775 = n1770 & ~\V1953(3) ;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = \V118(0)  & n1736;
  assign n1778 = \V132(2)  & n1737;
  assign \V1953(2)  = n1777 | n1778;
  assign n1780 = ~n1776 & \V1953(2) ;
  assign n1781 = n1776 & ~\V1953(2) ;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1761 & ~n1782;
  assign n1784 = n1761 & n1782;
  assign \V1613(1)  = n1783 | n1784;
  assign V373 = \V10(0)  & \V13(0) ;
  assign n1787 = \V203(0)  & ~\V165(0) ;
  assign n1788 = \V165(2)  & n1787;
  assign n1789 = \V165(1)  & n1788;
  assign n1790 = \V203(0)  & \V35(0) ;
  assign V377 = n1789 | n1790;
  assign n1792 = n531 & n782;
  assign n1793 = n495 & n917;
  assign n1794 = \V108(4)  & n1730;
  assign n1795 = \V124(4)  & n1737;
  assign n1796 = \V213(4)  & n1792;
  assign n1797 = \V100(4)  & n1793;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = ~n1795 & n1798;
  assign \V1921(4)  = n1794 | ~n1799;
  assign n1801 = \V124(5)  & n1737;
  assign n1802 = \V213(5)  & n1792;
  assign n1803 = \V100(5)  & n1793;
  assign n1804 = ~n1802 & ~n1803;
  assign \V1921(5)  = n1801 | ~n1804;
  assign n1806 = \V1921(4)  & ~\V1921(5) ;
  assign n1807 = ~\V1921(4)  & \V1921(5) ;
  assign n1808 = ~n1806 & ~n1807;
  assign \V1953(1)  = \V132(1)  & n1737;
  assign n1810 = ~n1808 & \V1953(1) ;
  assign n1811 = n1808 & ~\V1953(1) ;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = \V149(6)  & n918;
  assign n1814 = n917 & n1813;
  assign n1815 = \V132(0)  & n1737;
  assign n1816 = \V108(5)  & n1814;
  assign \V1953(0)  = n1815 | n1816;
  assign n1818 = ~n1812 & \V1953(0) ;
  assign n1819 = n1812 & ~\V1953(0) ;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = \V108(2)  & n1730;
  assign n1822 = \V124(2)  & n1737;
  assign n1823 = \V213(2)  & n1792;
  assign n1824 = \V100(2)  & n1793;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = ~n1822 & n1825;
  assign \V1921(2)  = n1821 | ~n1826;
  assign n1828 = \V108(3)  & n1730;
  assign n1829 = \V124(3)  & n1737;
  assign n1830 = \V213(3)  & n1792;
  assign n1831 = \V100(3)  & n1793;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1829 & n1832;
  assign \V1921(3)  = n1828 | ~n1833;
  assign n1835 = \V1921(2)  & ~\V1921(3) ;
  assign n1836 = ~\V1921(2)  & \V1921(3) ;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = \V108(1)  & n1730;
  assign n1839 = \V124(1)  & n1737;
  assign n1840 = \V213(1)  & n1792;
  assign n1841 = \V100(1)  & n1793;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1839 & n1842;
  assign \V1921(1)  = n1838 | ~n1843;
  assign n1845 = ~n1837 & \V1921(1) ;
  assign n1846 = n1837 & ~\V1921(1) ;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = \V108(0)  & n1730;
  assign n1849 = \V124(0)  & n1737;
  assign n1850 = \V213(0)  & n1792;
  assign n1851 = \V100(0)  & n1793;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~n1849 & n1852;
  assign \V1921(0)  = n1848 | ~n1853;
  assign n1855 = ~n1847 & \V1921(0) ;
  assign n1856 = n1847 & ~\V1921(0) ;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1820 & ~n1857;
  assign n1859 = n1820 & n1857;
  assign \V1613(0)  = n1858 | n1859;
  assign n1861 = ~\V43(0)  & \V45(0) ;
  assign \V511(0)  = \V40(0)  | n1861;
  assign n1863 = \V268(5)  & \V268(4) ;
  assign n1864 = \V268(3)  & \V268(1) ;
  assign n1865 = \V268(2)  & n1864;
  assign n1866 = n1863 & n1865;
  assign n1867 = ~\V56(0)  & ~\V62(0) ;
  assign n1868 = ~\V50(0)  & n1867;
  assign n1869 = ~n527 & ~n1868;
  assign n1870 = ~\V258(0)  & n1869;
  assign n1871 = \V258(0)  & \V268(0) ;
  assign n1872 = n1866 & n1871;
  assign n1873 = ~n1870 & ~n1872;
  assign n1874 = ~\V258(0)  & ~\V259(0) ;
  assign n1875 = ~n1873 & n1874;
  assign n1876 = \V258(0)  & \V259(0) ;
  assign n1877 = ~n1873 & n1876;
  assign n1878 = ~n1875 & ~n1877;
  assign n1879 = ~\V260(0)  & \V14(0) ;
  assign n1880 = ~n1878 & n1879;
  assign n1881 = \V260(0)  & \V14(0) ;
  assign n1882 = n1878 & n1881;
  assign \V1467(0)  = n1880 | n1882;
  assign n1884 = ~n493 & ~n501;
  assign n1885 = n869 & ~n1884;
  assign n1886 = \V14(0)  & ~n1793;
  assign n1887 = ~n1885 & n1886;
  assign n1888 = \V14(0)  & ~\V56(0) ;
  assign n1889 = ~n1885 & n1888;
  assign n1890 = ~n1887 & ~n1889;
  assign n1891 = \V100(2)  & ~n1890;
  assign n1892 = \V165(4)  & n1885;
  assign \V1709(1)  = n1891 | n1892;
  assign n1894 = \V100(1)  & ~n1890;
  assign n1895 = \V165(3)  & n1885;
  assign \V1709(0)  = n1894 | n1895;
  assign n1897 = \V100(4)  & ~n1890;
  assign n1898 = \V165(6)  & n1885;
  assign \V1709(3)  = n1897 | n1898;
  assign n1900 = \V100(3)  & ~n1890;
  assign n1901 = \V165(5)  & n1885;
  assign \V1709(2)  = n1900 | n1901;
  assign n1903 = ~\V214(0)  & ~\V43(0) ;
  assign n1904 = ~\V165(7)  & n867;
  assign n1905 = ~\V302(0)  & ~n1904;
  assign n1906 = ~\V172(0)  & \V240(0) ;
  assign V1719 = ~n867 & n1906;
  assign n1908 = ~n1789 & n1905;
  assign n1909 = V1719 & ~n1908;
  assign n1910 = \V215(0)  & \V66(0) ;
  assign n1911 = ~V763 & ~n542;
  assign n1912 = \V802(0)  & ~n1911;
  assign n1913 = ~\V32(0)  & \V32(2) ;
  assign n1914 = \V32(3)  & n1913;
  assign n1915 = n1055 & n1914;
  assign n1916 = n1019 & n1915;
  assign n1917 = n991 & n1916;
  assign n1918 = \V32(0)  & \V32(2) ;
  assign n1919 = \V32(3)  & n1918;
  assign n1920 = ~n1055 & n1919;
  assign n1921 = n1019 & n1920;
  assign n1922 = n991 & n1921;
  assign n1923 = ~\V32(0)  & \V32(1) ;
  assign n1924 = \V32(2)  & n1923;
  assign n1925 = \V32(3)  & n1924;
  assign n1926 = n1055 & n1925;
  assign n1927 = n991 & n1926;
  assign n1928 = \V32(0)  & \V32(1) ;
  assign n1929 = \V32(2)  & n1928;
  assign n1930 = \V32(3)  & n1929;
  assign n1931 = ~n1055 & n1930;
  assign n1932 = n991 & n1931;
  assign n1933 = ~\V32(0)  & \V32(3) ;
  assign n1934 = n1055 & n1933;
  assign n1935 = n1019 & n1934;
  assign n1936 = n989 & n1935;
  assign n1937 = \V32(0)  & \V32(3) ;
  assign n1938 = ~n1055 & n1937;
  assign n1939 = n1019 & n1938;
  assign n1940 = n989 & n1939;
  assign n1941 = \V32(3)  & n1923;
  assign n1942 = n1055 & n1941;
  assign n1943 = n989 & n1942;
  assign n1944 = \V32(3)  & n1928;
  assign n1945 = ~n1055 & n1944;
  assign n1946 = n989 & n1945;
  assign n1947 = n1055 & n1913;
  assign n1948 = n1019 & n1947;
  assign n1949 = n979 & n1948;
  assign n1950 = ~n1055 & n1918;
  assign n1951 = n1019 & n1950;
  assign n1952 = n979 & n1951;
  assign n1953 = n1055 & n1924;
  assign n1954 = n979 & n1953;
  assign n1955 = ~n1055 & n1929;
  assign n1956 = n979 & n1955;
  assign n1957 = n1055 & n1923;
  assign n1958 = n1019 & n1957;
  assign n1959 = ~n1055 & n1928;
  assign n1960 = n1019 & n1959;
  assign n1961 = \V32(0)  & n1055;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n1958 & n1962;
  assign n1964 = ~n1956 & n1963;
  assign n1965 = ~n1954 & n1964;
  assign n1966 = ~n1952 & n1965;
  assign n1967 = ~n1949 & n1966;
  assign n1968 = ~n1946 & n1967;
  assign n1969 = ~n1943 & n1968;
  assign n1970 = ~n1940 & n1969;
  assign n1971 = ~n1936 & n1970;
  assign n1972 = ~n1932 & n1971;
  assign n1973 = ~n1927 & n1972;
  assign n1974 = ~n1922 & n1973;
  assign n1975 = ~n1917 & n1974;
  assign n1976 = ~n783 & n1749;
  assign n1977 = n531 & n558;
  assign n1978 = \V66(0)  & n1977;
  assign n1979 = ~V763 & ~n1975;
  assign n1980 = ~n811 & n1979;
  assign n1981 = \V56(0)  & ~n1975;
  assign n1982 = ~n1976 & n1981;
  assign n1983 = n656 & n1981;
  assign n1984 = \V66(0)  & V763;
  assign n1985 = ~n1975 & n1984;
  assign n1986 = ~n1975 & n1978;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n1983 & n1987;
  assign n1989 = ~n1982 & n1988;
  assign n1990 = ~n1980 & n1989;
  assign n1991 = n542 & n545;
  assign n1992 = \V802(0)  & n551;
  assign n1993 = n550 & n874;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = n539 & ~n542;
  assign n1996 = ~n538 & n542;
  assign n1997 = ~n553 & ~n1996;
  assign n1998 = ~n1995 & n1997;
  assign n1999 = \V59(0)  & ~n1998;
  assign n2000 = ~n699 & ~n1999;
  assign n2001 = ~\V215(0)  & \V66(0) ;
  assign n2002 = V763 & n2001;
  assign n2003 = ~n867 & n2002;
  assign n2004 = \V802(0)  & n539;
  assign n2005 = \V56(0)  & n1991;
  assign n2006 = n543 & ~n1867;
  assign n2007 = \V802(0)  & n545;
  assign n2008 = \V802(0)  & ~n527;
  assign n2009 = \V70(0)  & ~n527;
  assign n2010 = \V59(0)  & ~n527;
  assign n2011 = \V802(0)  & n553;
  assign n2012 = \V56(0)  & \V174(0) ;
  assign n2013 = ~V1719 & n2000;
  assign n2014 = n1994 & n2013;
  assign n2015 = ~n2012 & n2014;
  assign n2016 = ~n2011 & n2015;
  assign n2017 = ~n2010 & n2016;
  assign n2018 = ~n2009 & n2017;
  assign n2019 = ~n2008 & n2018;
  assign n2020 = ~n2007 & n2019;
  assign n2021 = ~n2006 & n2020;
  assign n2022 = ~n2005 & n2021;
  assign n2023 = ~n2004 & n2022;
  assign \V423(0)  = n2003 | ~n2023;
  assign n2025 = \V32(9)  & n613;
  assign n2026 = \V199(2)  & n616;
  assign n2027 = \V239(2)  & n617;
  assign n2028 = \V84(5)  & n621;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~n2026 & n2029;
  assign \V1243(7)  = n2025 | ~n2030;
  assign n2032 = \V32(10)  & n613;
  assign n2033 = \V199(3)  & n616;
  assign n2034 = \V239(3)  & n617;
  assign n2035 = \V88(0)  & n621;
  assign n2036 = ~n2034 & ~n2035;
  assign n2037 = ~n2033 & n2036;
  assign \V1243(8)  = n2032 | ~n2037;
  assign n2039 = \V32(11)  & n613;
  assign n2040 = \V199(4)  & n616;
  assign n2041 = \V239(4)  & n617;
  assign n2042 = \V88(1)  & n621;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = ~n2040 & n2043;
  assign \V1243(9)  = n2039 | ~n2044;
  assign n2046 = n1421 & n1573;
  assign n2047 = n1486 & n1598;
  assign n2048 = \V288(7)  & \V288(6) ;
  assign n2049 = ~\V248(0)  & n2048;
  assign n2050 = \V1243(9)  & n2049;
  assign n2051 = \V1243(8)  & n2050;
  assign n2052 = \V1243(7)  & n2051;
  assign n2053 = V1719 & n2052;
  assign n2054 = ~n527 & n2053;
  assign n2055 = ~\V248(0)  & \V1243(9) ;
  assign n2056 = \V1243(8)  & n2055;
  assign n2057 = \V1243(7)  & n2056;
  assign n2058 = V1719 & n2057;
  assign n2059 = n994 & n2058;
  assign n2060 = ~n2046 & n2059;
  assign n2061 = n996 & n2058;
  assign n2062 = ~n2047 & n2061;
  assign n2063 = n993 & n2058;
  assign n2064 = ~n1230 & n2063;
  assign n2065 = ~n1711 & n2063;
  assign n2066 = ~\V248(0)  & \V288(7) ;
  assign n2067 = \V1243(9)  & n2066;
  assign n2068 = \V1243(8)  & n2067;
  assign n2069 = \V1243(7)  & n2068;
  assign n2070 = V1719 & n2069;
  assign n2071 = n1487 & n2070;
  assign n2072 = ~n527 & n2058;
  assign n2073 = n996 & n2072;
  assign n2074 = n994 & n2072;
  assign n2075 = ~\V248(0)  & \V243(0) ;
  assign n2076 = \V244(0)  & n2075;
  assign n2077 = \V245(0)  & n2076;
  assign n2078 = \V246(0)  & n2077;
  assign n2079 = \V247(0)  & n2078;
  assign n2080 = V1719 & n2079;
  assign n2081 = ~\V248(0)  & V1719;
  assign n2082 = n905 & n2081;
  assign n2083 = ~n2080 & ~n2082;
  assign n2084 = ~n2074 & n2083;
  assign n2085 = ~n2073 & n2084;
  assign n2086 = ~n2071 & n2085;
  assign n2087 = ~n2065 & n2086;
  assign n2088 = ~n2064 & n2087;
  assign n2089 = ~n2062 & n2088;
  assign n2090 = ~n2060 & n2089;
  assign \V393(0)  = n2054 | ~n2090;
  assign n2092 = ~\V15(0)  & ~\V393(0) ;
  assign n2093 = \V423(0)  & n2092;
  assign n2094 = n861 & n2093;
  assign n2095 = n527 & n2094;
  assign n2096 = n1990 & n2095;
  assign n2097 = n647 & n2096;
  assign n2098 = ~n1912 & n2097;
  assign n2099 = ~n1910 & n2098;
  assign n2100 = ~n1909 & n2099;
  assign V432 = n1903 & n2100;
  assign n2102 = \V100(5)  & ~n1890;
  assign n2103 = \V165(7)  & n1885;
  assign \V1709(4)  = n2102 | n2103;
  assign n2105 = n499 & n665;
  assign n2106 = \V108(2)  & ~n1731;
  assign \V1898(0)  = n2105 | n2106;
  assign n2108 = ~\V290(0)  & n867;
  assign n2109 = n691 & ~n2108;
  assign n2110 = n1905 & n2109;
  assign n2111 = \V14(0)  & n2110;
  assign n2112 = \V165(3)  & n2111;
  assign n2113 = n514 & n2112;
  assign n2114 = n487 & n2113;
  assign n2115 = \V65(0)  & ~n1748;
  assign n2116 = ~n543 & n2115;
  assign n2117 = n2111 & n2116;
  assign \V1392(0)  = n2114 | n2117;
  assign n2119 = \V32(11)  & n612;
  assign n2120 = \V32(8)  & n613;
  assign n2121 = \V199(1)  & n616;
  assign n2122 = \V239(1)  & n617;
  assign n2123 = \V84(4)  & n621;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = ~n2121 & n2124;
  assign n2126 = ~n2120 & n2125;
  assign \V1243(6)  = n2119 | ~n2126;
  assign n2128 = ~\V38(0)  & ~\V39(0) ;
  assign n2129 = ~\V42(0)  & n2128;
  assign n2130 = ~\V44(0)  & n2129;
  assign n2131 = \V38(0)  & \V39(0) ;
  assign n2132 = ~\V42(0)  & n2131;
  assign n2133 = ~\V44(0)  & n2132;
  assign n2134 = \V42(0)  & n2131;
  assign n2135 = \V44(0)  & n2134;
  assign n2136 = \V42(0)  & n2128;
  assign n2137 = \V44(0)  & n2136;
  assign n2138 = ~n2135 & ~n2137;
  assign n2139 = ~n2133 & n2138;
  assign V512 = n2130 | ~n2139;
  assign n2141 = \V246(0)  & ~\V247(0) ;
  assign n2142 = ~\V603(0)  & n2141;
  assign n2143 = ~n874 & n2142;
  assign n2144 = \V247(0)  & \V603(0) ;
  assign n2145 = ~\V246(0)  & \V247(0) ;
  assign n2146 = ~n874 & n2145;
  assign n2147 = ~n2144 & ~n2146;
  assign \V609(0)  = n2143 | ~n2147;
  assign n2149 = \V62(0)  & n543;
  assign n2150 = n2000 & ~n2149;
  assign n2151 = n647 & ~n867;
  assign n2152 = ~n2150 & n2151;
  assign V527 = n1903 & n2152;
  assign V537 = n547 & \V1213(0) ;
  assign V538 = n547 & \V1213(1) ;
  assign V539 = n547 & \V1213(2) ;
  assign V540 = n547 & \V1213(3) ;
  assign n2158 = \V183(4)  & n616;
  assign n2159 = \V223(4)  & n617;
  assign n2160 = \V32(4)  & n621;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n2158 & n2161;
  assign \V1213(4)  = n633 | ~n2162;
  assign V541 = n547 & \V1213(4) ;
  assign n2165 = \V257(0)  & n607;
  assign n2166 = \V183(5)  & n616;
  assign n2167 = \V223(5)  & n617;
  assign n2168 = \V32(5)  & n621;
  assign n2169 = ~n612 & ~n2168;
  assign n2170 = ~n2167 & n2169;
  assign n2171 = ~n2166 & n2170;
  assign \V1213(5)  = n2165 | ~n2171;
  assign V542 = n547 & \V1213(5) ;
  assign n2174 = \V257(1)  & n607;
  assign n2175 = \V189(0)  & n616;
  assign n2176 = \V229(0)  & n617;
  assign n2177 = \V32(6)  & n621;
  assign n2178 = ~n613 & ~n2177;
  assign n2179 = ~n2176 & n2178;
  assign n2180 = ~n2175 & n2179;
  assign \V1213(6)  = n2174 | ~n2180;
  assign V543 = n547 & \V1213(6) ;
  assign n2183 = \V257(2)  & n607;
  assign n2184 = \V189(1)  & n616;
  assign n2185 = \V229(1)  & n617;
  assign n2186 = \V32(7)  & n621;
  assign n2187 = \V32(0)  & n608;
  assign n2188 = ~n613 & ~n2187;
  assign n2189 = ~n2186 & n2188;
  assign n2190 = ~n2185 & n2189;
  assign n2191 = ~n2184 & n2190;
  assign \V1213(7)  = n2183 | ~n2191;
  assign V544 = n547 & \V1213(7) ;
  assign n2194 = \V257(3)  & n607;
  assign n2195 = \V189(2)  & n616;
  assign n2196 = \V229(2)  & n617;
  assign n2197 = \V32(8)  & n621;
  assign n2198 = \V32(1)  & n608;
  assign n2199 = ~n613 & ~n2198;
  assign n2200 = ~n2197 & n2199;
  assign n2201 = ~n2196 & n2200;
  assign n2202 = ~n2195 & n2201;
  assign \V1213(8)  = n2194 | ~n2202;
  assign V545 = n547 & \V1213(8) ;
  assign n2205 = \V257(4)  & n607;
  assign n2206 = \V189(3)  & n616;
  assign n2207 = \V229(3)  & n617;
  assign n2208 = \V32(9)  & n621;
  assign n2209 = \V32(2)  & n608;
  assign n2210 = ~n613 & ~n2209;
  assign n2211 = ~n2208 & n2210;
  assign n2212 = ~n2207 & n2211;
  assign n2213 = ~n2206 & n2212;
  assign \V1213(9)  = n2205 | ~n2213;
  assign V546 = n547 & \V1213(9) ;
  assign V547 = n547 & \V1213(10) ;
  assign V548 = n547 & \V1213(11) ;
  assign n2218 = ~n783 & ~n1747;
  assign n2219 = ~n1792 & ~n1793;
  assign n2220 = ~n1737 & n2219;
  assign n2221 = ~\V59(0)  & \V258(0) ;
  assign n2222 = ~\V259(0)  & n2221;
  assign n2223 = ~\V260(0)  & n2222;
  assign n2224 = n491 & n782;
  assign n2225 = ~n785 & ~n1736;
  assign n2226 = ~n2224 & n2225;
  assign n2227 = ~n2223 & n2226;
  assign n2228 = n2220 & n2227;
  assign n2229 = n527 & ~n785;
  assign n2230 = ~n1736 & n2229;
  assign n2231 = ~n2224 & n2230;
  assign n2232 = n2220 & n2231;
  assign n2233 = ~n2228 & ~n2232;
  assign n2234 = \V62(0)  & ~n2218;
  assign n2235 = \V65(0)  & n1748;
  assign n2236 = \V56(0)  & n2233;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n2234 & n2237;
  assign n2239 = ~n1789 & n2110;
  assign n2240 = \V149(0)  & ~n500;
  assign n2241 = \V14(0)  & ~\V289(0) ;
  assign n2242 = \V165(7)  & n2108;
  assign n2243 = ~\V1741(0)  & ~n2238;
  assign n2244 = ~n1904 & n2243;
  assign n2245 = n653 & ~n2239;
  assign n2246 = n527 & n2240;
  assign n2247 = \V290(0)  & ~n867;
  assign n2248 = ~\V302(0)  & ~\V214(0) ;
  assign n2249 = ~n2242 & n2248;
  assign n2250 = n2241 & n2249;
  assign n2251 = ~n2247 & n2250;
  assign n2252 = ~n2246 & n2251;
  assign n2253 = ~n2245 & n2252;
  assign \V798(0)  = n2244 | ~n2253;
  assign n2255 = \V149(5)  & n747;
  assign n2256 = \V32(6)  & n612;
  assign n2257 = \V32(3)  & n613;
  assign n2258 = \V194(1)  & n616;
  assign n2259 = \V234(1)  & n617;
  assign n2260 = \V78(5)  & n621;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2258 & n2261;
  assign n2263 = ~n2257 & n2262;
  assign n2264 = ~n2256 & n2263;
  assign \V1243(1)  = n2255 | ~n2264;
  assign n2266 = \V149(7)  & n747;
  assign n2267 = \V32(8)  & n612;
  assign n2268 = \V32(5)  & n613;
  assign n2269 = \V194(3)  & n616;
  assign n2270 = \V234(3)  & n617;
  assign n2271 = \V84(1)  & n621;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = ~n2269 & n2272;
  assign n2274 = ~n2268 & n2273;
  assign n2275 = ~n2267 & n2274;
  assign \V1243(3)  = n2266 | ~n2275;
  assign n2277 = \V149(6)  & n747;
  assign n2278 = \V32(7)  & n612;
  assign n2279 = \V32(4)  & n613;
  assign n2280 = \V194(2)  & n616;
  assign n2281 = \V234(2)  & n617;
  assign n2282 = \V84(0)  & n621;
  assign n2283 = ~n2281 & ~n2282;
  assign n2284 = ~n2280 & n2283;
  assign n2285 = ~n2279 & n2284;
  assign n2286 = ~n2278 & n2285;
  assign \V1243(2)  = n2277 | ~n2286;
  assign n2288 = n486 & \V802(0) ;
  assign n2289 = ~n807 & ~n2288;
  assign n2290 = \V271(0)  & ~\V274(0) ;
  assign n2291 = ~n560 & n2290;
  assign n2292 = \V134(1)  & \V134(0) ;
  assign n2293 = ~n550 & n2292;
  assign n2294 = ~n906 & n2293;
  assign n2295 = n2291 & n2294;
  assign n2296 = ~n651 & n686;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = n2289 & ~n2297;
  assign n2299 = n807 & n2297;
  assign n2300 = n2288 & n2297;
  assign n2301 = ~\V194(3)  & n2298;
  assign n2302 = n902 & n2301;
  assign n2303 = \V194(3)  & n2298;
  assign n2304 = ~n902 & n2303;
  assign n2305 = \V1243(3)  & n2299;
  assign n2306 = \V149(7)  & n2300;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2304 & n2307;
  assign \V572(3)  = n2302 | ~n2308;
  assign n2310 = \V32(10)  & n612;
  assign n2311 = \V32(7)  & n613;
  assign n2312 = \V199(0)  & n616;
  assign n2313 = \V239(0)  & n617;
  assign n2314 = \V84(3)  & n621;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n2312 & n2315;
  assign n2317 = ~n2311 & n2316;
  assign \V1243(5)  = n2310 | ~n2317;
  assign n2319 = ~\V194(2)  & n2298;
  assign n2320 = n903 & n2319;
  assign n2321 = \V194(2)  & n2298;
  assign n2322 = ~n903 & n2321;
  assign n2323 = \V1243(2)  & n2299;
  assign n2324 = \V149(6)  & n2300;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n2322 & n2325;
  assign \V572(2)  = n2320 | ~n2326;
  assign n2328 = \V32(9)  & n612;
  assign n2329 = \V32(6)  & n613;
  assign n2330 = \V194(4)  & n616;
  assign n2331 = \V234(4)  & n617;
  assign n2332 = \V84(2)  & n621;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = ~n2330 & n2333;
  assign n2335 = ~n2329 & n2334;
  assign \V1243(4)  = n2328 | ~n2335;
  assign n2337 = \V199(1)  & ~n901;
  assign n2338 = n2298 & n2337;
  assign n2339 = n899 & n2338;
  assign n2340 = \V199(0)  & ~n901;
  assign n2341 = n2298 & n2340;
  assign n2342 = n2299 & \V1243(5) ;
  assign n2343 = ~n2341 & ~n2342;
  assign \V572(5)  = n2339 | ~n2343;
  assign n2345 = \V194(4)  & ~n901;
  assign n2346 = n2298 & n2345;
  assign n2347 = ~\V194(4)  & n901;
  assign n2348 = n2298 & n2347;
  assign n2349 = n2299 & \V1243(4) ;
  assign n2350 = ~n2348 & ~n2349;
  assign \V572(4)  = n2346 | ~n2350;
  assign n2352 = n499 & n869;
  assign n2353 = \V14(0)  & ~n1792;
  assign n2354 = ~n2352 & n2353;
  assign n2355 = n1888 & ~n2352;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = ~\V165(7)  & ~\V165(6) ;
  assign n2358 = ~\V165(3)  & n2357;
  assign n2359 = n487 & n2358;
  assign n2360 = n647 & ~n2359;
  assign n2361 = n499 & n868;
  assign n2362 = \V213(0)  & ~n2356;
  assign n2363 = n2352 & ~n2360;
  assign n2364 = ~n2362 & ~n2363;
  assign \V1281(0)  = n2361 | ~n2364;
  assign n2366 = \V194(2)  & ~n905;
  assign n2367 = n2298 & n2366;
  assign n2368 = n903 & n2367;
  assign n2369 = \V194(1)  & ~n905;
  assign n2370 = n2298 & n2369;
  assign n2371 = \V149(5)  & n2300;
  assign n2372 = \V1243(1)  & n2299;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~n2370 & n2373;
  assign \V572(1)  = n2368 | ~n2374;
  assign n2376 = n783 & n861;
  assign n2377 = \V62(0)  & n1748;
  assign n2378 = ~n551 & ~n557;
  assign n2379 = \V56(0)  & ~n2378;
  assign n2380 = \V56(0)  & n2376;
  assign n2381 = ~n650 & ~n2380;
  assign n2382 = ~n2379 & n2381;
  assign n2383 = ~n2377 & n2382;
  assign n2384 = ~n2376 & n2383;
  assign n2385 = ~n1991 & n2384;
  assign n2386 = ~n647 & ~n2377;
  assign n2387 = ~n2376 & n2386;
  assign n2388 = ~n1991 & n2387;
  assign n2389 = ~\V59(0)  & n2382;
  assign n2390 = ~n2377 & n2389;
  assign n2391 = ~\V214(0)  & ~n867;
  assign n2392 = ~\V59(0)  & ~n647;
  assign n2393 = ~n2377 & n2392;
  assign n2394 = n2391 & ~n2393;
  assign n2395 = ~n2390 & n2394;
  assign n2396 = ~n2388 & n2395;
  assign V620 = n2385 | ~n2396;
  assign n2398 = \V41(0)  & \V45(0) ;
  assign n2399 = ~\V41(0)  & ~\V45(0) ;
  assign n2400 = ~n2398 & ~n2399;
  assign V621 = \V293(0)  & ~n2400;
  assign n2402 = \V194(0)  & ~n905;
  assign n2403 = n2298 & n2402;
  assign n2404 = ~\V194(0)  & n905;
  assign n2405 = n2298 & n2404;
  assign n2406 = ~\V321(2)  & n2299;
  assign n2407 = \V149(4)  & n2300;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = ~n2405 & n2408;
  assign \V572(0)  = n2403 | ~n2409;
  assign n2411 = \V59(0)  & ~\V302(0) ;
  assign n2412 = ~n550 & n2411;
  assign n2413 = n653 & n2412;
  assign n2414 = \V56(0)  & ~\V62(0) ;
  assign n2415 = ~\V302(0)  & n2414;
  assign n2416 = n560 & n2415;
  assign n2417 = ~\V302(0)  & ~n550;
  assign n2418 = n874 & n2417;
  assign n2419 = ~\V302(0)  & \V270(0) ;
  assign n2420 = ~n560 & n2419;
  assign n2421 = ~\V302(0)  & ~\V62(0) ;
  assign n2422 = \V270(0)  & n2421;
  assign n2423 = ~n2420 & ~n2422;
  assign n2424 = ~n2418 & n2423;
  assign n2425 = ~n2416 & n2424;
  assign V630 = n2413 | ~n2425;
  assign n2427 = n542 & n868;
  assign n2428 = n2241 & n2427;
  assign n2429 = n529 & n2428;
  assign n2430 = ~\V302(0)  & ~n867;
  assign n2431 = n692 & n2430;
  assign n2432 = n2241 & n2431;
  assign n2433 = n656 & n868;
  assign n2434 = n2241 & n2433;
  assign n2435 = n660 & n868;
  assign n2436 = n2241 & n2435;
  assign n2437 = ~n2434 & ~n2436;
  assign n2438 = ~n2432 & n2437;
  assign n2439 = ~n2429 & n2438;
  assign n2440 = \V100(0)  & ~n1890;
  assign n2441 = n1885 & ~n2360;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~n1724 & n2439;
  assign n2444 = ~n1884 & n2443;
  assign n2445 = n868 & n2444;
  assign \V1693(0)  = ~n2442 | n2445;
  assign n2447 = \V257(7)  & \V257(6) ;
  assign n2448 = \V257(3)  & \V257(5) ;
  assign n2449 = \V257(4)  & n2448;
  assign n2450 = n2447 & n2449;
  assign n2451 = \V257(2)  & n2450;
  assign n2452 = \V257(1)  & ~n2451;
  assign n2453 = ~\V257(1)  & n2451;
  assign V651 = n2452 | n2453;
  assign n2455 = \V257(1)  & ~V651;
  assign n2456 = \V257(0)  & ~n2455;
  assign n2457 = ~\V257(0)  & n2455;
  assign V650 = n2456 | n2457;
  assign n2459 = ~\V257(2)  & n2450;
  assign n2460 = \V257(2)  & ~n2450;
  assign V652 = n2459 | n2460;
  assign n2462 = \V257(5)  & ~n2447;
  assign n2463 = ~\V257(5)  & n2447;
  assign V655 = n2462 | n2463;
  assign n2465 = \V257(5)  & ~V655;
  assign n2466 = \V257(4)  & ~n2465;
  assign n2467 = ~\V257(4)  & n2465;
  assign V654 = n2466 | n2467;
  assign n2469 = \V257(4)  & ~V654;
  assign n2470 = ~n2450 & n2469;
  assign n2471 = \V257(3)  & ~n2450;
  assign V653 = n2470 | n2471;
  assign n2473 = ~\V257(7)  & \V257(6) ;
  assign n2474 = \V257(7)  & ~\V257(6) ;
  assign V656 = n2473 | n2474;
  assign n2476 = ~\V244(0)  & ~V587;
  assign n2477 = ~n874 & n2476;
  assign n2478 = \V244(0)  & V587;
  assign \V591(0)  = n2477 | n2478;
  assign n2480 = ~\V199(2)  & n2298;
  assign n2481 = n898 & n2480;
  assign n2482 = \V199(2)  & n2298;
  assign n2483 = ~n898 & n2482;
  assign n2484 = \V1243(7)  & n2299;
  assign n2485 = ~n2483 & ~n2484;
  assign \V572(7)  = n2481 | ~n2485;
  assign n2487 = ~\V199(1)  & n2298;
  assign n2488 = n899 & n2487;
  assign n2489 = \V199(1)  & n2298;
  assign n2490 = ~n899 & n2489;
  assign n2491 = \V1243(6)  & n2299;
  assign n2492 = ~n2490 & ~n2491;
  assign \V572(6)  = n2488 | ~n2492;
  assign n2494 = \V1243(9)  & n2299;
  assign n2495 = ~\V199(4)  & n2298;
  assign \V572(9)  = n2494 | n2495;
  assign n2497 = ~\V199(3)  & \V199(4) ;
  assign n2498 = n2298 & n2497;
  assign n2499 = \V199(3)  & ~\V199(4) ;
  assign n2500 = n2298 & n2499;
  assign n2501 = \V1243(8)  & n2299;
  assign n2502 = ~n2500 & ~n2501;
  assign \V572(8)  = n2498 | ~n2502;
  assign n2504 = \V134(1)  & n2289;
  assign n2505 = ~n2291 & n2504;
  assign n2506 = ~\V134(1)  & n2289;
  assign n2507 = n2291 & n2506;
  assign \V1992(1)  = n2505 | n2507;
  assign n2509 = ~\V134(0)  & ~\V1992(1) ;
  assign n2510 = n2289 & n2509;
  assign n2511 = n2291 & n2510;
  assign n2512 = \V134(0)  & \V1992(1) ;
  assign n2513 = \V134(0)  & n2289;
  assign n2514 = ~n2291 & n2513;
  assign n2515 = ~n2512 & ~n2514;
  assign \V1992(0)  = n2511 | ~n2515;
  assign n2517 = ~n526 & n2111;
  assign V775 = n514 & n2517;
  assign V778 = \V5(0)  & \V9(0) ;
  assign n2520 = \V10(0)  & ~\V13(0) ;
  assign V779 = \V6(0)  & n2520;
  assign V780 = \V9(0)  & \V6(0) ;
  assign n2523 = \V56(0)  & n496;
  assign n2524 = ~\V174(0)  & \V6(0) ;
  assign n2525 = \V12(0)  & n2524;
  assign n2526 = n2523 & n2525;
  assign n2527 = \V52(0)  & \V6(0) ;
  assign n2528 = \V12(0)  & n2527;
  assign V781 = n2526 | n2528;
  assign V782 = \V7(0)  & n2520;
  assign V783 = \V5(0)  & \V11(0) ;
  assign V784 = \V7(0)  & \V11(0) ;
  assign V787 = \V7(0)  & \V9(0) ;
  assign V1263 = \V9(0)  & \V4(0) ;
  assign n2535 = ~\V71(0)  & V1263;
  assign n2536 = ~\V202(0)  & V1263;
  assign n2537 = \V13(0)  & V1263;
  assign n2538 = ~n2536 & ~n2537;
  assign V789 = n2535 | ~n2538;
  assign V801 = n490 & ~n496;
  assign n2541 = ~n920 & ~n1730;
  assign n2542 = ~n1814 & n2541;
  assign n2543 = n918 & n2542;
  assign n2544 = ~n660 & ~n1737;
  assign n2545 = n659 & n2544;
  assign n2546 = ~n2543 & ~n2545;
  assign n2547 = ~\V174(0)  & V763;
  assign n2548 = n496 & n2547;
  assign n2549 = n2546 & ~n2548;
  assign n2550 = \V56(0)  & n2111;
  assign n2551 = ~n2549 & n2550;
  assign n2552 = \V802(0)  & n2111;
  assign n2553 = ~n2240 & n2552;
  assign n2554 = n490 & n496;
  assign n2555 = n2111 & n2554;
  assign n2556 = n2008 & n2111;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = ~n2553 & n2557;
  assign V966 = n2551 | ~n2558;
  assign n2560 = n651 & n2378;
  assign n2561 = \V62(0)  & n2111;
  assign n2562 = \V56(0)  & ~n2233;
  assign n2563 = n2111 & n2562;
  assign n2564 = n2549 & n2563;
  assign n2565 = ~n527 & n2561;
  assign n2566 = \V59(0)  & n2111;
  assign n2567 = ~n2560 & n2566;
  assign n2568 = ~n2565 & ~n2567;
  assign V986 = n2564 | ~n2568;
  assign n2570 = \V14(0)  & \V215(0) ;
  assign n2571 = \V69(0)  & n2570;
  assign n2572 = n672 & n2571;
  assign n2573 = \V68(0)  & n2570;
  assign n2574 = n672 & n2573;
  assign n2575 = \V215(0)  & \V70(0) ;
  assign n2576 = \V14(0)  & n2575;
  assign n2577 = n672 & n2576;
  assign n2578 = \V14(0)  & n672;
  assign n2579 = n1910 & n2578;
  assign n2580 = ~\V214(0)  & \V216(0) ;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2577 & n2581;
  assign n2583 = ~n2574 & n2582;
  assign \V1492(0)  = n2572 | ~n2583;
  assign \V500(0)  = \V271(0)  | ~\V14(0) ;
  assign n2586 = \V56(0)  & n1814;
  assign n2587 = \V16(0)  & ~\V15(0) ;
  assign n2588 = \V108(5)  & ~n2586;
  assign \V1901(0)  = n2587 | n2588;
  assign n2590 = ~n551 & V1719;
  assign n2591 = n2239 & n2590;
  assign n2592 = \V280(0)  & V1719;
  assign n2593 = n2239 & n2592;
  assign n2594 = n1994 & ~n2593;
  assign \V1717(0)  = n2591 | ~n2594;
  assign n2596 = ~\V271(0)  & ~\V202(0) ;
  assign n2597 = ~\V269(0)  & \V271(0) ;
  assign n2598 = ~n732 & ~n2597;
  assign \V634(0)  = n2596 | ~n2598;
  assign n2600 = \V277(0)  & \V14(0) ;
  assign n2601 = ~n547 & n2600;
  assign \V1439(0)  = n2224 | n2601;
  assign V1423 = \V1(0)  & \V9(0) ;
  assign V1387 = \V9(0)  & \V8(0) ;
  assign V1259 = \V3(0)  & \V9(0) ;
  assign V1258 = \V9(0)  & \V2(0) ;
  assign n2607 = ~V778 & ~V780;
  assign n2608 = ~V787 & n2607;
  assign n2609 = ~V1258 & n2608;
  assign n2610 = ~V1259 & n2609;
  assign n2611 = ~V1263 & n2610;
  assign n2612 = ~V1387 & n2611;
  assign \V375(0)  = V1423 | ~n2612;
  assign n2614 = ~\V1536(0)  & ~n1711;
  assign n2615 = ~\V1536(0)  & ~n1229;
  assign n2616 = n691 & ~n2615;
  assign n2617 = ~n2614 & n2616;
  assign n2618 = \V1536(0)  & ~n2523;
  assign n2619 = ~\V1536(0)  & ~n2046;
  assign n2620 = n2617 & ~n2619;
  assign \V1512(1)  = n2618 | ~n2620;
  assign n2622 = n691 & \V1536(0) ;
  assign n2623 = ~\V1536(0)  & n1713;
  assign n2624 = ~\V1536(0)  & n1489;
  assign n2625 = ~\V1536(0)  & ~n1657;
  assign n2626 = ~\V1536(0)  & ~n1121;
  assign n2627 = ~\V1536(0)  & ~n1529;
  assign n2628 = ~\V1536(0)  & ~n1319;
  assign n2629 = ~\V1536(0)  & ~n1584;
  assign n2630 = ~\V1536(0)  & ~n1456;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = ~n2628 & n2631;
  assign n2633 = ~n2627 & n2632;
  assign n2634 = ~n2626 & n2633;
  assign n2635 = ~n2625 & n2634;
  assign n2636 = ~n2624 & n2635;
  assign n2637 = ~n2623 & n2636;
  assign \V1512(3)  = n2622 | ~n2637;
  assign n2639 = ~\V15(0)  & ~n867;
  assign \V410(0)  = n2150 | ~n2639;
  assign n2641 = ~\V1536(0)  & ~n2047;
  assign n2642 = ~n694 & \V1536(0) ;
  assign n2643 = n2617 & ~n2642;
  assign \V1512(2)  = n2641 | ~n2643;
  assign V1256 = \V2(0)  & n2520;
  assign n2646 = ~\V35(0)  & ~\V174(0) ;
  assign n2647 = \V12(0)  & n2646;
  assign n2648 = \V2(0)  & n2647;
  assign n2649 = \V57(0)  & n2648;
  assign n2650 = ~V707 & n2649;
  assign n2651 = ~n545 & n2650;
  assign n2652 = ~n547 & n2651;
  assign n2653 = ~n560 & n2652;
  assign n2654 = n554 & n2653;
  assign n2655 = ~\V57(0)  & n2648;
  assign n2656 = ~n783 & n2655;
  assign n2657 = ~n560 & n2656;
  assign n2658 = ~\V60(0)  & n2648;
  assign n2659 = ~\V63(0)  & n2658;
  assign n2660 = n560 & n2659;
  assign n2661 = ~n2657 & ~n2660;
  assign V1257 = n2654 | ~n2661;
  assign n2663 = \V101(0)  & \V14(0) ;
  assign n2664 = ~n2586 & n2663;
  assign n2665 = ~n502 & n2587;
  assign \V1759(0)  = n2664 | n2665;
  assign V1260 = \V3(0)  & \V11(0) ;
  assign V1261 = ~\V62(0)  & V1260;
  assign V1262 = \V4(0)  & n2520;
  assign V1264 = \V12(0)  & \V4(0) ;
  assign V1265 = \V52(0)  & V1264;
  assign V1266 = \V4(0)  & \V11(0) ;
  assign V1267 = \V2(0)  & \V11(0) ;
  assign n2674 = ~\V802(0)  & n551;
  assign n2675 = ~n810 & \V1243(9) ;
  assign n2676 = ~\V239(4)  & n2674;
  assign \V1552(1)  = n2675 | n2676;
  assign n2678 = \V423(0)  & ~\V393(0) ;
  assign n2679 = ~n1912 & n2678;
  assign n2680 = ~n1909 & n2679;
  assign \V398(0)  = ~n1903 | ~n2680;
  assign n2682 = ~\V239(3)  & \V239(4) ;
  assign n2683 = n2674 & n2682;
  assign n2684 = \V239(3)  & ~\V239(4) ;
  assign n2685 = n2674 & n2684;
  assign n2686 = ~n810 & \V1243(8) ;
  assign n2687 = ~n2685 & ~n2686;
  assign \V1552(0)  = n2683 | ~n2687;
  assign n2689 = n527 & ~n660;
  assign n2690 = n1998 & n2689;
  assign n2691 = n2218 & n2690;
  assign V1365 = n2561 & n2691;
  assign n2693 = ~\V268(0)  & n1866;
  assign n2694 = \V268(0)  & ~n1866;
  assign V1370 = n2693 | n2694;
  assign n2696 = \V268(3)  & ~n1863;
  assign n2697 = ~\V268(3)  & n1863;
  assign V1373 = n2696 | n2697;
  assign n2699 = \V268(3)  & ~V1373;
  assign n2700 = \V268(2)  & ~n2699;
  assign n2701 = ~\V268(2)  & n2699;
  assign V1372 = n2700 | n2701;
  assign n2703 = \V268(2)  & ~V1372;
  assign n2704 = ~n1866 & n2703;
  assign n2705 = \V268(1)  & ~n1866;
  assign V1371 = n2704 | n2705;
  assign n2707 = \V59(0)  & n1991;
  assign n2708 = \V56(0)  & ~n1749;
  assign n2709 = n2383 & ~n2708;
  assign \V508(0)  = n2707 | ~n2709;
  assign n2711 = ~\V268(5)  & \V268(4) ;
  assign n2712 = \V268(5)  & ~\V268(4) ;
  assign V1374 = n2711 | n2712;
  assign V1378 = ~n2289 & V782;
  assign n2715 = ~\V248(0)  & V782;
  assign n2716 = ~n2297 & n2715;
  assign n2717 = ~n906 & n2716;
  assign n2718 = ~n654 & n2717;
  assign n2719 = n2295 & V782;
  assign n2720 = ~V1378 & ~n2719;
  assign V1380 = n2718 | ~n2720;
  assign n2722 = ~n810 & V782;
  assign n2723 = n551 & V782;
  assign V1382 = n2722 | n2723;
  assign n2725 = \V56(0)  & V782;
  assign n2726 = n861 & n2725;
  assign n2727 = ~n867 & n2726;
  assign V1384 = n785 & n2727;
  assign V1386 = n1869 & V782;
  assign n2730 = ~\V294(0)  & ~n1748;
  assign n2731 = ~n2376 & n2730;
  assign n2732 = \V62(0)  & \V91(1) ;
  assign n2733 = n783 & n2732;
  assign n2734 = \V59(0)  & \V91(0) ;
  assign n2735 = n783 & n2734;
  assign n2736 = ~n2400 & ~n2735;
  assign n2737 = ~n2733 & n2736;
  assign \V1629(0)  = n2731 | ~n2737;
  assign n2739 = \V59(0)  & ~V1719;
  assign n2740 = n698 & n2739;
  assign n2741 = ~n920 & n2740;
  assign n2742 = ~n1724 & n2741;
  assign n2743 = ~n656 & n2742;
  assign n2744 = n2111 & n2743;
  assign n2745 = n2560 & n2744;
  assign n2746 = \V59(0)  & \V174(0) ;
  assign n2747 = ~V1719 & n2746;
  assign n2748 = n698 & n2747;
  assign n2749 = ~n920 & n2748;
  assign n2750 = ~n656 & n2749;
  assign n2751 = n2111 & n2750;
  assign n2752 = n2560 & n2751;
  assign n2753 = n1991 & n2561;
  assign n2754 = ~n2752 & ~n2753;
  assign \V1274(0)  = n2745 | ~n2754;
  assign V1426 = \V1(0)  & n2520;
  assign V1428 = \V1(0)  & \V11(0) ;
  assign V1429 = \V1(0)  & \V12(0) ;
  assign n2759 = ~\V109(0)  & V1423;
  assign n2760 = \V13(0)  & V1423;
  assign V1431 = n2759 | n2760;
  assign V1432 = \V66(0)  & n2111;
  assign n2763 = ~\V279(0)  & ~\V280(0) ;
  assign n2764 = ~n1992 & n2763;
  assign n2765 = \V279(0)  & \V280(0) ;
  assign n2766 = ~n1992 & n2765;
  assign n2767 = \V149(4)  & n1992;
  assign n2768 = ~n2766 & ~n2767;
  assign \V826(0)  = n2764 | ~n2768;
  assign n2770 = \V67(0)  & ~n1977;
  assign V1470 = n2111 & n2770;
  assign \V435(0)  = V432 | V630;
  assign V1537 = \V68(0)  & n2111;
  assign n2774 = \V50(0)  & n2111;
  assign n2775 = \V69(0)  & n2111;
  assign V1539 = n2774 | n2775;
  assign n2777 = ~\V16(0)  & \V15(0) ;
  assign \V1758(0)  = n2587 | n2777;
  assign n2779 = \V14(0)  & \V110(0) ;
  assign n2780 = ~n1736 & n2779;
  assign n2781 = ~n2777 & n2780;
  assign n2782 = \V110(0)  & n1888;
  assign n2783 = ~n2777 & n2782;
  assign n2784 = \V14(0)  & \V108(4) ;
  assign n2785 = \V110(0)  & n2784;
  assign n2786 = ~n1736 & n2785;
  assign n2787 = ~\V101(0)  & \V14(0) ;
  assign n2788 = \V110(0)  & n2787;
  assign n2789 = ~n1736 & n2788;
  assign n2790 = \V108(4)  & n1888;
  assign n2791 = \V110(0)  & n2790;
  assign n2792 = ~\V101(0)  & n1888;
  assign n2793 = \V110(0)  & n2792;
  assign n2794 = ~\V110(0)  & \V1758(0) ;
  assign n2795 = n501 & n2794;
  assign n2796 = \V102(0)  & ~\V110(0) ;
  assign n2797 = n501 & n2796;
  assign n2798 = ~n2795 & ~n2797;
  assign n2799 = ~n2793 & n2798;
  assign n2800 = ~n2791 & n2799;
  assign n2801 = ~n2789 & n2800;
  assign n2802 = ~n2786 & n2801;
  assign n2803 = ~n2783 & n2802;
  assign \V1968(0)  = n2781 | ~n2803;
  assign n2805 = \V213(2)  & ~n2356;
  assign n2806 = \V165(4)  & n2352;
  assign \V1297(1)  = n2805 | n2806;
  assign n2808 = \V213(1)  & ~n2356;
  assign n2809 = \V165(3)  & n2352;
  assign \V1297(0)  = n2808 | n2809;
  assign n2811 = \V213(4)  & ~n2356;
  assign n2812 = \V165(6)  & n2352;
  assign \V1297(3)  = n2811 | n2812;
  assign n2814 = \V213(3)  & ~n2356;
  assign n2815 = \V165(5)  & n2352;
  assign \V1297(2)  = n2814 | n2815;
  assign n2817 = \V213(5)  & ~n2356;
  assign n2818 = \V165(7)  & n2352;
  assign \V1297(4)  = n2817 | n2818;
  assign n2820 = \V274(0)  & ~\V202(0) ;
  assign \V640(0)  = \V271(0)  | n2820;
  assign n2822 = ~\V802(0)  & n1904;
  assign n2823 = \V14(0)  & \V262(0) ;
  assign n2824 = ~n2223 & n2823;
  assign \V1679(0)  = ~n526 | n2824;
  assign n2826 = ~n785 & ~\V1679(0) ;
  assign n2827 = ~n1736 & n2826;
  assign n2828 = ~n2224 & n2827;
  assign n2829 = n2220 & n2828;
  assign n2830 = ~\V1741(0)  & n2829;
  assign n2831 = ~n1978 & n2830;
  assign n2832 = ~n2822 & n2831;
  assign n2833 = n1976 & n2832;
  assign n2834 = ~n2238 & ~n2829;
  assign n2835 = ~n1978 & n2834;
  assign n2836 = ~n2822 & n2835;
  assign n2837 = ~n691 & ~n2829;
  assign n2838 = ~n1978 & n2837;
  assign n2839 = ~n2822 & n2838;
  assign n2840 = ~n1978 & n2243;
  assign n2841 = ~n2822 & n2840;
  assign n2842 = ~n691 & ~\V1741(0) ;
  assign n2843 = ~n1978 & n2842;
  assign n2844 = ~n2822 & n2843;
  assign n2845 = \V289(0)  & ~n1978;
  assign n2846 = ~\V1741(0)  & n2242;
  assign n2847 = ~n1978 & n2846;
  assign n2848 = ~n2845 & ~n2847;
  assign n2849 = ~n2844 & n2848;
  assign n2850 = ~n2841 & n2849;
  assign n2851 = ~n2839 & n2850;
  assign n2852 = ~n2836 & n2851;
  assign V1669 = n2833 | ~n2852;
  assign n2854 = ~\V290(0)  & ~\V289(0) ;
  assign n2855 = ~n653 & n2854;
  assign V1736 = n2822 & n2855;
  assign n2857 = \V14(0)  & \V261(0) ;
  assign n2858 = n1868 & n2857;
  assign n2859 = ~n2223 & n2857;
  assign n2860 = \V14(0)  & \V268(0) ;
  assign n2861 = n1866 & n2860;
  assign n2862 = ~\V262(0)  & n2857;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = ~n2859 & n2863;
  assign V1832 = n2858 | ~n2864;
  assign n2866 = \V108(1)  & ~n1731;
  assign n2867 = n547 & ~n861;
  assign \V1897(0)  = n2866 | n2867;
  assign n2869 = ~n550 & ~n651;
  assign n2870 = ~\V249(0)  & ~\V289(0) ;
  assign n2871 = ~\V290(0)  & n2870;
  assign n2872 = \V295(0)  & n2871;
  assign n2873 = n527 & n2872;
  assign \V1652(0)  = n2869 | ~n2873;
  assign n2875 = n501 & n665;
  assign n2876 = \V108(3)  & ~n1731;
  assign \V1899(0)  = n2875 | n2876;
  assign n2878 = \V258(0)  & \V14(0) ;
  assign n2879 = n1873 & n2878;
  assign n2880 = ~n1869 & n2879;
  assign n2881 = ~\V258(0)  & \V14(0) ;
  assign n2882 = ~n1873 & n2881;
  assign n2883 = ~V1370 & n2881;
  assign n2884 = n1866 & n2883;
  assign n2885 = ~n2882 & ~n2884;
  assign \V1451(0)  = n2880 | ~n2885;
  assign n2887 = \V37(0)  & ~\V1243(7) ;
  assign n2888 = ~\V37(0)  & ~\V1213(10) ;
  assign \V1829(7)  = n2887 | n2888;
  assign n2890 = \V37(0)  & ~\V1243(6) ;
  assign n2891 = ~\V37(0)  & ~\V1213(9) ;
  assign \V1829(6)  = n2890 | n2891;
  assign n2893 = ~\V37(0)  & \V321(2) ;
  assign n2894 = \V37(0)  & ~\V1243(9) ;
  assign \V1829(9)  = n2893 | n2894;
  assign n2896 = \V37(0)  & ~\V1243(8) ;
  assign n2897 = ~\V37(0)  & ~\V1213(11) ;
  assign \V1829(8)  = n2896 | n2897;
  assign n2899 = ~\V134(1)  & ~n560;
  assign n2900 = ~\V88(3)  & n560;
  assign \V1771(1)  = n2899 | n2900;
  assign n2902 = \V174(0)  & ~n691;
  assign n2903 = \V174(0)  & n867;
  assign n2904 = ~\V302(0)  & \V292(0) ;
  assign n2905 = ~n490 & ~n2904;
  assign n2906 = ~n2903 & n2905;
  assign \V1620(0)  = n2902 | ~n2906;
  assign n2908 = ~\V134(0)  & ~n560;
  assign n2909 = ~\V88(2)  & n560;
  assign \V1771(0)  = n2908 | n2909;
  assign n2911 = \V37(0)  & ~\V1243(1) ;
  assign n2912 = ~\V37(0)  & ~\V1213(4) ;
  assign \V1829(1)  = n2911 | n2912;
  assign n2914 = \V37(0)  & ~\V1213(2) ;
  assign \V1829(0)  = n2893 | n2914;
  assign n2916 = \V37(0)  & ~\V1243(3) ;
  assign n2917 = ~\V37(0)  & ~\V1213(6) ;
  assign \V1829(3)  = n2916 | n2917;
  assign n2919 = \V37(0)  & ~\V1243(2) ;
  assign n2920 = ~\V37(0)  & ~\V1213(5) ;
  assign \V1829(2)  = n2919 | n2920;
  assign n2922 = \V37(0)  & ~\V1243(5) ;
  assign n2923 = ~\V37(0)  & ~\V1213(8) ;
  assign \V1829(5)  = n2922 | n2923;
  assign n2925 = \V37(0)  & ~\V1243(4) ;
  assign n2926 = ~\V37(0)  & ~\V1213(7) ;
  assign \V1829(4)  = n2925 | n2926;
  assign n2928 = \V108(4)  & ~n1731;
  assign \V1900(0)  = n2777 | n2928;
  assign n2930 = \V14(0)  & ~\V259(0) ;
  assign n2931 = ~n1873 & n2930;
  assign n2932 = \V14(0)  & \V259(0) ;
  assign n2933 = n1873 & n2932;
  assign \V1459(0)  = n2931 | n2933;
  assign n2935 = \V149(5)  & n1992;
  assign n2936 = ~\V279(0)  & ~n1992;
  assign \V821(0)  = n2935 | n2936;
  assign n2938 = \V149(7)  & \V802(0) ;
  assign n2939 = n540 & n2938;
  assign n2940 = n1990 & n2439;
  assign \V1645(0)  = n2939 | ~n2940;
  assign \V1833(0)  = ~\V261(0) ;
  assign \V585(0)  = ~\V34(0) ;
  assign \V1760(0)  = ~\V101(0) ;
  assign \V1243(0)  = ~\V321(2) ;
  assign V657 = ~\V257(7) ;
  assign \V1864(0)  = ~\V302(0) ;
  assign V1375 = ~\V268(5) ;
  assign \V1481(0)  = ~\V214(0) ;
  assign \V1671(0)  = ~\V205(0) ;
  assign \V1863(0)  = ~\V301(0) ;
  assign \V1495(0)  = ~\V175(0) ;
  assign \V1757(0)  = \V15(0) ;
endmodule


