// Benchmark "TOP" written by ABC on Sun Apr 24 20:32:42 2016

module TOP ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_;
  wire n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n124, n125,
    n126, n127, n128, n129, n131, n132, n134, n135, n137, n139, n142, n143,
    n145, n146, n147, n149, n150, n152, n153, n156, n161, n164, n165, n169,
    n170, n172, n175, n178, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n466, n467, n468, n469, n470, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n551, n552, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n645, n646, n647, n648,
    n649, n650, n651, n652, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687,
    n689, n690, n691, n692, n693, n695, n696, n697, n698, n699, n700, n701,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n787, n788, n789, n790,
    n791, n792, n794, n795, n796, n797, n798, n799, n800, n801, n802, n804,
    n805, n806, n807, n808, n809, n810, n811, n813, n814, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n831,
    n832, n833, n834, n836, n837, n838, n839, n840, n841, n843, n844, n845;
  assign n72 = ~i_3_ & ~i_4_;
  assign n73 = ~i_5_ & n72;
  assign n74 = ~i_6_ & n73;
  assign n75 = i_0_ & i_2_;
  assign n76 = ~i_1_ & n75;
  assign n77 = n74 & n76;
  assign n78 = i_3_ & ~i_4_;
  assign n79 = ~i_5_ & n78;
  assign n80 = ~i_6_ & n79;
  assign n81 = i_0_ & i_1_;
  assign n82 = n80 & n81;
  assign n83 = ~n77 & ~n82;
  assign n84 = ~i_0_ & ~i_1_;
  assign n85 = ~i_2_ & n84;
  assign n86 = i_1_ & i_2_;
  assign n87 = ~i_0_ & n86;
  assign n88 = ~n85 & ~n87;
  assign n89 = i_1_ & ~i_2_;
  assign n90 = ~i_0_ & n89;
  assign n91 = ~n76 & ~n90;
  assign n92 = n88 & n91;
  assign n93 = n80 & ~n92;
  assign n94 = n83 & ~n93;
  assign n95 = ~i_7_ & ~n94;
  assign n96 = i_7_ & n77;
  assign n97 = ~i_0_ & ~i_2_;
  assign n98 = ~i_1_ & ~n97;
  assign n99 = ~n75 & n98;
  assign n100 = n80 & n99;
  assign n101 = i_7_ & n80;
  assign n102 = ~n90 & ~n98;
  assign n103 = n101 & n102;
  assign n104 = ~n100 & ~n103;
  assign n105 = ~n96 & n104;
  assign n106 = i_0_ & ~i_1_;
  assign n107 = ~i_2_ & n106;
  assign o_20_ = n74 & n107;
  assign n109 = ~i_3_ & n85;
  assign n110 = ~i_4_ & n109;
  assign n111 = ~i_5_ & n110;
  assign n112 = ~i_6_ & n111;
  assign n113 = ~o_20_ & ~n112;
  assign n114 = n90 & n101;
  assign n115 = n113 & ~n114;
  assign n116 = i_2_ & n84;
  assign n117 = ~i_1_ & ~n116;
  assign n118 = n74 & ~n117;
  assign n119 = n76 & n101;
  assign n120 = ~n118 & ~n119;
  assign n121 = n115 & n120;
  assign n122 = n105 & n121;
  assign o_0_ = n95 | ~n122;
  assign n124 = i_4_ & ~i_5_;
  assign n125 = ~i_6_ & n124;
  assign n126 = n113 & ~n125;
  assign n127 = ~n100 & ~n118;
  assign n128 = n126 & n127;
  assign n129 = ~i_7_ & ~n128;
  assign o_1_ = n95 | n129;
  assign n131 = ~i_6_ & ~i_7_;
  assign n132 = i_5_ & n72;
  assign o_2_ = n131 & n132;
  assign n134 = i_5_ & n78;
  assign n135 = ~i_6_ & n134;
  assign o_3_ = ~i_7_ & n135;
  assign n137 = i_6_ & ~i_7_;
  assign o_4_ = n79 & n137;
  assign n139 = i_5_ & n137;
  assign o_5_ = ~i_4_ & n139;
  assign o_6_ = n80 & n116;
  assign n142 = i_6_ & n90;
  assign n143 = n132 & n142;
  assign o_7_ = i_7_ & n143;
  assign n145 = i_6_ & i_7_;
  assign n146 = n132 & n145;
  assign n147 = i_2_ & n81;
  assign o_8_ = n146 & n147;
  assign n149 = i_6_ & n73;
  assign n150 = i_7_ & n149;
  assign o_9_ = n116 & n150;
  assign n152 = n87 & n146;
  assign n153 = n134 & n145;
  assign o_15_ = n87 & n153;
  assign o_10_ = n152 | o_15_;
  assign n156 = n89 & n146;
  assign o_11_ = i_0_ & n156;
  assign o_12_ = n76 & n146;
  assign o_13_ = n90 & n153;
  assign o_14_ = n107 & n153;
  assign n161 = ~i_2_ & n81;
  assign o_16_ = n153 & n161;
  assign o_17_ = n107 & n124;
  assign n164 = i_3_ & i_4_;
  assign n165 = n116 & n164;
  assign o_18_ = ~i_5_ & n165;
  assign o_19_ = i_4_ & n109;
  assign o_21_ = n80 & n107;
  assign n169 = n79 & n145;
  assign n170 = ~n150 & ~n169;
  assign o_22_ = n107 & ~n170;
  assign n172 = i_3_ & i_5_;
  assign o_23_ = n85 & n172;
  assign o_24_ = n111 & n137;
  assign n175 = n73 & n90;
  assign o_25_ = n137 & n175;
  assign o_26_ = n75 & n150;
  assign n178 = n73 & n87;
  assign o_27_ = n137 & n178;
  assign o_28_ = n76 & n169;
  assign o_29_ = i_7_ & n112;
  assign o_30_ = n147 & n150;
  assign n183 = ~i_3_ & i_4_;
  assign n184 = n147 & n183;
  assign n185 = n147 & n164;
  assign n186 = n79 & n147;
  assign n187 = ~o_4_ & ~n186;
  assign n188 = ~n185 & n187;
  assign n189 = ~n184 & n188;
  assign n190 = ~n131 & n132;
  assign n191 = ~n145 & n190;
  assign n192 = n147 & n191;
  assign n193 = n134 & n147;
  assign n194 = ~n192 & ~n193;
  assign n195 = n189 & n194;
  assign n196 = ~o_8_ & n195;
  assign n197 = i_5_ & n164;
  assign n198 = n161 & n197;
  assign n199 = ~n73 & ~o_2_;
  assign n200 = n147 & ~n199;
  assign n201 = ~n198 & ~n200;
  assign n202 = n196 & n201;
  assign n203 = ~n135 & ~n169;
  assign n204 = ~n80 & n203;
  assign n205 = n161 & ~n204;
  assign n206 = i_6_ & n134;
  assign n207 = i_3_ & n124;
  assign n208 = ~n206 & ~n207;
  assign n209 = n161 & ~n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = n202 & n210;
  assign n212 = ~o_4_ & ~o_28_;
  assign n213 = i_5_ & n183;
  assign n214 = ~n80 & ~n213;
  assign n215 = n76 & ~n214;
  assign n216 = n212 & ~n215;
  assign n217 = ~n146 & ~n183;
  assign n218 = n161 & ~n217;
  assign n219 = n74 & n161;
  assign n220 = n149 & n161;
  assign n221 = ~n191 & ~n220;
  assign n222 = ~o_2_ & n221;
  assign n223 = ~n219 & n222;
  assign n224 = ~n218 & n223;
  assign n225 = ~n131 & n134;
  assign n226 = ~n164 & ~n225;
  assign n227 = n76 & ~n226;
  assign n228 = n224 & ~n227;
  assign n229 = n216 & n228;
  assign n230 = n211 & n229;
  assign n231 = n84 & n169;
  assign n232 = i_2_ & n231;
  assign n233 = ~n80 & ~n183;
  assign n234 = n116 & ~n233;
  assign n235 = ~n232 & ~n234;
  assign n236 = n116 & n153;
  assign n237 = ~o_18_ & ~n236;
  assign n238 = n235 & n237;
  assign n239 = ~i_5_ & n183;
  assign n240 = n85 & n239;
  assign n241 = ~n110 & ~n240;
  assign n242 = ~o_2_ & ~n149;
  assign n243 = ~n191 & n242;
  assign n244 = n107 & ~n243;
  assign n245 = ~n146 & ~n239;
  assign n246 = n107 & ~n245;
  assign n247 = ~n244 & ~n246;
  assign n248 = n241 & n247;
  assign n249 = n238 & n248;
  assign n250 = n87 & n164;
  assign n251 = n90 & ~n226;
  assign n252 = ~o_3_ & ~n169;
  assign n253 = n90 & ~n252;
  assign n254 = ~n251 & ~n253;
  assign n255 = ~n250 & n254;
  assign n256 = ~n178 & n255;
  assign n257 = n249 & n256;
  assign n258 = i_3_ & ~n80;
  assign n259 = n90 & ~n258;
  assign n260 = ~i_2_ & n231;
  assign n261 = ~i_3_ & n116;
  assign n262 = n124 & n261;
  assign n263 = ~i_4_ & n261;
  assign n264 = n85 & ~n226;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n262 & n265;
  assign n267 = ~n260 & n266;
  assign n268 = n80 & n85;
  assign n269 = n267 & ~n268;
  assign n270 = ~n259 & n269;
  assign n271 = n87 & n206;
  assign n272 = n87 & ~n252;
  assign n273 = i_7_ & n135;
  assign n274 = n87 & n273;
  assign n275 = n87 & ~n214;
  assign n276 = ~n274 & ~n275;
  assign n277 = ~n272 & n276;
  assign n278 = n87 & ~n245;
  assign n279 = n277 & ~n278;
  assign n280 = ~n271 & n279;
  assign n281 = ~n150 & n245;
  assign n282 = n76 & ~n281;
  assign n283 = n107 & n169;
  assign n284 = i_7_ & ~n107;
  assign n285 = n206 & ~n284;
  assign n286 = n73 & ~n145;
  assign n287 = n76 & n286;
  assign n288 = ~n285 & ~n287;
  assign n289 = ~n135 & n288;
  assign n290 = ~n283 & n289;
  assign n291 = ~o_17_ & n290;
  assign n292 = ~n282 & n291;
  assign n293 = n280 & n292;
  assign n294 = n270 & n293;
  assign n295 = n257 & n294;
  assign o_31_ = ~n230 | ~n295;
  assign n297 = n85 & ~n203;
  assign n298 = n230 & ~n297;
  assign n299 = i_5_ & n110;
  assign n300 = ~o_19_ & ~n268;
  assign n301 = ~n299 & n300;
  assign n302 = n298 & n301;
  assign n303 = n111 & ~n137;
  assign n304 = ~n175 & ~n303;
  assign n305 = ~n236 & n304;
  assign n306 = n90 & n169;
  assign n307 = ~n114 & ~n306;
  assign n308 = n79 & n131;
  assign n309 = ~n183 & ~n308;
  assign n310 = n90 & ~n309;
  assign n311 = n307 & ~n310;
  assign n312 = ~o_20_ & ~n274;
  assign n313 = n247 & n312;
  assign n314 = n80 & n87;
  assign n315 = n87 & n169;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~n164 & ~n206;
  assign n318 = n87 & ~n317;
  assign n319 = n316 & ~n318;
  assign n320 = ~n153 & ~n164;
  assign n321 = n90 & ~n320;
  assign n322 = ~n178 & ~n321;
  assign n323 = n87 & ~n217;
  assign n324 = n322 & ~n323;
  assign n325 = n319 & n324;
  assign n326 = n313 & n325;
  assign n327 = n311 & n326;
  assign n328 = n85 & ~n317;
  assign n329 = n235 & ~n263;
  assign n330 = ~n328 & n329;
  assign n331 = n327 & n330;
  assign n332 = n305 & n331;
  assign n333 = ~o_7_ & n292;
  assign n334 = n332 & n333;
  assign o_32_ = ~n302 | ~n334;
  assign n336 = n116 & n146;
  assign n337 = ~o_9_ & ~n336;
  assign n338 = ~n234 & n337;
  assign n339 = n116 & n286;
  assign n340 = n85 & ~n320;
  assign n341 = ~n339 & ~n340;
  assign n342 = n338 & n341;
  assign n343 = ~n260 & n342;
  assign n344 = n300 & n343;
  assign n345 = n87 & ~n199;
  assign n346 = n90 & n197;
  assign n347 = ~n345 & ~n346;
  assign n348 = n87 & n191;
  assign n349 = n347 & ~n348;
  assign n350 = ~n323 & n349;
  assign n351 = n90 & ~n214;
  assign n352 = n90 & n207;
  assign n353 = ~n351 & ~n352;
  assign n354 = n90 & n134;
  assign n355 = ~n306 & ~n354;
  assign n356 = n353 & n355;
  assign n357 = n350 & n356;
  assign n358 = ~n183 & ~n190;
  assign n359 = n76 & ~n358;
  assign n360 = ~n161 & ~n359;
  assign n361 = ~i_7_ & n314;
  assign n362 = n360 & ~n361;
  assign n363 = n147 & n286;
  assign n364 = n362 & ~n363;
  assign n365 = n357 & n364;
  assign n366 = n76 & n80;
  assign n367 = ~n107 & ~n366;
  assign n368 = n365 & n367;
  assign n369 = n344 & n368;
  assign n370 = n90 & ~n245;
  assign n371 = ~n175 & ~n370;
  assign n372 = ~n165 & n371;
  assign n373 = ~n232 & ~n236;
  assign n374 = n372 & n373;
  assign n375 = n289 & n374;
  assign n376 = n228 & n375;
  assign n377 = ~n87 & ~n110;
  assign n378 = n376 & n377;
  assign n379 = n189 & n378;
  assign o_33_ = ~n369 | ~n379;
  assign n381 = i_4_ & n87;
  assign n382 = ~n314 & ~n381;
  assign n383 = n107 & n286;
  assign n384 = n101 & n107;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~o_15_ & ~n278;
  assign n387 = n385 & n386;
  assign n388 = n382 & n387;
  assign n389 = ~n178 & ~n251;
  assign n390 = n311 & n389;
  assign n391 = n388 & n390;
  assign n392 = n107 & n197;
  assign n393 = n107 & n146;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n213 & n394;
  assign n396 = n338 & n395;
  assign n397 = ~n165 & ~n175;
  assign n398 = ~o_7_ & n397;
  assign n399 = ~n213 & ~n308;
  assign n400 = n107 & ~n399;
  assign n401 = n398 & ~n400;
  assign n402 = n396 & n401;
  assign n403 = n391 & n402;
  assign n404 = n161 & n225;
  assign n405 = n224 & ~n404;
  assign n406 = n85 & n286;
  assign n407 = n85 & ~n214;
  assign n408 = ~n406 & ~n407;
  assign n409 = n73 & n116;
  assign n410 = ~i_6_ & n409;
  assign n411 = ~n328 & ~n410;
  assign n412 = n408 & n411;
  assign n413 = ~n282 & n412;
  assign n414 = n405 & n413;
  assign n415 = n85 & n150;
  assign n416 = ~n260 & ~n315;
  assign n417 = ~n415 & n416;
  assign n418 = ~n240 & ~n299;
  assign n419 = n216 & n418;
  assign n420 = n417 & n419;
  assign n421 = n80 & n161;
  assign n422 = n76 & ~n320;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n186 & n423;
  assign n425 = i_4_ & n161;
  assign n426 = i_3_ & n425;
  assign n427 = n147 & ~n358;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n200 & n428;
  assign n430 = n161 & n169;
  assign n431 = n145 & n193;
  assign n432 = ~n185 & ~n431;
  assign n433 = ~n430 & n432;
  assign n434 = n429 & n433;
  assign n435 = n424 & n434;
  assign n436 = n420 & n435;
  assign n437 = n414 & n436;
  assign n438 = ~n273 & n288;
  assign n439 = n373 & n438;
  assign n440 = n437 & n439;
  assign o_34_ = ~n403 | ~n440;
  assign n442 = n350 & ~n361;
  assign n443 = ~o_21_ & ~n306;
  assign n444 = ~n87 & ~o_13_;
  assign n445 = ~n135 & ~n383;
  assign n446 = n444 & n445;
  assign n447 = n443 & n446;
  assign n448 = ~n282 & ~n287;
  assign n449 = ~o_22_ & n353;
  assign n450 = n448 & n449;
  assign n451 = n447 & n450;
  assign n452 = n442 & n451;
  assign n453 = n298 & n452;
  assign n454 = n116 & n134;
  assign n455 = ~n145 & n454;
  assign n456 = n330 & ~n455;
  assign n457 = n107 & n207;
  assign n458 = ~n285 & ~n457;
  assign n459 = ~n246 & n458;
  assign n460 = ~n268 & n459;
  assign n461 = n456 & n460;
  assign n462 = n237 & n371;
  assign n463 = n461 & n462;
  assign n464 = ~n110 & n463;
  assign o_35_ = ~n453 | ~n464;
  assign n466 = n374 & n396;
  assign n467 = ~n285 & n466;
  assign n468 = ~n109 & ~n268;
  assign n469 = n467 & n468;
  assign n470 = n411 & n469;
  assign o_36_ = ~n453 | ~n470;
  assign n472 = n76 & ~n242;
  assign n473 = ~n165 & ~n236;
  assign n474 = ~n472 & n473;
  assign n475 = ~n231 & n474;
  assign n476 = n76 & o_3_;
  assign n477 = ~n457 & ~n476;
  assign n478 = ~n119 & ~n259;
  assign n479 = n477 & n478;
  assign n480 = ~n455 & n479;
  assign n481 = n475 & n480;
  assign n482 = ~o_3_ & ~n359;
  assign n483 = n88 & n360;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n109 & ~n484;
  assign n486 = n481 & n485;
  assign n487 = n83 & ~n366;
  assign n488 = ~n268 & n487;
  assign n489 = ~i_7_ & ~n488;
  assign n490 = ~n145 & n193;
  assign n491 = n105 & ~n490;
  assign n492 = n266 & n491;
  assign n493 = ~n489 & n492;
  assign n494 = n486 & n493;
  assign n495 = n313 & n442;
  assign n496 = n99 & n213;
  assign n497 = ~n404 & ~n496;
  assign n498 = n145 & n186;
  assign n499 = n355 & ~n498;
  assign n500 = ~n87 & ~n106;
  assign n501 = n169 & ~n500;
  assign n502 = ~n352 & ~n501;
  assign n503 = ~n318 & n502;
  assign n504 = n499 & n503;
  assign n505 = ~n227 & n504;
  assign n506 = n497 & n505;
  assign n507 = n434 & n506;
  assign n508 = n495 & n507;
  assign o_37_ = ~n494 | ~n508;
  assign n510 = n254 & n349;
  assign n511 = n280 & n510;
  assign n512 = ~n259 & n511;
  assign n513 = n211 & n512;
  assign n514 = ~n282 & ~n303;
  assign n515 = n290 & n301;
  assign n516 = n514 & n515;
  assign n517 = n229 & n516;
  assign n518 = ~n132 & ~n149;
  assign n519 = n107 & ~n518;
  assign n520 = ~o_20_ & ~n519;
  assign n521 = ~n250 & n520;
  assign n522 = n342 & n521;
  assign n523 = ~n231 & ~n236;
  assign n524 = n522 & n523;
  assign n525 = n517 & n524;
  assign o_38_ = ~n513 | ~n525;
  assign n527 = n116 & ~n518;
  assign n528 = n437 & ~n527;
  assign n529 = n107 & n149;
  assign n530 = ~i_7_ & n529;
  assign n531 = ~n236 & ~n530;
  assign n532 = ~n152 & ~n271;
  assign n533 = n382 & n532;
  assign n534 = n531 & n533;
  assign n535 = ~o_20_ & n443;
  assign n536 = n235 & n535;
  assign n537 = ~n213 & n459;
  assign n538 = n536 & n537;
  assign n539 = n534 & n538;
  assign n540 = ~n321 & ~n351;
  assign n541 = n87 & n286;
  assign n542 = ~n273 & ~n541;
  assign n543 = n540 & n542;
  assign n544 = n87 & n150;
  assign n545 = n372 & ~n544;
  assign n546 = n543 & n545;
  assign n547 = ~n287 & ~n392;
  assign n548 = n546 & n547;
  assign n549 = n539 & n548;
  assign o_39_ = ~n528 | ~n549;
  assign n551 = ~n87 & ~n260;
  assign n552 = ~n268 & n551;
  assign n553 = n305 & n552;
  assign n554 = n365 & n553;
  assign n555 = n196 & n235;
  assign n556 = n85 & n146;
  assign n557 = ~n519 & ~n556;
  assign n558 = n266 & ~n370;
  assign n559 = n557 & n558;
  assign n560 = n555 & n559;
  assign n561 = ~n404 & ~n430;
  assign n562 = ~n227 & ~n476;
  assign n563 = n212 & ~n366;
  assign n564 = n562 & n563;
  assign n565 = ~n421 & n564;
  assign n566 = n224 & n565;
  assign n567 = n561 & n566;
  assign n568 = n560 & n567;
  assign n569 = n291 & n568;
  assign o_40_ = ~n554 | ~n569;
  assign n571 = n456 & ~n457;
  assign n572 = n474 & n571;
  assign n573 = ~n297 & n521;
  assign n574 = n468 & n564;
  assign n575 = n107 & ~n233;
  assign n576 = ~n77 & ~n359;
  assign n577 = ~n575 & n576;
  assign n578 = n574 & n577;
  assign n579 = n573 & n578;
  assign n580 = ~n283 & n579;
  assign n581 = n572 & n580;
  assign o_41_ = ~n513 | ~n581;
  assign n583 = ~n219 & n432;
  assign n584 = i_4_ & o_23_;
  assign n585 = ~n262 & ~n584;
  assign n586 = n89 & n169;
  assign n587 = ~n268 & ~n586;
  assign n588 = n585 & n587;
  assign n589 = n583 & n588;
  assign n590 = n342 & n589;
  assign n591 = ~n427 & ~n544;
  assign n592 = n221 & ~n232;
  assign n593 = n591 & n592;
  assign n594 = n107 & n190;
  assign n595 = n416 & ~n594;
  assign n596 = n187 & ~n363;
  assign n597 = n595 & n596;
  assign n598 = n593 & n597;
  assign n599 = n590 & n598;
  assign n600 = ~n392 & n448;
  assign n601 = ~o_30_ & n600;
  assign n602 = ~o_19_ & ~n556;
  assign n603 = ~n111 & n602;
  assign n604 = n458 & n603;
  assign n605 = n388 & n604;
  assign n606 = n601 & n605;
  assign n607 = n599 & n606;
  assign n608 = n107 & ~n309;
  assign n609 = ~n218 & ~n608;
  assign n610 = n543 & n609;
  assign n611 = n473 & n610;
  assign n612 = ~o_16_ & ~n215;
  assign n613 = n423 & n612;
  assign n614 = ~n426 & n613;
  assign n615 = n611 & n614;
  assign n616 = n371 & n615;
  assign o_42_ = ~n607 | ~n616;
  assign n618 = n89 & ~n233;
  assign n619 = n304 & ~n618;
  assign n620 = n85 & n190;
  assign n621 = ~n366 & ~n620;
  assign n622 = n161 & ~n317;
  assign n623 = ~n143 & ~n541;
  assign n624 = ~n622 & n623;
  assign n625 = n621 & n624;
  assign n626 = n438 & n625;
  assign n627 = n619 & n626;
  assign n628 = ~n251 & ~n359;
  assign n629 = n534 & n628;
  assign n630 = ~o_11_ & ~n422;
  assign n631 = n629 & n630;
  assign n632 = n627 & n631;
  assign o_43_ = ~n599 | ~n632;
  assign n634 = ~n135 & n458;
  assign n635 = ~n283 & n634;
  assign n636 = ~n575 & n635;
  assign n637 = n600 & n636;
  assign n638 = n230 & n637;
  assign n639 = n342 & n374;
  assign n640 = n357 & n639;
  assign n641 = n552 & n640;
  assign n642 = ~n110 & ~n519;
  assign n643 = n641 & n642;
  assign o_44_ = ~n638 | ~n643;
  assign n645 = ~o_10_ & n520;
  assign n646 = i_6_ & n178;
  assign n647 = n645 & ~n646;
  assign n648 = ~n406 & n639;
  assign n649 = n647 & n648;
  assign n650 = n301 & ~n315;
  assign n651 = ~n90 & n650;
  assign n652 = n649 & n651;
  assign o_45_ = ~n638 | ~n652;
  assign n654 = ~n165 & ~o_25_;
  assign n655 = ~n114 & n373;
  assign n656 = n654 & n655;
  assign n657 = ~n260 & n468;
  assign n658 = n90 & n308;
  assign n659 = ~o_7_ & ~n658;
  assign n660 = n657 & n659;
  assign n661 = n656 & n660;
  assign n662 = n522 & n661;
  assign n663 = n511 & n662;
  assign o_46_ = ~n638 | ~n663;
  assign n665 = n429 & n567;
  assign n666 = ~o_15_ & n188;
  assign n667 = n313 & n666;
  assign n668 = ~n272 & n667;
  assign n669 = n665 & n668;
  assign n670 = ~n197 & n214;
  assign n671 = n107 & ~n670;
  assign n672 = ~n472 & n576;
  assign n673 = n635 & n672;
  assign n674 = ~n671 & n673;
  assign n675 = n456 & n674;
  assign n676 = n418 & n473;
  assign n677 = n408 & n676;
  assign n678 = n675 & n677;
  assign n679 = n254 & ~n646;
  assign n680 = ~n152 & n679;
  assign n681 = ~n259 & n680;
  assign n682 = n678 & n681;
  assign o_47_ = ~n669 | ~n682;
  assign n684 = n473 & n573;
  assign n685 = n512 & n684;
  assign n686 = n638 & n685;
  assign n687 = n329 & n686;
  assign o_48_ = n109 | ~n687;
  assign n689 = ~n232 & n337;
  assign n690 = n137 & n409;
  assign n691 = ~n328 & ~n690;
  assign n692 = n468 & n691;
  assign n693 = n686 & n692;
  assign o_49_ = ~n689 | ~n693;
  assign n695 = n90 & n286;
  assign n696 = ~n370 & ~n695;
  assign n697 = n566 & n696;
  assign n698 = ~n209 & ~n351;
  assign n699 = n202 & n698;
  assign n700 = n326 & n699;
  assign n701 = n678 & n700;
  assign o_50_ = ~n697 | ~n701;
  assign n703 = n327 & n674;
  assign n704 = n147 & n149;
  assign n705 = ~n426 & ~n704;
  assign n706 = n222 & ~n430;
  assign n707 = ~o_16_ & n706;
  assign n708 = n705 & n707;
  assign n709 = n565 & n708;
  assign n710 = n703 & n709;
  assign n711 = n85 & n153;
  assign n712 = n603 & ~n711;
  assign n713 = ~i_5_ & ~n175;
  assign n714 = ~n398 & ~n713;
  assign n715 = n712 & ~n714;
  assign n716 = ~n231 & n237;
  assign n717 = n715 & n716;
  assign n718 = ~o_8_ & ~n498;
  assign n719 = ~n431 & n718;
  assign n720 = ~n261 & n719;
  assign n721 = n717 & n720;
  assign o_51_ = ~n710 | ~n721;
  assign n723 = n636 & ~n690;
  assign n724 = ~o_8_ & n187;
  assign n725 = n432 & n724;
  assign n726 = n705 & n725;
  assign n727 = n212 & n389;
  assign n728 = n521 & n727;
  assign n729 = n726 & n728;
  assign n730 = n280 & n729;
  assign n731 = n723 & n730;
  assign n732 = ~n190 & ~n308;
  assign n733 = n76 & ~n732;
  assign n734 = ~n392 & ~n733;
  assign n735 = n337 & n734;
  assign n736 = ~n253 & n735;
  assign n737 = ~o_11_ & ~n404;
  assign n738 = n423 & n737;
  assign n739 = n706 & n738;
  assign n740 = n712 & n739;
  assign n741 = n481 & n740;
  assign n742 = n736 & n741;
  assign o_52_ = ~n731 | ~n742;
  assign n744 = ~o_30_ & n561;
  assign n745 = n355 & ~n646;
  assign n746 = ~n363 & n745;
  assign n747 = n744 & n746;
  assign n748 = n637 & n747;
  assign n749 = n229 & n748;
  assign n750 = n312 & n749;
  assign n751 = ~n111 & n397;
  assign n752 = ~n232 & n751;
  assign n753 = n344 & n752;
  assign n754 = n90 & n183;
  assign n755 = ~n184 & ~n754;
  assign n756 = n319 & n718;
  assign n757 = ~n152 & ~n244;
  assign n758 = n756 & n757;
  assign n759 = n755 & n758;
  assign n760 = n753 & n759;
  assign o_53_ = ~n750 | ~n760;
  assign n762 = ~n106 & n289;
  assign n763 = n659 & n762;
  assign n764 = n73 & n147;
  assign n765 = n347 & ~n764;
  assign n766 = ~n425 & n765;
  assign n767 = n763 & n766;
  assign n768 = n97 & n207;
  assign n769 = ~i_3_ & n381;
  assign n770 = ~n409 & ~n584;
  assign n771 = ~n769 & n770;
  assign n772 = ~n114 & n771;
  assign n773 = n195 & n772;
  assign n774 = ~n768 & n773;
  assign n775 = i_6_ & n175;
  assign n776 = n235 & ~n775;
  assign n777 = ~n315 & n473;
  assign n778 = n776 & n777;
  assign n779 = ~n297 & n468;
  assign n780 = n778 & n779;
  assign n781 = n774 & n780;
  assign n782 = ~n421 & n561;
  assign n783 = n223 & n782;
  assign n784 = ~n253 & n783;
  assign n785 = n781 & n784;
  assign o_54_ = ~n767 | ~n785;
  assign n787 = ~o_7_ & n749;
  assign n788 = n189 & n778;
  assign n789 = n645 & n788;
  assign n790 = n267 & ~n407;
  assign n791 = n603 & n790;
  assign n792 = n789 & n791;
  assign o_55_ = ~n787 | ~n792;
  assign n794 = n238 & ~n714;
  assign n795 = n316 & ~n345;
  assign n796 = ~o_13_ & ~n754;
  assign n797 = ~n340 & n796;
  assign n798 = n795 & n797;
  assign n799 = n657 & n771;
  assign n800 = n798 & n799;
  assign n801 = n794 & n800;
  assign n802 = n521 & n801;
  assign o_56_ = ~n638 | ~n802;
  assign n804 = n277 & ~n764;
  assign n805 = n322 & n804;
  assign n806 = n555 & n805;
  assign n807 = n791 & n806;
  assign n808 = n307 & ~n381;
  assign n809 = n654 & n763;
  assign n810 = n405 & n809;
  assign n811 = n808 & n810;
  assign o_57_ = ~n807 | ~n811;
  assign n813 = n468 & n640;
  assign n814 = n674 & n813;
  assign o_58_ = ~n669 | ~n814;
  assign n816 = ~o_7_ & n602;
  assign n817 = n74 & n90;
  assign n818 = ~n336 & ~n817;
  assign n819 = n547 & n818;
  assign n820 = n816 & n819;
  assign n821 = ~n234 & ~n421;
  assign n822 = ~n153 & ~n213;
  assign n823 = n76 & ~n822;
  assign n824 = ~n310 & ~n823;
  assign n825 = n821 & n824;
  assign n826 = n820 & n825;
  assign n827 = n656 & n826;
  assign n828 = n414 & n827;
  assign o_59_ = ~n731 | ~n828;
  assign n830 = n74 & n147;
  assign n831 = n724 & ~n830;
  assign n832 = n583 & n831;
  assign n833 = ~n156 & n832;
  assign n834 = n753 & n833;
  assign o_60_ = ~n710 | ~n834;
  assign n836 = n212 & ~n823;
  assign n837 = n794 & n836;
  assign n838 = n790 & n837;
  assign n839 = n224 & n241;
  assign n840 = n838 & n839;
  assign n841 = n703 & n840;
  assign o_61_ = ~n211 | ~n841;
  assign n843 = n726 & n739;
  assign n844 = n762 & n843;
  assign n845 = n551 & n844;
  assign o_62_ = ~n813 | ~n845;
endmodule


