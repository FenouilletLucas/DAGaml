// Benchmark "i5" written by ABC on Tue May 16 16:07:50 2017

module i5 ( 
    \V124(2) , \V40(3) , \V88(11) , \V40(5) , \V88(10) , \V40(6) ,
    \V40(7) , \V124(1) , \V40(9) , \V112(3) , \V112(2) , \V112(1) ,
    \V40(13) , \V40(15) , \V40(14) , \V100(3) , \V100(2) , \V100(5) ,
    \V40(11) , \V40(10) , \V128(3) , \V100(1) , \V128(2) , \V115(3) ,
    \V115(2) , \V128(1) , \V100(7) , \V128(0) , \V76(13) , \V100(6) ,
    \V100(9) , \V76(15) , \V115(1) , \V76(14) , \V76(11) , \V103(3) ,
    \V76(10) , \V103(2) , \V103(1) , \V2(0) , \V2(1) , \V118(3) ,
    \V118(2) , \V118(1) , \V106(3) , \V4(0) , \V106(2) , \V100(11) ,
    \V4(1) , \V100(10) , \V100(13) , \V100(15) , \V106(1) , \V100(14) ,
    \V28(13) , \V28(15) , \V28(14) , \V64(13) , \V28(11) , \V64(15) ,
    \V28(10) , \V64(14) , \V64(11) , \V64(10) , \V109(3) , \V109(2) ,
    \V109(1) , \V88(1) , \V88(2) , \V88(3) , \V88(5) , \V88(6) , \V132(3) ,
    \V88(7) , \V132(2) , \V88(9) , \V76(1) , \V76(2) , \V132(1) , \V28(1) ,
    \V76(3) , \V132(0) , \V28(2) , \V28(3) , \V76(5) , \V76(6) , \V28(5) ,
    \V76(7) , \V28(6) , \V16(13) , \V28(7) , \V76(9) , \V133(0) ,
    \V16(15) , \V28(9) , \V64(1) , \V16(14) , \V64(2) , \V52(13) ,
    \V121(3) , \V16(1) , \V64(3) , \V121(2) , \V16(2) , \V16(11) ,
    \V52(15) , \V16(3) , \V64(5) , \V16(10) , \V52(14) , \V64(6) ,
    \V16(5) , \V64(7) , \V16(6) , \V52(11) , \V121(1) , \V16(7) , \V64(9) ,
    \V52(10) , \V16(9) , \V52(1) , \V52(2) , \V52(3) , \V52(5) , \V52(6) ,
    \V52(7) , \V88(13) , \V52(9) , \V88(15) , \V40(1) , \V88(14) ,
    \V124(3) , \V40(2) ,
    \V199(1) , \V199(0) , \V199(7) , \V199(6) , \V199(9) , \V199(8) ,
    \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) , \V151(0) ,
    \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V167(3) , \V167(2) ,
    \V167(5) , \V167(4) , \V167(1) , \V167(0) , \V199(11) , \V167(7) ,
    \V199(10) , \V167(6) , \V199(13) , \V183(11) , \V167(9) , \V199(12) ,
    \V183(10) , \V167(8) , \V199(15) , \V183(13) , \V199(14) , \V183(12) ,
    \V183(15) , \V183(14) , \V167(11) , \V167(10) , \V167(13) , \V151(11) ,
    \V167(12) , \V151(10) , \V167(15) , \V151(13) , \V167(14) , \V151(12) ,
    \V151(15) , \V151(14) , \V183(3) , \V183(2) , \V183(5) , \V183(4) ,
    \V183(1) , \V183(0) , \V135(1) , \V135(0) , \V183(7) , \V183(6) ,
    \V183(9) , \V183(8) , \V199(3) , \V199(2) , \V199(5) , \V199(4)   );
  input  \V124(2) , \V40(3) , \V88(11) , \V40(5) , \V88(10) , \V40(6) ,
    \V40(7) , \V124(1) , \V40(9) , \V112(3) , \V112(2) , \V112(1) ,
    \V40(13) , \V40(15) , \V40(14) , \V100(3) , \V100(2) , \V100(5) ,
    \V40(11) , \V40(10) , \V128(3) , \V100(1) , \V128(2) , \V115(3) ,
    \V115(2) , \V128(1) , \V100(7) , \V128(0) , \V76(13) , \V100(6) ,
    \V100(9) , \V76(15) , \V115(1) , \V76(14) , \V76(11) , \V103(3) ,
    \V76(10) , \V103(2) , \V103(1) , \V2(0) , \V2(1) , \V118(3) ,
    \V118(2) , \V118(1) , \V106(3) , \V4(0) , \V106(2) , \V100(11) ,
    \V4(1) , \V100(10) , \V100(13) , \V100(15) , \V106(1) , \V100(14) ,
    \V28(13) , \V28(15) , \V28(14) , \V64(13) , \V28(11) , \V64(15) ,
    \V28(10) , \V64(14) , \V64(11) , \V64(10) , \V109(3) , \V109(2) ,
    \V109(1) , \V88(1) , \V88(2) , \V88(3) , \V88(5) , \V88(6) , \V132(3) ,
    \V88(7) , \V132(2) , \V88(9) , \V76(1) , \V76(2) , \V132(1) , \V28(1) ,
    \V76(3) , \V132(0) , \V28(2) , \V28(3) , \V76(5) , \V76(6) , \V28(5) ,
    \V76(7) , \V28(6) , \V16(13) , \V28(7) , \V76(9) , \V133(0) ,
    \V16(15) , \V28(9) , \V64(1) , \V16(14) , \V64(2) , \V52(13) ,
    \V121(3) , \V16(1) , \V64(3) , \V121(2) , \V16(2) , \V16(11) ,
    \V52(15) , \V16(3) , \V64(5) , \V16(10) , \V52(14) , \V64(6) ,
    \V16(5) , \V64(7) , \V16(6) , \V52(11) , \V121(1) , \V16(7) , \V64(9) ,
    \V52(10) , \V16(9) , \V52(1) , \V52(2) , \V52(3) , \V52(5) , \V52(6) ,
    \V52(7) , \V88(13) , \V52(9) , \V88(15) , \V40(1) , \V88(14) ,
    \V124(3) , \V40(2) ;
  output \V199(1) , \V199(0) , \V199(7) , \V199(6) , \V199(9) , \V199(8) ,
    \V151(3) , \V151(2) , \V151(5) , \V151(4) , \V151(1) , \V151(0) ,
    \V151(7) , \V151(6) , \V151(9) , \V151(8) , \V167(3) , \V167(2) ,
    \V167(5) , \V167(4) , \V167(1) , \V167(0) , \V199(11) , \V167(7) ,
    \V199(10) , \V167(6) , \V199(13) , \V183(11) , \V167(9) , \V199(12) ,
    \V183(10) , \V167(8) , \V199(15) , \V183(13) , \V199(14) , \V183(12) ,
    \V183(15) , \V183(14) , \V167(11) , \V167(10) , \V167(13) , \V151(11) ,
    \V167(12) , \V151(10) , \V167(15) , \V151(13) , \V167(14) , \V151(12) ,
    \V151(15) , \V151(14) , \V183(3) , \V183(2) , \V183(5) , \V183(4) ,
    \V183(1) , \V183(0) , \V135(1) , \V135(0) , \V183(7) , \V183(6) ,
    \V183(9) , \V183(8) , \V199(3) , \V199(2) , \V199(5) , \V199(4) ;
  wire n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n212, n213, n214, n215, n216, n218, n220, n221, n223, n225, n226, n227,
    n228, n230, n231, n232, n233, n235, n236, n237, n238, n239, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n253, n254, n255,
    n256, n257, n259, n261, n262, n263, n264, n266, n267, n268, n269, n270,
    n272, n273, n274, n275, n276, n278, n279, n280, n281, n282, n283, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n297, n299,
    n300, n302, n303, n304, n305, n307, n308, n309, n310, n311, n313, n314,
    n315, n316, n317, n319, n320, n321, n322, n323, n325, n327, n328, n329,
    n330, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342, n344,
    n345, n346, n347, n348, n349, n351, n353, n355, n356, n358, n359, n361,
    n362, n363, n364, n365, n366, n367, n368, n370, n372, n374, n375, n376,
    n377, n379, n380, n381, n382, n383, n385, n386, n387, n388, n390, n392,
    n393, n394, n395, n396, n397, n398, n399, n401, n402, n404, n406, n407,
    n409, n411, n412, n414, n415, n416, n417, n418, n419, n420, n421, n423,
    n425, n426, n428, n430, n431, n432, n433, n434, n435, n436, n437, n439,
    n440, n442, n444, n445, n447, n448, n449, n450, n451, n452, n453, n454,
    n456, n458, n459, n460, n461, n463, n464, n465, n466, n467, n469, n470,
    n471, n472, n473, n475, n476, n477, n478, n479, n480, n482, n484, n485,
    n486, n487, n489, n491, n492, n494, n495, n496, n497, n498, n499, n501,
    n503, n504, n506, n507, n508, n509, n510, n511;
  assign n200 = \V100(2)  & \V88(3) ;
  assign n201 = \V100(1)  & n200;
  assign n202 = \V100(1)  & \V88(2) ;
  assign n203 = \V124(2)  & \V121(3) ;
  assign n204 = \V124(1)  & n203;
  assign n205 = \V124(1)  & \V121(2) ;
  assign n206 = \V124(2)  & \V133(0) ;
  assign n207 = \V124(1)  & n206;
  assign n208 = \V124(3)  & n207;
  assign n209 = ~n205 & ~n208;
  assign n210 = ~\V121(1)  & n209;
  assign \V199(4)  = n204 | ~n210;
  assign n212 = \V100(2)  & \V199(4) ;
  assign n213 = \V100(1)  & n212;
  assign n214 = \V100(3)  & n213;
  assign n215 = ~n202 & ~n214;
  assign n216 = ~\V88(1)  & n215;
  assign \V199(1)  = n201 | ~n216;
  assign n218 = \V132(3)  & \V133(0) ;
  assign \V199(0)  = \V128(3)  | n218;
  assign n220 = \V124(3)  & n206;
  assign n221 = ~\V121(2)  & ~n220;
  assign \V199(8)  = n203 | ~n221;
  assign n223 = \V100(7)  & \V199(8) ;
  assign \V199(7)  = \V88(7)  | n223;
  assign n225 = \V100(6)  & \V88(7) ;
  assign n226 = \V100(6)  & \V199(8) ;
  assign n227 = \V100(7)  & n226;
  assign n228 = ~\V88(6)  & ~n227;
  assign \V199(6)  = n225 | ~n228;
  assign n230 = \V88(11)  & \V100(10) ;
  assign n231 = \V100(9)  & n230;
  assign n232 = \V88(10)  & \V100(9) ;
  assign n233 = \V133(0)  & \V124(3) ;
  assign \V199(12)  = \V121(3)  | n233;
  assign n235 = \V100(10)  & \V199(12) ;
  assign n236 = \V100(9)  & n235;
  assign n237 = \V100(11)  & n236;
  assign n238 = ~n232 & ~n237;
  assign n239 = ~\V88(9)  & n238;
  assign \V199(9)  = n231 | ~n239;
  assign n241 = \V103(3)  & \V106(2) ;
  assign n242 = \V106(1)  & n241;
  assign n243 = \V103(2)  & \V106(1) ;
  assign n244 = \V128(3)  & \V132(2) ;
  assign n245 = \V132(1)  & n244;
  assign n246 = \V128(2)  & \V132(1) ;
  assign n247 = \V132(2)  & \V133(0) ;
  assign n248 = \V132(1)  & n247;
  assign n249 = \V132(3)  & n248;
  assign n250 = ~n246 & ~n249;
  assign n251 = ~\V128(1)  & n250;
  assign \V167(0)  = n245 | ~n251;
  assign n253 = \V106(2)  & \V167(0) ;
  assign n254 = \V106(1)  & n253;
  assign n255 = \V106(3)  & n254;
  assign n256 = ~n243 & ~n255;
  assign n257 = ~\V103(1)  & n256;
  assign \V151(4)  = n242 | ~n257;
  assign n259 = \V28(3)  & \V151(4) ;
  assign \V151(3)  = \V16(3)  | n259;
  assign n261 = \V28(2)  & \V16(3) ;
  assign n262 = \V28(2)  & \V151(4) ;
  assign n263 = \V28(3)  & n262;
  assign n264 = ~\V16(2)  & ~n263;
  assign \V151(2)  = n261 | ~n264;
  assign n266 = \V28(6)  & \V16(7) ;
  assign n267 = \V28(5)  & n266;
  assign n268 = \V28(5)  & \V16(6) ;
  assign n269 = \V106(3)  & n253;
  assign n270 = ~\V103(2)  & ~n269;
  assign \V151(8)  = n241 | ~n270;
  assign n272 = \V28(6)  & \V151(8) ;
  assign n273 = \V28(5)  & n272;
  assign n274 = \V28(7)  & n273;
  assign n275 = ~n268 & ~n274;
  assign n276 = ~\V16(5)  & n275;
  assign \V151(5)  = n267 | ~n276;
  assign n278 = \V28(1)  & n261;
  assign n279 = \V28(1)  & \V16(2) ;
  assign n280 = \V28(1)  & n262;
  assign n281 = \V28(3)  & n280;
  assign n282 = ~n279 & ~n281;
  assign n283 = ~\V16(1)  & n282;
  assign \V151(1)  = n278 | ~n283;
  assign n285 = \V132(2)  & \V132(0) ;
  assign n286 = \V128(3)  & n285;
  assign n287 = \V132(1)  & n286;
  assign n288 = \V128(1)  & \V132(0) ;
  assign n289 = \V132(0)  & n246;
  assign n290 = \V132(0)  & n247;
  assign n291 = \V132(1)  & n290;
  assign n292 = \V132(3)  & n291;
  assign n293 = ~n289 & ~n292;
  assign n294 = ~\V128(0)  & n293;
  assign n295 = ~n288 & n294;
  assign \V151(0)  = n287 | ~n295;
  assign n297 = \V28(7)  & \V151(8) ;
  assign \V151(7)  = \V16(7)  | n297;
  assign n299 = \V28(7)  & n272;
  assign n300 = ~\V16(6)  & ~n299;
  assign \V151(6)  = n266 | ~n300;
  assign n302 = \V28(10)  & \V16(11) ;
  assign n303 = \V28(9)  & n302;
  assign n304 = \V28(9)  & \V16(10) ;
  assign n305 = \V106(3)  & \V167(0) ;
  assign \V151(12)  = \V103(3)  | n305;
  assign n307 = \V28(10)  & \V151(12) ;
  assign n308 = \V28(9)  & n307;
  assign n309 = \V28(11)  & n308;
  assign n310 = ~n304 & ~n309;
  assign n311 = ~\V16(9)  & n310;
  assign \V151(9)  = n303 | ~n311;
  assign n313 = \V112(2)  & \V109(3) ;
  assign n314 = \V112(1)  & n313;
  assign n315 = \V112(1)  & \V109(2) ;
  assign n316 = \V132(3)  & n247;
  assign n317 = ~\V128(2)  & ~n316;
  assign \V183(0)  = n244 | ~n317;
  assign n319 = \V112(2)  & \V183(0) ;
  assign n320 = \V112(1)  & n319;
  assign n321 = \V112(3)  & n320;
  assign n322 = ~n315 & ~n321;
  assign n323 = ~\V109(1)  & n322;
  assign \V167(4)  = n314 | ~n323;
  assign n325 = \V52(3)  & \V167(4) ;
  assign \V167(3)  = \V40(3)  | n325;
  assign n327 = \V40(3)  & \V52(2) ;
  assign n328 = \V52(2)  & \V167(4) ;
  assign n329 = \V52(3)  & n328;
  assign n330 = ~\V40(2)  & ~n329;
  assign \V167(2)  = n327 | ~n330;
  assign n332 = \V40(7)  & \V52(6) ;
  assign n333 = \V52(5)  & n332;
  assign n334 = \V40(6)  & \V52(5) ;
  assign n335 = \V112(3)  & n319;
  assign n336 = ~\V109(2)  & ~n335;
  assign \V167(8)  = n313 | ~n336;
  assign n338 = \V52(6)  & \V167(8) ;
  assign n339 = \V52(5)  & n338;
  assign n340 = \V52(7)  & n339;
  assign n341 = ~n334 & ~n340;
  assign n342 = ~\V40(5)  & n341;
  assign \V167(5)  = n333 | ~n342;
  assign n344 = \V52(1)  & n327;
  assign n345 = \V52(1)  & \V40(2) ;
  assign n346 = \V52(1)  & n328;
  assign n347 = \V52(3)  & n346;
  assign n348 = ~n345 & ~n347;
  assign n349 = ~\V40(1)  & n348;
  assign \V167(1)  = n344 | ~n349;
  assign n351 = \V100(11)  & \V199(12) ;
  assign \V199(11)  = \V88(11)  | n351;
  assign n353 = \V52(7)  & \V167(8) ;
  assign \V167(7)  = \V40(7)  | n353;
  assign n355 = \V100(11)  & n235;
  assign n356 = ~\V88(10)  & ~n355;
  assign \V199(10)  = n230 | ~n356;
  assign n358 = \V52(7)  & n338;
  assign n359 = ~\V40(6)  & ~n358;
  assign \V167(6)  = n332 | ~n359;
  assign n361 = \V100(14)  & \V88(15) ;
  assign n362 = \V100(13)  & n361;
  assign n363 = \V100(13)  & \V88(14) ;
  assign n364 = \V100(14)  & \V133(0) ;
  assign n365 = \V100(13)  & n364;
  assign n366 = \V100(15)  & n365;
  assign n367 = ~n363 & ~n366;
  assign n368 = ~\V88(13)  & n367;
  assign \V199(13)  = n362 | ~n368;
  assign n370 = \V118(3)  & \V199(0) ;
  assign \V183(12)  = \V115(3)  | n370;
  assign n372 = \V76(11)  & \V183(12) ;
  assign \V183(11)  = \V64(11)  | n372;
  assign n374 = \V40(11)  & \V52(10) ;
  assign n375 = \V52(9)  & n374;
  assign n376 = \V40(10)  & \V52(9) ;
  assign n377 = \V112(3)  & \V183(0) ;
  assign \V167(12)  = \V109(3)  | n377;
  assign n379 = \V52(10)  & \V167(12) ;
  assign n380 = \V52(9)  & n379;
  assign n381 = \V52(11)  & n380;
  assign n382 = ~n376 & ~n381;
  assign n383 = ~\V40(9)  & n382;
  assign \V167(9)  = n375 | ~n383;
  assign n385 = \V76(10)  & \V64(11) ;
  assign n386 = \V76(10)  & \V183(12) ;
  assign n387 = \V76(11)  & n386;
  assign n388 = ~\V64(10)  & ~n387;
  assign \V183(10)  = n385 | ~n388;
  assign n390 = \V100(15)  & \V133(0) ;
  assign \V199(15)  = \V88(15)  | n390;
  assign n392 = \V76(14)  & \V64(15) ;
  assign n393 = \V76(13)  & n392;
  assign n394 = \V76(13)  & \V64(14) ;
  assign n395 = \V76(14)  & \V199(0) ;
  assign n396 = \V76(13)  & n395;
  assign n397 = \V76(15)  & n396;
  assign n398 = ~n394 & ~n397;
  assign n399 = ~\V64(13)  & n398;
  assign \V183(13)  = n393 | ~n399;
  assign n401 = \V100(15)  & n364;
  assign n402 = ~\V88(14)  & ~n401;
  assign \V199(14)  = n361 | ~n402;
  assign n404 = \V76(15)  & \V199(0) ;
  assign \V183(15)  = \V64(15)  | n404;
  assign n406 = \V76(15)  & n395;
  assign n407 = ~\V64(14)  & ~n406;
  assign \V183(14)  = n392 | ~n407;
  assign n409 = \V52(11)  & \V167(12) ;
  assign \V167(11)  = \V40(11)  | n409;
  assign n411 = \V52(11)  & n379;
  assign n412 = ~\V40(10)  & ~n411;
  assign \V167(10)  = n374 | ~n412;
  assign n414 = \V40(15)  & \V52(14) ;
  assign n415 = \V52(13)  & n414;
  assign n416 = \V40(14)  & \V52(13) ;
  assign n417 = \V52(14)  & \V183(0) ;
  assign n418 = \V52(13)  & n417;
  assign n419 = \V52(15)  & n418;
  assign n420 = ~n416 & ~n419;
  assign n421 = ~\V40(13)  & n420;
  assign \V167(13)  = n415 | ~n421;
  assign n423 = \V28(11)  & \V151(12) ;
  assign \V151(11)  = \V16(11)  | n423;
  assign n425 = \V28(11)  & n307;
  assign n426 = ~\V16(10)  & ~n425;
  assign \V151(10)  = n302 | ~n426;
  assign n428 = \V52(15)  & \V183(0) ;
  assign \V167(15)  = \V40(15)  | n428;
  assign n430 = \V28(14)  & \V16(15) ;
  assign n431 = \V28(13)  & n430;
  assign n432 = \V28(13)  & \V16(14) ;
  assign n433 = \V28(14)  & \V167(0) ;
  assign n434 = \V28(13)  & n433;
  assign n435 = \V28(15)  & n434;
  assign n436 = ~n432 & ~n435;
  assign n437 = ~\V16(13)  & n436;
  assign \V151(13)  = n431 | ~n437;
  assign n439 = \V52(15)  & n417;
  assign n440 = ~\V40(14)  & ~n439;
  assign \V167(14)  = n414 | ~n440;
  assign n442 = \V28(15)  & \V167(0) ;
  assign \V151(15)  = \V16(15)  | n442;
  assign n444 = \V28(15)  & n433;
  assign n445 = ~\V16(14)  & ~n444;
  assign \V151(14)  = n430 | ~n445;
  assign n447 = \V115(3)  & \V118(2) ;
  assign n448 = \V118(1)  & n447;
  assign n449 = \V115(2)  & \V118(1) ;
  assign n450 = \V118(2)  & \V199(0) ;
  assign n451 = \V118(1)  & n450;
  assign n452 = \V118(3)  & n451;
  assign n453 = ~n449 & ~n452;
  assign n454 = ~\V115(1)  & n453;
  assign \V183(4)  = n448 | ~n454;
  assign n456 = \V76(3)  & \V183(4) ;
  assign \V183(3)  = \V64(3)  | n456;
  assign n458 = \V76(2)  & \V64(3) ;
  assign n459 = \V76(2)  & \V183(4) ;
  assign n460 = \V76(3)  & n459;
  assign n461 = ~\V64(2)  & ~n460;
  assign \V183(2)  = n458 | ~n461;
  assign n463 = \V76(6)  & \V64(7) ;
  assign n464 = \V76(5)  & n463;
  assign n465 = \V76(5)  & \V64(6) ;
  assign n466 = \V118(3)  & n450;
  assign n467 = ~\V115(2)  & ~n466;
  assign \V183(8)  = n447 | ~n467;
  assign n469 = \V76(6)  & \V183(8) ;
  assign n470 = \V76(5)  & n469;
  assign n471 = \V76(7)  & n470;
  assign n472 = ~n465 & ~n471;
  assign n473 = ~\V64(5)  & n472;
  assign \V183(5)  = n464 | ~n473;
  assign n475 = \V76(1)  & n458;
  assign n476 = \V76(1)  & \V64(2) ;
  assign n477 = \V76(1)  & n459;
  assign n478 = \V76(3)  & n477;
  assign n479 = ~n476 & ~n478;
  assign n480 = ~\V64(1)  & n479;
  assign \V183(1)  = n475 | ~n480;
  assign n482 = \V4(1)  & \V151(0) ;
  assign \V135(1)  = \V2(1)  | n482;
  assign n484 = \V2(1)  & \V4(0) ;
  assign n485 = \V4(0)  & \V151(0) ;
  assign n486 = \V4(1)  & n485;
  assign n487 = ~\V2(0)  & ~n486;
  assign \V135(0)  = n484 | ~n487;
  assign n489 = \V76(7)  & \V183(8) ;
  assign \V183(7)  = \V64(7)  | n489;
  assign n491 = \V76(7)  & n469;
  assign n492 = ~\V64(6)  & ~n491;
  assign \V183(6)  = n463 | ~n492;
  assign n494 = \V76(9)  & n385;
  assign n495 = \V64(10)  & \V76(9) ;
  assign n496 = \V76(9)  & n386;
  assign n497 = \V76(11)  & n496;
  assign n498 = ~n495 & ~n497;
  assign n499 = ~\V64(9)  & n498;
  assign \V183(9)  = n494 | ~n499;
  assign n501 = \V100(3)  & \V199(4) ;
  assign \V199(3)  = \V88(3)  | n501;
  assign n503 = \V100(3)  & n212;
  assign n504 = ~\V88(2)  & ~n503;
  assign \V199(2)  = n200 | ~n504;
  assign n506 = \V100(5)  & n225;
  assign n507 = \V100(5)  & \V88(6) ;
  assign n508 = \V100(5)  & n226;
  assign n509 = \V100(7)  & n508;
  assign n510 = ~n507 & ~n509;
  assign n511 = ~\V88(5)  & n510;
  assign \V199(5)  = n506 | ~n511;
endmodule


