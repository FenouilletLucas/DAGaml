// Benchmark "k2" written by ABC on Tue May 16 16:07:51 2017

module k2 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, r0, s0,
    z0, z1, a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1, h2,
    i1, i2, j1, j2, k1, k2, l1, l2, m1, n1, o1, p1, q1, r1, s1, t0, t1, u0,
    u1, v0, v1, w0, w1, x0, x1, y0, y1  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0, p0, q0, r0, s0;
  output z0, z1, a1, a2, b1, b2, c1, c2, d1, d2, e1, e2, f1, f2, g1, g2, h1,
    h2, i1, i2, j1, j2, k1, k2, l1, l2, m1, n1, o1, p1, q1, r1, s1, t0, t1,
    u0, u1, v0, v1, w0, w1, x0, x1, y0, y1;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n235, n236, n237, n238, n240, n241, n242,
    n243, n245, n246, n247, n248, n249, n250, n251, n252, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n368, n369, n370, n371, n372, n373, n374, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n471, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n744, n745, n746, n747, n748, n749, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n841, n842, n843, n844, n845, n846, n848, n849, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n936, n937, n938, n940, n942, n943, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n957, n958, n959;
  assign n92 = ~b0 & ~c0;
  assign n93 = s & t;
  assign n94 = u & ~v;
  assign n95 = n93 & n94;
  assign n96 = n92 & n95;
  assign n97 = d0 & e0;
  assign n98 = n96 & n97;
  assign n99 = a & ~f;
  assign n100 = n98 & n99;
  assign n101 = b0 & n95;
  assign n102 = ~d0 & ~e0;
  assign n103 = a & d;
  assign n104 = n102 & n103;
  assign n105 = n101 & n104;
  assign n106 = d0 & ~e0;
  assign n107 = ~s & n106;
  assign n108 = a & n107;
  assign n109 = x & ~c0;
  assign n110 = ~t & n94;
  assign n111 = n109 & n110;
  assign n112 = n108 & n111;
  assign n113 = ~d0 & e0;
  assign n114 = ~s & n113;
  assign n115 = ~d & n114;
  assign n116 = c & n115;
  assign n117 = ~u & ~v;
  assign n118 = ~t & n117;
  assign n119 = c0 & n118;
  assign n120 = a & n119;
  assign n121 = n116 & n120;
  assign n122 = ~n112 & ~n121;
  assign c1 = n105 | ~n122;
  assign n124 = ~n100 & ~c1;
  assign n125 = ~l & a0;
  assign n126 = c0 & n110;
  assign n127 = s & n126;
  assign n128 = a & n113;
  assign n129 = n93 & n117;
  assign n130 = c0 & n129;
  assign n131 = l & a0;
  assign n132 = w & c0;
  assign n133 = t & n94;
  assign n134 = n132 & n133;
  assign n135 = ~b0 & c0;
  assign n136 = n95 & n135;
  assign n137 = ~a & ~e;
  assign n138 = n106 & n137;
  assign n139 = n136 & n138;
  assign n140 = n108 & n134;
  assign n141 = ~n139 & ~n140;
  assign n142 = n128 & n130;
  assign n143 = n125 & n142;
  assign n144 = n128 & n131;
  assign n145 = n127 & n144;
  assign n146 = n127 & n128;
  assign n147 = n125 & n146;
  assign n148 = ~n143 & ~n145;
  assign n149 = n141 & n148;
  assign n150 = n130 & n144;
  assign n151 = n149 & ~n150;
  assign y1 = n147 | ~n151;
  assign n153 = ~f & ~p;
  assign n154 = n128 & n153;
  assign n155 = s & ~c0;
  assign n156 = ~t & v;
  assign n157 = u & n156;
  assign n158 = n155 & n157;
  assign n159 = ~l & n158;
  assign n160 = k & z;
  assign n161 = n114 & n157;
  assign n162 = a & n161;
  assign n163 = n159 & n160;
  assign n164 = n154 & n163;
  assign n165 = ~l & n160;
  assign n166 = n162 & n165;
  assign n167 = ~n164 & ~n166;
  assign n168 = n106 & n129;
  assign n169 = a & n168;
  assign n170 = n160 & n169;
  assign n171 = ~l & n170;
  assign n172 = l & n158;
  assign n173 = n154 & n160;
  assign n174 = n172 & n173;
  assign n175 = l & n160;
  assign n176 = n162 & n175;
  assign n177 = ~n174 & ~n176;
  assign n178 = ~n170 & n177;
  assign n179 = ~n171 & n178;
  assign a1 = ~n167 | ~n179;
  assign n181 = ~y1 & ~a1;
  assign n182 = n110 & n155;
  assign n183 = a0 & n106;
  assign n184 = r & n183;
  assign n185 = n182 & n184;
  assign n186 = a & ~c0;
  assign n187 = n129 & n186;
  assign n188 = n183 & n187;
  assign n189 = w & ~c0;
  assign n190 = n133 & n189;
  assign n191 = ~f & n190;
  assign n192 = n108 & n191;
  assign n193 = a & n185;
  assign n194 = ~n188 & ~n192;
  assign n195 = ~n193 & n194;
  assign n196 = n131 & n158;
  assign n197 = n154 & n196;
  assign n198 = n131 & n162;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~r & n182;
  assign n201 = a & n183;
  assign n202 = n200 & n201;
  assign n203 = w & n158;
  assign n204 = ~c & n115;
  assign n205 = n126 & n204;
  assign n206 = a & n205;
  assign n207 = ~c0 & n118;
  assign n208 = ~d & n207;
  assign n209 = ~f & n108;
  assign n210 = n208 & n209;
  assign n211 = t & v;
  assign n212 = n114 & n211;
  assign n213 = n189 & n212;
  assign n214 = u & n213;
  assign n215 = a & n153;
  assign i2 = n214 & n215;
  assign n217 = a0 & n159;
  assign n218 = n154 & n217;
  assign n219 = n154 & n203;
  assign n220 = n125 & n162;
  assign n221 = w & n162;
  assign n222 = ~n210 & ~i2;
  assign n223 = ~n206 & n222;
  assign n224 = ~n221 & n223;
  assign n225 = ~n220 & n224;
  assign n226 = ~n219 & n225;
  assign n227 = ~n218 & n226;
  assign n228 = w & n169;
  assign n229 = ~n145 & ~n228;
  assign n230 = ~n171 & n229;
  assign n231 = ~n143 & n230;
  assign n232 = n227 & n231;
  assign n233 = n167 & n232;
  assign b1 = ~n141 | ~n233;
  assign n235 = ~n202 & ~b1;
  assign n236 = n199 & n235;
  assign n237 = n195 & n236;
  assign n238 = n181 & n237;
  assign z0 = ~n124 | ~n238;
  assign n240 = ~o & n92;
  assign n241 = n102 & n240;
  assign n242 = ~m & ~n;
  assign n243 = v & n242;
  assign z1 = n241 & n243;
  assign n245 = e & n106;
  assign n246 = n136 & n245;
  assign n247 = f & n98;
  assign n248 = ~n246 & ~n247;
  assign n249 = n101 & n113;
  assign n250 = n97 & n136;
  assign n251 = ~n105 & ~n250;
  assign n252 = ~n249 & n251;
  assign a2 = ~n248 | ~n252;
  assign n254 = ~s & n102;
  assign n255 = ~j & n189;
  assign n256 = ~u & n156;
  assign n257 = n107 & n256;
  assign n258 = n255 & n257;
  assign n259 = ~m0 & n258;
  assign n260 = ~p0 & n259;
  assign n261 = ~q0 & n260;
  assign n262 = ~n0 & n261;
  assign n263 = n114 & n256;
  assign n264 = j & n189;
  assign n265 = n263 & n264;
  assign n266 = o0 & n262;
  assign n267 = h0 & n265;
  assign n268 = ~n266 & ~n267;
  assign n269 = s & c0;
  assign n270 = n102 & n256;
  assign n271 = n269 & n270;
  assign n272 = n268 & ~n271;
  assign n273 = ~c0 & n212;
  assign n274 = y & n273;
  assign n275 = n119 & n254;
  assign n276 = n134 & n254;
  assign n277 = n272 & ~n274;
  assign n278 = n126 & n254;
  assign n279 = n277 & ~n278;
  assign n280 = ~n276 & n279;
  assign n281 = ~n275 & n280;
  assign n282 = ~f0 & ~h0;
  assign n283 = ~s & n97;
  assign n284 = n0 & n282;
  assign n285 = n265 & n284;
  assign n286 = n189 & n256;
  assign n287 = n283 & n286;
  assign n288 = n0 & n261;
  assign n289 = ~n287 & ~n288;
  assign n290 = ~n285 & n289;
  assign n291 = p0 & n259;
  assign n292 = n290 & ~n291;
  assign n293 = ~o0 & n262;
  assign n294 = ~r0 & s0;
  assign n295 = n293 & n294;
  assign n296 = ~n0 & q0;
  assign n297 = n260 & n296;
  assign n298 = ~n295 & ~n297;
  assign n299 = m0 & n258;
  assign n300 = n292 & n298;
  assign n301 = ~n299 & n300;
  assign n302 = n155 & n256;
  assign n303 = u & n211;
  assign n304 = a0 & n97;
  assign n305 = n159 & n304;
  assign n306 = n189 & n283;
  assign n307 = n303 & n306;
  assign n308 = ~n305 & ~n307;
  assign n309 = z & n97;
  assign n310 = n159 & n309;
  assign n311 = n97 & n203;
  assign n312 = n97 & n302;
  assign n313 = n308 & ~n310;
  assign n314 = ~n312 & n313;
  assign n315 = ~n311 & n314;
  assign n316 = a0 & ~c0;
  assign n317 = n97 & n129;
  assign n318 = n316 & n317;
  assign n319 = n190 & n283;
  assign n320 = n207 & n283;
  assign n321 = ~n185 & ~n320;
  assign n322 = ~n319 & n321;
  assign n323 = ~n318 & n322;
  assign n324 = ~c0 & n110;
  assign n325 = n283 & n324;
  assign n326 = n323 & ~n325;
  assign n327 = d & n114;
  assign n328 = n134 & n204;
  assign n329 = n134 & n327;
  assign n330 = ~n328 & ~n329;
  assign n331 = r & a0;
  assign n332 = n102 & n331;
  assign n333 = n127 & n332;
  assign n334 = a0 & n102;
  assign n335 = n130 & n334;
  assign n336 = ~n333 & ~n335;
  assign n337 = ~n0 & n282;
  assign n338 = n265 & n337;
  assign n339 = f0 & n265;
  assign n340 = n113 & n136;
  assign n341 = r0 & ~s0;
  assign n342 = n293 & n341;
  assign n343 = n102 & n136;
  assign n344 = n107 & n211;
  assign n345 = c0 & n344;
  assign n346 = a & c0;
  assign n347 = n212 & n346;
  assign n348 = a0 & n273;
  assign n349 = n160 & n273;
  assign w0 = n348 | n349;
  assign n351 = ~y1 & ~w0;
  assign n352 = ~n347 & n351;
  assign n353 = ~n121 & n352;
  assign n354 = ~n206 & n353;
  assign n355 = ~n100 & n354;
  assign n356 = ~n345 & n355;
  assign n357 = ~n343 & n356;
  assign n358 = ~n342 & n357;
  assign n359 = ~n340 & n358;
  assign n360 = ~n339 & n359;
  assign n361 = ~n338 & n360;
  assign n362 = n336 & n361;
  assign n363 = n330 & n362;
  assign n364 = n326 & n363;
  assign n365 = n315 & n364;
  assign n366 = n301 & n365;
  assign b2 = ~n281 | ~n366;
  assign n368 = v & n93;
  assign n369 = u & n368;
  assign n370 = n128 & n302;
  assign n371 = n128 & n369;
  assign n372 = y & n162;
  assign n373 = ~n347 & ~n370;
  assign n374 = ~n372 & n373;
  assign y0 = n371 | ~n374;
  assign n376 = n199 & ~y0;
  assign n377 = n227 & n376;
  assign n378 = ~n202 & ~n228;
  assign n379 = n96 & n106;
  assign n380 = x & n263;
  assign n381 = ~n379 & ~n380;
  assign n382 = b & ~u;
  assign n383 = n212 & n382;
  assign n384 = n109 & n383;
  assign n385 = n213 & n382;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n249 & n386;
  assign n388 = n107 & n157;
  assign n389 = n107 & n189;
  assign n390 = n303 & n389;
  assign n391 = z & n106;
  assign n392 = n159 & n391;
  assign n393 = ~a0 & n388;
  assign n394 = y & n388;
  assign n395 = n106 & n203;
  assign n396 = n106 & n369;
  assign n397 = n106 & n302;
  assign n398 = ~n345 & ~n397;
  assign n399 = ~n396 & n398;
  assign n400 = ~n395 & n399;
  assign n401 = ~n394 & n400;
  assign n402 = ~n393 & n401;
  assign n403 = ~n392 & n402;
  assign n404 = ~n390 & n403;
  assign n405 = a0 & n388;
  assign n406 = n172 & n183;
  assign n407 = n159 & n183;
  assign n408 = ~n405 & ~n407;
  assign q1 = n406 | ~n408;
  assign n410 = n404 & ~q1;
  assign n411 = n387 & n410;
  assign n412 = n0 & q0;
  assign n413 = n260 & n412;
  assign n414 = n255 & n263;
  assign n415 = ~n413 & ~n414;
  assign n416 = t & n117;
  assign n417 = n113 & n129;
  assign n418 = a0 & n113;
  assign n419 = n200 & n418;
  assign n420 = n160 & n417;
  assign n421 = w & n417;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~n419 & n422;
  assign n424 = n110 & n114;
  assign n425 = n96 & n113;
  assign n426 = n114 & n190;
  assign n427 = n109 & n424;
  assign n428 = n114 & n207;
  assign n429 = ~n425 & ~n428;
  assign n430 = ~n427 & n429;
  assign t1 = n426 | ~n430;
  assign n432 = x & n114;
  assign n433 = n416 & n432;
  assign n434 = n423 & ~t1;
  assign n435 = ~n433 & n434;
  assign n436 = n113 & n331;
  assign n437 = n182 & n436;
  assign n438 = n316 & n417;
  assign n439 = ~n437 & ~n438;
  assign n440 = w & n114;
  assign n441 = n416 & n440;
  assign n442 = n439 & ~n441;
  assign n443 = n134 & n283;
  assign n444 = n172 & n391;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~g & n205;
  assign n447 = ~g & n126;
  assign n448 = n327 & n447;
  assign n449 = n119 & n204;
  assign n450 = y & n424;
  assign n451 = ~d & n102;
  assign n452 = n101 & n451;
  assign n453 = n122 & ~n452;
  assign n454 = ~n450 & n453;
  assign n455 = ~n340 & n454;
  assign n456 = ~n449 & n455;
  assign n457 = ~n448 & n456;
  assign n458 = ~n446 & n457;
  assign n459 = n445 & n458;
  assign n460 = n330 & n459;
  assign n461 = n442 & n460;
  assign n462 = n435 & n461;
  assign n463 = n415 & n462;
  assign n464 = n411 & n463;
  assign n465 = n381 & n464;
  assign n466 = n195 & n465;
  assign n467 = n181 & n466;
  assign n468 = n248 & n467;
  assign n469 = n378 & n468;
  assign c2 = ~n377 | ~n469;
  assign n471 = n301 & n415;
  assign o1 = n127 & n183;
  assign n1 = n200 & n304;
  assign n474 = z & n317;
  assign n475 = w & n317;
  assign n476 = ~o1 & ~n1;
  assign n477 = n130 & n183;
  assign n478 = n476 & ~n477;
  assign n479 = ~n475 & n478;
  assign n480 = ~n474 & n479;
  assign n481 = n445 & n480;
  assign n482 = n107 & n416;
  assign n483 = b & x;
  assign n484 = n482 & n483;
  assign n485 = b & w;
  assign n486 = n482 & n485;
  assign n487 = ~n484 & ~n486;
  assign n488 = n481 & n487;
  assign n489 = n107 & n126;
  assign n490 = n107 & n119;
  assign n491 = ~n489 & ~n490;
  assign n492 = n326 & n491;
  assign n493 = n157 & n283;
  assign n494 = n97 & n158;
  assign n495 = n131 & n494;
  assign n496 = a0 & n493;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n305 & ~n343;
  assign n499 = ~n250 & n498;
  assign n500 = n497 & n499;
  assign n501 = n492 & n500;
  assign n502 = n488 & n501;
  assign n503 = n411 & n502;
  assign d1 = ~n471 | ~n503;
  assign n505 = n157 & n269;
  assign n506 = h & ~q;
  assign n507 = i & q;
  assign n508 = ~n506 & ~n507;
  assign n509 = n & ~v;
  assign n510 = n241 & n509;
  assign n511 = ~w0 & ~n510;
  assign n512 = n336 & ~n452;
  assign n513 = ~n343 & n512;
  assign n514 = n113 & n158;
  assign n515 = ~f & p;
  assign n516 = n514 & n515;
  assign n517 = n132 & n254;
  assign n518 = n303 & n517;
  assign n519 = ~h & ~q;
  assign n520 = n518 & n519;
  assign n521 = ~i & q;
  assign n522 = n518 & n521;
  assign n523 = n214 & n515;
  assign n524 = ~o & ~b0;
  assign n525 = n155 & n524;
  assign n526 = n102 & n525;
  assign n527 = n118 & n526;
  assign n528 = ~x & n110;
  assign n529 = n254 & n528;
  assign n530 = n240 & n529;
  assign n531 = ~n170 & ~n171;
  assign n532 = n141 & n531;
  assign x1 = ~n378 | ~n532;
  assign n534 = n505 & n508;
  assign n535 = ~z1 & ~x1;
  assign n536 = ~n210 & n535;
  assign n537 = ~n112 & n536;
  assign n538 = ~n105 & n537;
  assign n539 = ~n444 & n538;
  assign n540 = ~n413 & n539;
  assign n541 = ~n310 & n540;
  assign n542 = ~n379 & n541;
  assign n543 = ~n530 & n542;
  assign n544 = ~n527 & n543;
  assign n545 = ~n523 & n544;
  assign n546 = ~n522 & n545;
  assign n547 = ~n520 & n546;
  assign n548 = ~n516 & n547;
  assign n549 = n410 & n548;
  assign n550 = n513 & n549;
  assign n551 = n511 & n550;
  assign n552 = n195 & n551;
  assign n553 = n281 & n552;
  assign d2 = n534 | ~n553;
  assign n555 = c0 & n211;
  assign n556 = n283 & n555;
  assign n557 = n497 & ~n556;
  assign n558 = ~u & n109;
  assign n559 = n344 & n558;
  assign n560 = ~u & n189;
  assign n561 = n344 & n560;
  assign n562 = n172 & n309;
  assign n563 = ~n493 & n557;
  assign n564 = ~n562 & n563;
  assign n565 = ~n561 & n564;
  assign n566 = ~n559 & n565;
  assign n567 = n315 & n566;
  assign n568 = n513 & n567;
  assign n569 = ~n342 & n492;
  assign n570 = n411 & n569;
  assign e1 = ~n568 | ~n570;
  assign n572 = e0 & n368;
  assign n573 = ~k & z;
  assign n574 = f & n514;
  assign n575 = s & e0;
  assign n576 = n118 & n575;
  assign n577 = ~u & n572;
  assign n578 = n160 & n576;
  assign n579 = n158 & n573;
  assign n580 = n154 & n579;
  assign n581 = ~s & n157;
  assign n582 = n573 & n581;
  assign n583 = n573 & n574;
  assign n584 = n573 & n576;
  assign n585 = n273 & n573;
  assign n586 = n573 & n577;
  assign n587 = ~n578 & ~n586;
  assign n588 = ~n585 & n587;
  assign n589 = ~n584 & n588;
  assign n590 = ~n583 & n589;
  assign n591 = ~n582 & n590;
  assign n592 = ~n580 & n591;
  assign n593 = x & n257;
  assign n594 = ~g0 & n593;
  assign n595 = n282 & n594;
  assign n596 = ~i0 & n595;
  assign n597 = ~j0 & n596;
  assign n598 = n113 & n256;
  assign n599 = n269 & n598;
  assign n600 = k0 & n597;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~k0 & l0;
  assign n603 = n597 & n602;
  assign n604 = i0 & n595;
  assign n605 = ~n603 & ~n604;
  assign n606 = n601 & n605;
  assign n607 = j0 & n596;
  assign n608 = ~f0 & g0;
  assign n609 = n593 & n608;
  assign n610 = ~n607 & ~n609;
  assign n611 = f0 & n593;
  assign n612 = n610 & ~n611;
  assign n613 = y & n107;
  assign n614 = n110 & n613;
  assign n615 = ~f0 & h0;
  assign n616 = n594 & n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = n612 & n617;
  assign n619 = n606 & n618;
  assign n620 = n592 & n619;
  assign n621 = ~r0 & ~s0;
  assign n622 = n293 & n621;
  assign n623 = w & n577;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~s & e0;
  assign n626 = n256 & n625;
  assign n627 = n132 & n626;
  assign n628 = ~n342 & ~n627;
  assign n629 = n624 & n628;
  assign n630 = n381 & n629;
  assign n631 = n160 & n574;
  assign n632 = ~z & n574;
  assign n633 = f & n214;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n631 & n634;
  assign n636 = u & w;
  assign n637 = n572 & n636;
  assign n638 = a0 & n424;
  assign n639 = w & n576;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n637 & n640;
  assign n642 = x & n110;
  assign n643 = n575 & n642;
  assign n644 = n442 & ~n643;
  assign n645 = n435 & n644;
  assign n646 = n114 & n133;
  assign n647 = n109 & n646;
  assign n648 = w & n110;
  assign n649 = n575 & n648;
  assign n650 = ~n647 & ~n649;
  assign n651 = n316 & n646;
  assign n652 = n650 & ~n651;
  assign n653 = n645 & n652;
  assign l2 = w & n424;
  assign k2 = n450 | l2;
  assign n656 = n417 & n573;
  assign n657 = n653 & ~k2;
  assign n658 = ~n656 & n657;
  assign n659 = f & n107;
  assign n660 = n208 & n659;
  assign n661 = d & n107;
  assign n662 = n207 & n661;
  assign n663 = ~n660 & ~n662;
  assign n664 = ~n250 & n330;
  assign n665 = ~c0 & n106;
  assign n666 = n101 & n665;
  assign n667 = o & n102;
  assign n668 = n92 & n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = n97 & n369;
  assign n671 = n160 & n577;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~k0 & ~l0;
  assign n674 = n597 & n673;
  assign n675 = n506 & n518;
  assign n676 = n507 & n518;
  assign n677 = g & n205;
  assign n678 = g & n126;
  assign n679 = n327 & n678;
  assign n680 = n116 & n134;
  assign n681 = n190 & n659;
  assign n682 = ~n325 & ~n444;
  assign n683 = ~n681 & n682;
  assign n684 = ~n680 & n683;
  assign n685 = ~n246 & n684;
  assign n686 = n487 & n685;
  assign n687 = n480 & n686;
  assign n688 = n491 & n687;
  assign g2 = ~n411 | ~n688;
  assign n690 = a0 & n572;
  assign n691 = ~z1 & ~g2;
  assign n692 = ~n192 & n691;
  assign n693 = ~n188 & n692;
  assign n694 = ~n443 & n693;
  assign n695 = ~n679 & n694;
  assign n696 = ~n677 & n695;
  assign n697 = ~n247 & n696;
  assign n698 = ~n676 & n697;
  assign n699 = ~n675 & n698;
  assign n700 = ~n674 & n699;
  assign n701 = ~n340 & n700;
  assign n702 = ~n339 & n701;
  assign n703 = ~n338 & n702;
  assign n704 = ~n449 & n703;
  assign n705 = ~n448 & n704;
  assign n706 = ~n446 & n705;
  assign n707 = ~n530 & n706;
  assign n708 = ~n527 & n707;
  assign n709 = ~n523 & n708;
  assign n710 = ~n522 & n709;
  assign n711 = ~n520 & n710;
  assign n712 = ~n516 & n711;
  assign n713 = n323 & n712;
  assign n714 = n672 & n713;
  assign n715 = n669 & n714;
  assign n716 = n511 & n715;
  assign n717 = n664 & n716;
  assign n718 = n568 & n717;
  assign n719 = n471 & n718;
  assign n720 = n181 & n719;
  assign n721 = n124 & n720;
  assign n722 = n663 & n721;
  assign n723 = n378 & n722;
  assign n724 = n658 & n723;
  assign n725 = n641 & n724;
  assign n726 = n635 & n725;
  assign n727 = n377 & n726;
  assign n728 = n630 & n727;
  assign n729 = n620 & n728;
  assign n730 = n281 & n729;
  assign n731 = ~n505 & n730;
  assign e2 = n690 | ~n731;
  assign n733 = n410 & n488;
  assign n734 = a0 & n577;
  assign n735 = n672 & ~n734;
  assign n736 = ~n249 & ~n250;
  assign n737 = ~n414 & n736;
  assign n738 = ~n295 & n737;
  assign n739 = ~n622 & n738;
  assign n740 = n492 & n739;
  assign n741 = n735 & n740;
  assign n742 = n568 & n741;
  assign f1 = ~n733 | ~n742;
  assign n744 = ~a & n113;
  assign n745 = n302 & n744;
  assign n746 = y & n369;
  assign n747 = n744 & n746;
  assign n748 = ~a & y;
  assign n749 = n161 & n748;
  assign u0 = n747 | n749;
  assign n751 = ~a & u;
  assign n752 = v & n751;
  assign n753 = w & n752;
  assign n754 = n114 & n753;
  assign n755 = n153 & n754;
  assign n756 = ~a & ~f;
  assign n757 = w & n756;
  assign n758 = n107 & n757;
  assign n759 = n133 & n758;
  assign n760 = n107 & n756;
  assign n761 = n208 & n760;
  assign n762 = n155 & n156;
  assign n763 = n153 & n762;
  assign n764 = n744 & n763;
  assign n765 = ~a & a0;
  assign n766 = c0 & n765;
  assign n767 = n417 & n766;
  assign n768 = ~a & d;
  assign n769 = ~d0 & n768;
  assign n770 = n101 & n769;
  assign n771 = ~b & ~u;
  assign n772 = n212 & n771;
  assign n773 = n109 & n772;
  assign n774 = ~a & n107;
  assign n775 = n110 & n774;
  assign n776 = n109 & n775;
  assign n777 = ~a & ~c0;
  assign n778 = n129 & n777;
  assign n779 = n183 & n778;
  assign n780 = ~b & x;
  assign n781 = n482 & n780;
  assign n782 = ~b & w;
  assign n783 = n482 & n782;
  assign n784 = n98 & n756;
  assign n785 = ~a & n126;
  assign n786 = n116 & n785;
  assign n787 = n127 & n131;
  assign n788 = n744 & n787;
  assign n789 = ~a & z;
  assign n790 = n168 & n789;
  assign n791 = ~a & w;
  assign n792 = n168 & n791;
  assign n793 = n213 & n771;
  assign n794 = ~a & n183;
  assign n795 = n182 & n794;
  assign n796 = n134 & n774;
  assign n797 = n161 & n765;
  assign n798 = n161 & n789;
  assign n799 = n161 & n791;
  assign n800 = ~a & c0;
  assign n801 = n212 & n800;
  assign n802 = ~a & n449;
  assign n803 = ~n745 & ~u0;
  assign n804 = ~n139 & n803;
  assign n805 = ~n802 & n804;
  assign n806 = ~n801 & n805;
  assign n807 = ~n799 & n806;
  assign n808 = ~n798 & n807;
  assign n809 = ~n797 & n808;
  assign n810 = ~n796 & n809;
  assign n811 = ~n795 & n810;
  assign n812 = ~n793 & n811;
  assign n813 = ~n792 & n812;
  assign n814 = ~n790 & n813;
  assign n815 = ~n788 & n814;
  assign n816 = ~n786 & n815;
  assign n817 = ~n784 & n816;
  assign n818 = ~n783 & n817;
  assign n819 = ~n781 & n818;
  assign n820 = ~n779 & n819;
  assign n821 = ~n776 & n820;
  assign n822 = ~n773 & n821;
  assign n823 = ~n770 & n822;
  assign n824 = ~n767 & n823;
  assign n825 = ~n764 & n824;
  assign n826 = ~n761 & n825;
  assign n827 = ~n759 & n826;
  assign f2 = n755 | ~n827;
  assign n829 = n488 & n664;
  assign n830 = n & v;
  assign n831 = n241 & n830;
  assign n832 = ~n413 & ~n668;
  assign n833 = ~n831 & n832;
  assign n834 = n386 & n833;
  assign n835 = n512 & n834;
  assign n836 = n290 & n835;
  assign n837 = n298 & n836;
  assign n838 = n735 & n837;
  assign n839 = n653 & n838;
  assign g1 = ~n829 | ~n839;
  assign n841 = ~n384 & ~n734;
  assign n842 = n512 & n841;
  assign n843 = n308 & n842;
  assign n844 = n557 & n843;
  assign n845 = n268 & n844;
  assign n846 = n292 & n845;
  assign h1 = ~n829 | ~n846;
  assign n848 = ~n247 & ~n681;
  assign n849 = n663 & n848;
  assign h2 = ~n635 | ~n849;
  assign n851 = n669 & ~n831;
  assign n852 = ~n450 & n851;
  assign n853 = ~n370 & n492;
  assign n854 = ~n121 & ~n206;
  assign n855 = ~n105 & n854;
  assign n856 = ~n679 & n855;
  assign n857 = ~n677 & n856;
  assign n858 = ~n681 & n857;
  assign n859 = ~n680 & n858;
  assign n860 = n663 & n859;
  assign u1 = ~n248 | ~n860;
  assign n862 = ~a2 & ~u1;
  assign n863 = ~n343 & n862;
  assign n864 = ~n271 & n863;
  assign n865 = ~n380 & n864;
  assign n866 = n386 & n865;
  assign n867 = n442 & n866;
  assign n868 = n628 & n867;
  assign n869 = n605 & n868;
  assign n870 = n612 & n869;
  assign n871 = n853 & n870;
  assign n872 = n733 & n871;
  assign i1 = ~n852 | ~n872;
  assign n874 = ~q1 & ~u1;
  assign n875 = ~n425 & n874;
  assign n876 = ~l2 & n875;
  assign n877 = ~n614 & n876;
  assign n878 = ~n379 & n877;
  assign n879 = n439 & n878;
  assign n880 = n423 & n879;
  assign n881 = n513 & n880;
  assign n882 = n652 & n881;
  assign n883 = n851 & n882;
  assign n884 = n471 & n883;
  assign j1 = ~n829 | ~n884;
  assign n886 = ~n405 & ~n603;
  assign n887 = n336 & n886;
  assign n888 = n404 & n887;
  assign n889 = n481 & n888;
  assign n890 = n650 & n889;
  assign n891 = n387 & n890;
  assign n892 = n492 & n891;
  assign n893 = n268 & n892;
  assign n894 = n644 & n893;
  assign n895 = n601 & n894;
  assign n896 = n664 & n895;
  assign n897 = n735 & n896;
  assign n898 = n567 & n897;
  assign n899 = n852 & n898;
  assign k1 = ~n630 | ~n899;
  assign n901 = ~n441 & ~n452;
  assign n902 = ~n607 & n901;
  assign n903 = ~n578 & n902;
  assign n904 = n404 & n903;
  assign n905 = n487 & n904;
  assign n906 = n387 & n905;
  assign n907 = n435 & n906;
  assign n908 = n652 & n907;
  assign n909 = n606 & n908;
  assign n910 = n853 & n909;
  assign l1 = ~n852 | ~n910;
  assign n912 = ~n484 & ~n647;
  assign n913 = ~n666 & n912;
  assign n914 = ~l2 & n913;
  assign n915 = n330 & n914;
  assign n916 = n513 & n915;
  assign n917 = n628 & n916;
  assign n918 = n610 & n917;
  assign n919 = n411 & n918;
  assign n920 = n645 & n919;
  assign n921 = n617 & n920;
  assign m1 = ~n853 | ~n921;
  assign n923 = ~n370 & n862;
  assign n924 = n386 & n923;
  assign n925 = n330 & n924;
  assign n926 = n326 & n925;
  assign n927 = n669 & n926;
  assign n928 = n735 & n927;
  assign n929 = n272 & n928;
  assign n930 = n568 & n929;
  assign n931 = n471 & n930;
  assign n932 = n733 & n931;
  assign n933 = n658 & n932;
  assign n934 = n630 & n933;
  assign p1 = ~n620 | ~n934;
  assign n936 = ~n380 & ~n831;
  assign n937 = n592 & n936;
  assign n938 = n658 & n937;
  assign s1 = ~n641 | ~n938;
  assign n940 = ~n274 & ~n348;
  assign x0 = n747 | ~n940;
  assign n942 = ~n749 & ~x0;
  assign n943 = ~n349 & n942;
  assign t0 = n745 | ~n943;
  assign n945 = n505 & ~n508;
  assign n946 = ~n627 & ~l2;
  assign n947 = ~n676 & n946;
  assign n948 = ~n675 & n947;
  assign n949 = ~n674 & n948;
  assign n950 = n566 & n949;
  assign n951 = n735 & n950;
  assign n952 = n624 & n951;
  assign n953 = n641 & n952;
  assign n954 = n635 & n953;
  assign n955 = n620 & n954;
  assign v1 = n945 | ~n955;
  assign n957 = n177 & n195;
  assign n958 = n124 & n957;
  assign n959 = n167 & n958;
  assign w1 = ~n377 | ~n959;
  assign j2 = 1'b0;
  assign v0 = 1'b0;
  assign r1 = l2;
endmodule


