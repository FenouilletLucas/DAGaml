// Benchmark "top" written by ABC on Sun Apr 24 20:32:55 2016

module top ( clock, 
    tin_pv10_4_4_, tin_pv11_4_4_, tin_pv6_7_7_, tin_pv2_0_0_,
    tin_pv10_3_3_, tin_pv1_2_2_, tin_pv11_3_3_, tin_pv4_3_3_,
    tin_pv10_2_2_, tin_pv11_2_2_, tin_pv6_0_0_, tin_pv2_1_1_,
    tin_pv10_1_1_, tin_pv1_3_3_, preset_0_0_, tin_pv11_1_1_, tin_pv4_4_4_,
    tin_pready_0_0_, tin_pv10_0_0_, tin_pv11_0_0_, tin_pv6_1_1_,
    tin_pv2_2_2_, tin_pv1_4_4_, tin_pv4_5_5_, tin_pv6_2_2_, tin_pv2_3_3_,
    tin_pv1_5_5_, tin_pv4_6_6_, tin_pv6_3_3_, tin_pv2_4_4_, tin_pv1_6_6_,
    pclk, tin_pv4_7_7_, tin_pv6_4_4_, tin_pv2_5_5_, tin_pv1_7_7_,
    tin_pv4_0_0_, tin_pv6_5_5_, tin_pv2_6_6_, tin_pv10_7_7_, tin_pv1_0_0_,
    tin_pv11_7_7_, tin_pv4_1_1_, tin_pv10_6_6_, tin_pv11_6_6_,
    tin_pv6_6_6_, tin_pv2_7_7_, preset, tin_pv10_5_5_, tin_pv1_1_1_,
    tin_pv11_5_5_, tin_pv4_2_2_,
    pv14_2_2_, pv12_3_3_, pv10_4_4_, pv7_5_5_, pv3_6_6_, pv15_2_2_,
    pv13_3_3_, pv11_4_4_, pv6_7_7_, pv2_0_0_, pv14_1_1_, pv12_2_2_,
    pv10_3_3_, pv9_0_0_, pv5_1_1_, pv1_2_2_, pv15_1_1_, pv13_2_2_,
    pv11_3_3_, pv8_2_2_, pv4_3_3_, pv14_0_0_, pv12_1_1_, pv10_2_2_,
    pv7_6_6_, pv3_7_7_, pv15_0_0_, pv13_1_1_, pv11_2_2_, pv6_0_0_,
    pv2_1_1_, pv12_0_0_, pv10_1_1_, pv9_1_1_, pv5_2_2_, pv1_3_3_,
    pv13_0_0_, pv11_1_1_, pv8_3_3_, pv4_4_4_, pready_0_0_, pv10_0_0_,
    pv7_7_7_, pv3_0_0_, pv11_0_0_, pv6_1_1_, pv2_2_2_, pv9_2_2_, pv5_3_3_,
    pv1_4_4_, pv8_4_4_, pv4_5_5_, pv7_0_0_, pv3_1_1_, pv6_2_2_, pv2_3_3_,
    pv9_3_3_, pv5_4_4_, pv1_5_5_, pv8_5_5_, pv4_6_6_, pv7_1_1_, pv3_2_2_,
    pv6_3_3_, pv2_4_4_, pv9_4_4_, pv5_5_5_, pv1_6_6_, pv8_6_6_, pv4_7_7_,
    pv7_2_2_, pv3_3_3_, pv6_4_4_, pv2_5_5_, pv14_7_7_, pv9_5_5_, pv5_6_6_,
    pv1_7_7_, pv15_7_7_, pv8_7_7_, pv4_0_0_, pv14_6_6_, pv12_7_7_,
    pv7_3_3_, pv3_4_4_, pv15_6_6_, pv13_7_7_, pv6_5_5_, pv2_6_6_, pdn,
    pv14_5_5_, pv12_6_6_, pv10_7_7_, pv9_6_6_, pv5_7_7_, pv1_0_0_,
    pv15_5_5_, pv13_6_6_, pv11_7_7_, pv8_0_0_, pv4_1_1_, pv14_4_4_,
    pv12_5_5_, pv10_6_6_, pv7_4_4_, pv3_5_5_, pv15_4_4_, pv13_5_5_,
    pv11_6_6_, pv6_6_6_, pv2_7_7_, pv14_3_3_, pv12_4_4_, pv10_5_5_,
    pv9_7_7_, pv5_0_0_, pv1_1_1_, pv15_3_3_, pv13_4_4_, pv11_5_5_,
    pv8_1_1_, pv4_2_2_  );
  input  clock;
  input  tin_pv10_4_4_, tin_pv11_4_4_, tin_pv6_7_7_, tin_pv2_0_0_,
    tin_pv10_3_3_, tin_pv1_2_2_, tin_pv11_3_3_, tin_pv4_3_3_,
    tin_pv10_2_2_, tin_pv11_2_2_, tin_pv6_0_0_, tin_pv2_1_1_,
    tin_pv10_1_1_, tin_pv1_3_3_, preset_0_0_, tin_pv11_1_1_, tin_pv4_4_4_,
    tin_pready_0_0_, tin_pv10_0_0_, tin_pv11_0_0_, tin_pv6_1_1_,
    tin_pv2_2_2_, tin_pv1_4_4_, tin_pv4_5_5_, tin_pv6_2_2_, tin_pv2_3_3_,
    tin_pv1_5_5_, tin_pv4_6_6_, tin_pv6_3_3_, tin_pv2_4_4_, tin_pv1_6_6_,
    pclk, tin_pv4_7_7_, tin_pv6_4_4_, tin_pv2_5_5_, tin_pv1_7_7_,
    tin_pv4_0_0_, tin_pv6_5_5_, tin_pv2_6_6_, tin_pv10_7_7_, tin_pv1_0_0_,
    tin_pv11_7_7_, tin_pv4_1_1_, tin_pv10_6_6_, tin_pv11_6_6_,
    tin_pv6_6_6_, tin_pv2_7_7_, preset, tin_pv10_5_5_, tin_pv1_1_1_,
    tin_pv11_5_5_, tin_pv4_2_2_;
  output pv14_2_2_, pv12_3_3_, pv10_4_4_, pv7_5_5_, pv3_6_6_, pv15_2_2_,
    pv13_3_3_, pv11_4_4_, pv6_7_7_, pv2_0_0_, pv14_1_1_, pv12_2_2_,
    pv10_3_3_, pv9_0_0_, pv5_1_1_, pv1_2_2_, pv15_1_1_, pv13_2_2_,
    pv11_3_3_, pv8_2_2_, pv4_3_3_, pv14_0_0_, pv12_1_1_, pv10_2_2_,
    pv7_6_6_, pv3_7_7_, pv15_0_0_, pv13_1_1_, pv11_2_2_, pv6_0_0_,
    pv2_1_1_, pv12_0_0_, pv10_1_1_, pv9_1_1_, pv5_2_2_, pv1_3_3_,
    pv13_0_0_, pv11_1_1_, pv8_3_3_, pv4_4_4_, pready_0_0_, pv10_0_0_,
    pv7_7_7_, pv3_0_0_, pv11_0_0_, pv6_1_1_, pv2_2_2_, pv9_2_2_, pv5_3_3_,
    pv1_4_4_, pv8_4_4_, pv4_5_5_, pv7_0_0_, pv3_1_1_, pv6_2_2_, pv2_3_3_,
    pv9_3_3_, pv5_4_4_, pv1_5_5_, pv8_5_5_, pv4_6_6_, pv7_1_1_, pv3_2_2_,
    pv6_3_3_, pv2_4_4_, pv9_4_4_, pv5_5_5_, pv1_6_6_, pv8_6_6_, pv4_7_7_,
    pv7_2_2_, pv3_3_3_, pv6_4_4_, pv2_5_5_, pv14_7_7_, pv9_5_5_, pv5_6_6_,
    pv1_7_7_, pv15_7_7_, pv8_7_7_, pv4_0_0_, pv14_6_6_, pv12_7_7_,
    pv7_3_3_, pv3_4_4_, pv15_6_6_, pv13_7_7_, pv6_5_5_, pv2_6_6_, pdn,
    pv14_5_5_, pv12_6_6_, pv10_7_7_, pv9_6_6_, pv5_7_7_, pv1_0_0_,
    pv15_5_5_, pv13_6_6_, pv11_7_7_, pv8_0_0_, pv4_1_1_, pv14_4_4_,
    pv12_5_5_, pv10_6_6_, pv7_4_4_, pv3_5_5_, pv15_4_4_, pv13_5_5_,
    pv11_6_6_, pv6_6_6_, pv2_7_7_, pv14_3_3_, pv12_4_4_, pv10_5_5_,
    pv9_7_7_, pv5_0_0_, pv1_1_1_, pv15_3_3_, pv13_4_4_, pv11_5_5_,
    pv8_1_1_, pv4_2_2_;
  reg n_n4142, n_n3936, n_n3574, n_n3008, n_n3726, n_n3604, n_n3144,
    n_n3782, n_n3067, n_n4258, n_n3225, n_n3180, n_n3274, n_n3475, n_n3687,
    n_n3381, n_n3098, n_n4108, n_n3497, n_n3793, n_n4316, n_n4349, n_n3029,
    n_n3619, n_n3264, n_n3780, ndn3_4, n_n4114, n_n3146, n_n3511, n_n3152,
    n_n3833, n_n4282, n_n3305, n_n4392, n_n4224, n_n3198, n_n3204, n_n3024,
    n_n4139, ndn3_15, n_n3133, n_n4074, n_n3270, n_n3858, n_n3456, n_n3521,
    n_n3081, n_n4381, n_n3670, n_n4211, n_n3493, n_n3495, n_n3916, n_n3195,
    n_n3525, n_n3729, n_n3876, ndn3_5, n_n3549, n_n3489, n_n3764, n_n3281,
    n_n3707, n_n3517, n_n4160, n_n4222, n_n3012, n_n4071, n_n3372, n_n3344,
    n_n3688, n_n3079, n_n3313, n_n3411, n_n3231, n_n3396, n_n3432, n_n3606,
    n_n3733, n_n3556, n_n4040, n_n3120, n_n3221, n_n3173, n_n3851, n_n3113,
    n_n3242, n_n3118, n_n3376, n_n4089, n_n3044, n_n3627, n_n3035, n_n3111,
    n_n3321, n_n3443, n_n3215, ndn3_10, n_n4172, nlc1_2, n_n3590, n_n4110,
    nlc3_3, n_n3576, n_n4129, n_n4189, n_n4286, n_n4383, pdn, n_n3567,
    n_n3892, n_n3075, n_n3354, n_n3465, ndn3_6, n_n3617, n_n4162, n_n3207,
    n_n4120, n_n3065, n_n4005, n_n3266, n_n4337, n_n3600, n_n3415, n_n4243,
    n_n3872, n_n3648, n_n3358, n_n3350, ndn3_7, n_n3116, n_n3583, n_n3906,
    n_n4131, n_n3316, n_n3061, n_n3048, n_n3886, n_n3919, n_n3128, n_n3995,
    n_n4213, n_n3761, ndn3_8, n_n3252, n_n4366, n_n3328, n_n3988, n_n3348,
    n_n3544, n_n3101, n_n4279, n_n3896, n_n3736, n_n4251, n_n3650, n_n3307,
    n_n4294, n_n4334, n_n3955, n_n4164, n_n3155, n_n3749, n_n4233, n_n4347,
    n_n3826, n_n3360, n_n3458, n_n3093, n_n3157, n_n3506, n_n3161, n_n3319,
    n_n3429, n_n3971, n_n3449, n_n4270, n_n4288, n_n3183, n_n3130, nlak4_2,
    n_n4047, n_n3978, n_n3239, n_n4145, n_n3890, n_n4003, n_n3091, n_n3985,
    n_n3326, n_n4052, nsr4_2, n_n4099, n_n4375, n_n4067, n_n4290, n_n3898,
    n_n4122, n_n3774, n_n3014, n_n4241, n_n3952, n_n3237, n_n3968, n_n3922,
    n_n3551, n_n3379, n_n4275, n_n3570, n_n3854, n_n4057, n_n3451, n_n4037,
    n_n3408, n_n4229, n_n4201, n_n3339, n_n4362, n_n3483, n_n3557, n_n4185,
    n_n3069, n_n3643, n_n3404, n_n3057, n_n3020, n_n3828, n_n3631, n_n3138,
    nsr1_2, n_n4065, n_n3679, n_n3287, n_n4351, n_n4059, n_n3436, nen3_10,
    n_n3461, n_n4012, n_n3051, n_n3073, n_n3777, n_n3709, n_n3946, n_n3085,
    n_n3259, n_n3504, n_n4045, n_n3954, n_n3136, n_n4372, n_n4236, n_n3040,
    n_n3874, n_n3999, n_n3223, ndn1_34, n_n3743, n_n3657, n_n3213, n_n3095,
    n_n3663, n_n3724, n_n3038, n_n3370, n_n3624, n_n3578, n_n3713, n_n3089,
    n_n3211, n_n3367, n_n3434, n_n3126, n_n4192, n_n4136, n_n3053, n_n3938,
    n_n3769, n_n4390, nsr3_17, n_n3903, n_n3658, nrq3_11, n_n3818, n_n3533,
    n_n3463, n_n3175, n_n3055, n_n3202, n_n3385, n_n4077, n_n3142, n_n3901,
    n_n3934, n_n3823, n_n3722, n_n4309, n_n4159, n_n4330, n_n3836, n_n3470,
    n_n3331, n_n3883, n_n4299, n_n4157, ndn3_9, n_n3208, n_n3190, n_n4029,
    n_n3042, nsr3_14, n_n4151, n_n3188, n_n4303, n_n3250, n_n3170, n_n3758,
    n_n3910, n_n3108, n_n3150, n_n4320, n_n4360, n_n4247, n_n4199, n_n3966,
    n_n3766, n_n4021, n_n4062, n_n3514, n_n3572, n_n4166, n_n3976, n_n3394,
    n_n4095, n_n3863, n_n3720, ngfdn_3, n_n3756, n_n3667, n_n3342, n_n3529,
    n_n4209, n_n4324, n_n3337, n_n4227, n_n4153, n_n3831, n_n3233, n_n4263,
    n_n3413, n_n4182, n_n3841, n_n3441, n_n4026, n_n4342, n_n4102, n_n3277,
    n_n4180, n_n3878, n_n3931, n_n3845, n_n3865, n_n3486, n_n4056, n_n3674,
    n_n3959, n_n3608, n_n4080, n_n4018, n_n4354, n_n3797, n_n3739, n_n3646,
    n_n3099, n_n3537, n_n3806, n_n3087, n_n4105, n_n3262, n_n4125, n_n3814,
    n_n4093, nsr3_3;
  wire n1333, n1334_1, n1340, n1341, n1343, n1344_1, n1346, n1347, n1351,
    n1352, n1356, n1357, n1361, n1362, n1365, n1366, n1370, n1371, n1377,
    n1378, n1380, n1381, n1383, n1384_1, n1387, n1388, n1392, n1393, n1396,
    n1397, n1400, n1401, n1403, n1404_1, n1406, n1407, n1411, n1412,
    n1414_1, n1415, n1417, n1418, n1422, n1423, n1426, n1427, n1431, n1432,
    n1434_1, n1435, n1439_1, n1440, n1443, n1444_1, n1448, n1449_1, n1451,
    n1452, n1456, n1457, n1460, n1461, n1465, n1466, n1468, n1469_1,
    n1474_1, n1475, n1479_1, n1480, n1488, n1489_1, n1491, n1492, n1496,
    n1497, n1501, n1502, n1506, n1507, n1510, n1511, n1515, n1516, n1522,
    n1523, n1525, n1526, n1528, n1529_1, n1533, n1534_1, n1538, n1539_1,
    n1543, n1544_1, n1547, n1548, n1550, n1551, n1552, n1553, n1554_1,
    n1555, n1556, n1557, n1558, n1559_1, n1560, n1561, n1562, n1563,
    n1564_1, n1565, n1566, n1567, n1568, n1569_1, n1570, n1571, n1572,
    n1573, n1574_1, n1575, n1576, n1577, n1578, n1579_1, n1580, n1581,
    n1582, n1583, n1584_1, n1585, n1586, n1587, n1588, n1589_1, n1590,
    n1591, n1592, n1593, n1594_1, n1595, n1596, n1597, n1598, n1599_1,
    n1600, n1601, n1602, n1603, n1604_1, n1605, n1606, n1607, n1608,
    n1609_1, n1610, n1611, n1612, n1613, n1614_1, n1615, n1616, n1617,
    n1618, n1619_1, n1620, n1621, n1622, n1623, n1624_1, n1625, n1626,
    n1627, n1628, n1629_1, n1630, n1631, n1632, n1633, n1634_1, n1635,
    n1636, n1637, n1638, n1639_1, n1640, n1641, n1642, n1643, n1644_1,
    n1645, n1646, n1647, n1648, n1649_1, n1650, n1651, n1652, n1653,
    n1654_1, n1655, n1656, n1657, n1658, n1659_1, n1660, n1661, n1662,
    n1663, n1664_1, n1665, n1666, n1667, n1668, n1669_1, n1670, n1671,
    n1672, n1673, n1674_1, n1676, n1677, n1678, n1679_1, n1681, n1682,
    n1683, n1684_1, n1685, n1686, n1687, n1688, n1689_1, n1690, n1691,
    n1692, n1693, n1694_1, n1695, n1696, n1697, n1698, n1699_1, n1700,
    n1701, n1702, n1703, n1704_1, n1705, n1707, n1708, n1709_1, n1711,
    n1712, n1713, n1714_1, n1715, n1716, n1717, n1718, n1719_1, n1720,
    n1721, n1722, n1723, n1724_1, n1725, n1726, n1727, n1728, n1729_1,
    n1730, n1731, n1732, n1733, n1734_1, n1735, n1736, n1737, n1738,
    n1739_1, n1740, n1741, n1742, n1743, n1745, n1746, n1747, n1748,
    n1749_1, n1750, n1751, n1752, n1753, n1754_1, n1755, n1756, n1758,
    n1760, n1762, n1764_1, n1765, n1766, n1767, n1768, n1770, n1771, n1773,
    n1775, n1777, n1778, n1779_1, n1780, n1781, n1782, n1783, n1784_1,
    n1785, n1786, n1787, n1788, n1789_1, n1790, n1791, n1792, n1793,
    n1794_1, n1795, n1796, n1797, n1798, n1799_1, n1800, n1801, n1802,
    n1803, n1804_1, n1805, n1806, n1807, n1808, n1809_1, n1810, n1811,
    n1812, n1813, n1814_1, n1815, n1817, n1818, n1820, n1822, n1823,
    n1824_1, n1826, n1827, n1828, n1830, n1831, n1832, n1834_1, n1835,
    n1837, n1838, n1839_1, n1840, n1841, n1842, n1843, n1844_1, n1845,
    n1846, n1847, n1848, n1849_1, n1850, n1851, n1852, n1853, n1854_1,
    n1855, n1856, n1857, n1858, n1859_1, n1860, n1861, n1862, n1863,
    n1864_1, n1865, n1866, n1867, n1868, n1869_1, n1870, n1871, n1872,
    n1873, n1874_1, n1875, n1876, n1877, n1878, n1879_1, n1880, n1881,
    n1882, n1883, n1884_1, n1885, n1886, n1887, n1888, n1890, n1891, n1892,
    n1893, n1895, n1897, n1899_1, n1901, n1902, n1903, n1905, n1906, n1907,
    n1908, n1909_1, n1911, n1913, n1915, n1916, n1917, n1918, n1920, n1922,
    n1923, n1924_1, n1925, n1927, n1929_1, n1931, n1932, n1933, n1934_1,
    n1935, n1936, n1937, n1938, n1940, n1941, n1942, n1943, n1945, n1946,
    n1947, n1948, n1949_1, n1950, n1951, n1952, n1953, n1954_1, n1955,
    n1956, n1957, n1958, n1959_1, n1960, n1961, n1962, n1963, n1964_1,
    n1965, n1966, n1967, n1968, n1969_1, n1970, n1971, n1972, n1973,
    n1974_1, n1975, n1976, n1977, n1978, n1979_1, n1981, n1983, n1985,
    n1988, n1989_1, n1990, n1991, n1994_1, n1995, n1996, n1997, n1998,
    n1999_1, n2000, n2001, n2002, n2003, n2004_1, n2005, n2006, n2007,
    n2008, n2009_1, n2010, n2011, n2012, n2013, n2014_1, n2015, n2016,
    n2017, n2018, n2019_1, n2020, n2021, n2022, n2023, n2024_1, n2025,
    n2026, n2027, n2028, n2029_1, n2030, n2032, n2033, n2035, n2036, n2037,
    n2039_1, n2041, n2043, n2045, n2046, n2047, n2048, n2049_1, n2050,
    n2051, n2052, n2053, n2054_1, n2055, n2056, n2057, n2058, n2059_1,
    n2060, n2061, n2062, n2063, n2064_1, n2065, n2066, n2067, n2068,
    n2069_1, n2071, n2072, n2074_1, n2075, n2076, n2078, n2080, n2081,
    n2083, n2084_1, n2086, n2088, n2089_1, n2091, n2092, n2094_1, n2095,
    n2096, n2098, n2100, n2101, n2103, n2105, n2106, n2108, n2109_1, n2110,
    n2111, n2113, n2114_1, n2115, n2116, n2117, n2119_1, n2120, n2122,
    n2123, n2124_1, n2126, n2127, n2129_1, n2130, n2131, n2133, n2134_1,
    n2135, n2137, n2139_1, n2141, n2142, n2143, n2144_1, n2146, n2147,
    n2148, n2150, n2152, n2154_1, n2156, n2158, n2160, n2162, n2163, n2165,
    n2166, n2167, n2169_1, n2170, n2171, n2172, n2173, n2174_1, n2176,
    n2178, n2179_1, n2181, n2182, n2184_1, n2185, n2186, n2187, n2188,
    n2190, n2191, n2192, n2193, n2194_1, n2196, n2197, n2198, n2199_1,
    n2200, n2201, n2202, n2203, n2204_1, n2205, n2206, n2207, n2208,
    n2209_1, n2210, n2211, n2212, n2213, n2214_1, n2215, n2216, n2217,
    n2218, n2219_1, n2220, n2221, n2222, n2223, n2224_1, n2225, n2226,
    n2227, n2228, n2229_1, n2230, n2231, n2232, n2233, n2234_1, n2235,
    n2236, n2237, n2238, n2239_1, n2240, n2241, n2242, n2243, n2244_1,
    n2245, n2246, n2248, n2249_1, n2250, n2252, n2253, n2255, n2257, n2258,
    n2260, n2261, n2263, n2264_1, n2265, n2267, n2268, n2270, n2272, n2274,
    n2276, n2278, n2279, n2280, n2281, n2282, n2284, n2285, n2287, n2289,
    n2291, n2292, n2294, n2296, n2298, n2299, n2301, n2302, n2304, n2305,
    n2306, n2309, n2311, n2312, n2313, n2315, n2317, n2318, n2320, n2322,
    n2324, n2326, n2328, n2329, n2331, n2333, n2335, n2337, n2339, n2340,
    n2341, n2343, n2345, n2347, n2348, n2350, n2352, n2354, n2356, n2358,
    n2360, n2362, n2363, n2365, n2367, n2369, n2371, n2373, n2375, n2376,
    n2377, n2379, n2380, n2381, n2383, n2384, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2394, n2396, n2398, n2400, n2402, n2403, n2404,
    n2405, n2406, n2407, n2409, n2410, n2411, n2413, n2414, n2415, n2416,
    n2417, n2419, n2421, n2423, n2425, n2426, n2428, n2430, n2432, n2433,
    n2434, n2436, n2438, n2440, n2441, n2442, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2467, n2469, n2470,
    n2472, n2474, n2475, n2477, n2479, n2481, n2483, n2484, n2486, n2488,
    n2490, n2491, n2493, n2495, n2497, n2498, n2500, n2501, n2503, n2505,
    n2506, n2507, n2509, n2510, n2511, n2512, n2513, n2514, n2516, n2518,
    n2520, n2521, n2522, n2523, n2524, n2525, n2527, n2528, n2529, n2531,
    n2533, n2534, n2535, n2536, n2537, n2538, n2540, n2542, n2543, n2545,
    n2547, n2549, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2574, n2576, n2578, n2580, n2581, n2583, n2584, n2586,
    n2588, n2590, n2592, n2593, n2595, n2596, n2598, n2599, n2600, n2602,
    n2603, n2604, n2606, n2608, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2622, n2624, n2625, n2626, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2641, n2642, n2643, n2645, n2647, n2648, n2650, n2651, n2652,
    n2653, n2654, n2655, n2657, n2658, n2659, n2661, n2663, n2664, n2666,
    n2667, n2668, n2669, n2672, n2674, n2675, n2677, n2679, n2680, n2682,
    n2684, n2685, n2687, n2689, n2691, n2692, n2694, n2696, n2697, n2699,
    n2700, n2702, n2703, n2705, n2706, n2708, n2710, n2711, n2713, n2715,
    n2717, n2718, n2720, n2722, n2723, n2725, n2727, n2728, n2729, n2731,
    n2732, n2734, n2735, n2737, n2738, n2739, n2741, n2744, n2745, n2746,
    n2747, n2748, n2750, n2751, n2753, n2754, n2756, n2757, n2759, n2761,
    n2763, n2765, n2768, n2769, n2771, n2772, n2774, n2775, n2777, n2779,
    n2781, n2782, n2784, n2786, n2787, n2789, n2790, n2791, n2793, n2794,
    n2795, n2797, n2799, n2801, n2803, n2805, n2807, n2809, n2811, n2812,
    n2814, n2816, n2818, n2819, n2820, n2821, n2822, n2823, n2825, n2827,
    n2828, n2830, n2832, n2834, n2836, n2837, n2838, n2839, n2841, n2842,
    n2843, n2845, n2846, n2848, n2850, n2852, n2854, n2856, n2858, n2860,
    n2861, n2862, n2863, n2864, n2865, n2867, n2868, n2869, n2870, n2872,
    n2873, n2875, n2876, n2878, n2879, n2881, n2882, n2883, n2885, n2886,
    n2887, n2889, n2891, n2893, n2895, n2897, n2898, n2899, n2901, n2902,
    n2904, n2906, n2907, n2908, n2910, n2912, n2913, n2914, n2915, n2916,
    n2918, n2920, n2921, n2923, n2924, n2926, n2928, n2929, n2931, n2932,
    n2933, n2935, n2936, n2937, n2939, n2941, n2943, n2944, n2946, n2948,
    n2950, n2951, n2953, n2954, n2956, n2958, n2959, n2961, n2962, n2964,
    n2965, n2966, n2968, n2969, n2970, n2972, n2973, n2975, n2976, n2978,
    n2979, n2981, n2982, n2984, n2985, n2987, n2988, n2990, n2992, n2994,
    n2995, n2996, n2998, n3000, n3001, n3003, n3005, n3006, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3019, n3021,
    n3022, n3024, n3026, n3027, n3028, n3030, n3032, n3033, n3035, n3036,
    n3038, n3039, n3040, n3042, n3043, n3045, n3047, n3049, n3051, n3053,
    n3055, n3057, n3058, n3059, n3061, n3062, n3063, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3081, n3082, n3084, n3085, n3087, n3089, n3090, n3091, n3092,
    n3093, n3094, n3096, n3097, n3099, n3100, n3101, n3102, n3103, n3104,
    n3106, n3108, n3110, n3112, n3114, n3116, n3117, n3119, n3121, n3123,
    n3125, n3127, n3129, n3130, n3131, n3132, n3133, n3134, n3136, n3138,
    n3139, n3141, n3142, n350, n355, n360, n365, n370, n375, n380, n385,
    n390, n395, n400, n405, n410, n415, n420, n425, n430, n435, n440, n445,
    n450, n455, n460, n465, n470, n475, n480, n485, n490, n495, n500, n505,
    n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560, n565,
    n570, n575, n580, n585, n590, n595, n600, n605, n610, n615, n620, n625,
    n630, n635, n640, n645, n650, n655, n660, n665, n670, n675, n680, n685,
    n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740, n745,
    n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800, n805,
    n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860, n865,
    n870, n875, n880, n885, n890, n895, n899, n904, n909, n914, n919, n924,
    n929, n934, n939, n944, n949, n954, n959, n964, n969, n974, n979, n984,
    n989, n994, n999, n1004, n1009, n1014, n1019, n1024, n1029, n1034,
    n1039, n1044, n1049, n1054, n1059, n1064, n1069, n1074, n1079, n1084,
    n1089, n1094, n1099, n1104, n1109, n1114, n1119, n1124, n1129, n1134,
    n1139, n1144, n1149, n1154, n1159, n1164, n1169, n1174, n1179, n1184,
    n1189, n1194, n1199, n1204, n1209, n1214, n1219, n1224, n1229, n1234,
    n1239, n1244, n1249, n1254, n1259, n1264, n1269, n1274, n1279, n1284,
    n1289, n1294, n1299, n1304, n1309, n1314, n1319, n1324, n1329, n1334,
    n1339, n1344, n1349, n1354, n1359, n1364, n1369, n1374, n1379, n1384,
    n1389, n1394, n1399, n1404, n1409, n1414, n1419, n1424, n1429, n1434,
    n1439, n1444, n1449, n1454, n1459, n1464, n1469, n1474, n1479, n1484,
    n1489, n1494, n1499, n1504, n1509, n1514, n1519, n1524, n1529, n1534,
    n1539, n1544, n1549, n1554, n1559, n1564, n1569, n1574, n1579, n1584,
    n1589, n1594, n1599, n1604, n1609, n1614, n1619, n1624, n1629, n1634,
    n1639, n1644, n1649, n1654, n1659, n1664, n1669, n1674, n1679, n1684,
    n1689, n1694, n1699, n1704, n1709, n1714, n1719, n1724, n1729, n1734,
    n1739, n1744, n1749, n1754, n1759, n1764, n1769, n1774, n1779, n1784,
    n1789, n1794, n1799, n1804, n1809, n1814, n1819, n1824, n1829, n1834,
    n1839, n1844, n1849, n1854, n1859, n1864, n1869, n1874, n1879, n1884,
    n1889, n1894, n1899, n1904, n1909, n1914, n1919, n1924, n1929, n1934,
    n1939, n1944, n1949, n1954, n1959, n1964, n1969, n1974, n1979, n1984,
    n1989, n1994, n1999, n2004, n2009, n2014, n2019, n2024, n2029, n2034,
    n2039, n2044, n2049, n2054, n2059, n2064, n2069, n2074, n2079, n2084,
    n2089, n2094, n2099, n2104, n2109, n2114, n2119, n2124, n2129, n2134,
    n2139, n2144, n2149, n2154, n2159, n2164, n2169, n2174, n2179, n2184,
    n2189, n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2229, n2234,
    n2239, n2244, n2249, n2254, n2259, n2264, n2269;
  assign pv14_2_2_ = n_n3358 & n_n4153;
  assign pv12_3_3_ = n_n3631 & n_n3367;
  assign n1333 = n_n4136 & n_n3042;
  assign n1334_1 = tin_pv10_4_4_ & ~n_n3042;
  assign pv10_4_4_ = n1333 | n1334_1;
  assign pv7_5_5_ = n_n3130 & n_n3679;
  assign pv3_6_6_ = n_n3252 & n_n3057;
  assign pv15_2_2_ = n_n3113 & n_n4037;
  assign pv13_3_3_ = n_n3600 & n_n3404;
  assign n1340 = n_n4120 & n_n3966;
  assign n1341 = tin_pv11_4_4_ & ~n_n4120;
  assign pv11_4_4_ = n1340 | n1341;
  assign n1343 = n_n4164 & n_n3370;
  assign n1344_1 = tin_pv6_7_7_ & ~n_n4164;
  assign pv6_7_7_ = n1343 | n1344_1;
  assign n1346 = n_n3211 & n_n3910;
  assign n1347 = tin_pv2_0_0_ & ~n_n3211;
  assign pv2_0_0_ = n1346 | n1347;
  assign pv14_1_1_ = n_n3012 & n_n3038;
  assign pv12_2_2_ = n_n3067 & n_n3576;
  assign n1351 = n_n4129 & n_n3213;
  assign n1352 = tin_pv10_3_3_ & ~n_n4129;
  assign pv10_3_3_ = n1351 | n1352;
  assign pv9_0_0_ = n_n3128 & n_n3890;
  assign pv5_1_1_ = n_n3443 & n_n3287;
  assign n1356 = n_n3470 & n_n3537;
  assign n1357 = tin_pv1_2_2_ & ~n_n3470;
  assign pv1_2_2_ = n1356 | n1357;
  assign pv15_1_1_ = n_n3606 & n_n3108;
  assign pv13_2_2_ = n_n3379 & n_n3463;
  assign n1361 = n_n3432 & n_n3583;
  assign n1362 = tin_pv11_3_3_ & ~n_n3432;
  assign pv11_3_3_ = n1361 | n1362;
  assign pv8_2_2_ = n_n3456 & n_n3055;
  assign n1365 = n_n3489 & n_n4309;
  assign n1366 = tin_pv4_3_3_ & ~n_n3489;
  assign pv4_3_3_ = n1365 | n1366;
  assign pv14_0_0_ = n_n3761 & n_n3903;
  assign pv12_1_1_ = n_n3264 & n_n4390;
  assign n1370 = n_n3549 & n_n3065;
  assign n1371 = tin_pv10_2_2_ & ~n_n3065;
  assign pv10_2_2_ = n1370 | n1371;
  assign pv7_6_6_ = n_n3670 & n_n3617;
  assign pv3_7_7_ = n_n3590 & n_n4102;
  assign pv15_0_0_ = n_n4003 & n_n3188;
  assign pv13_1_1_ = n_n3221 & n_n3150;
  assign n1377 = n_n3152 & n_n3823;
  assign n1378 = tin_pv11_2_2_ & ~n_n3152;
  assign pv11_2_2_ = n1377 | n1378;
  assign n1380 = n_n3029 & n_n3506;
  assign n1381 = tin_pv6_0_0_ & ~n_n3029;
  assign pv6_0_0_ = n1380 | n1381;
  assign n1383 = n_n3999 & n_n3646;
  assign n1384_1 = tin_pv2_1_1_ & ~n_n3999;
  assign pv2_1_1_ = n1383 | n1384_1;
  assign pv12_0_0_ = n_n3098 & n_n3339;
  assign n1387 = n_n3270 & n_n3872;
  assign n1388 = tin_pv10_1_1_ & ~n_n3872;
  assign pv10_1_1_ = n1387 | n1388;
  assign pv9_1_1_ = n_n3024 & n_n3044;
  assign pv5_2_2_ = n_n4286 & n_n3350;
  assign n1392 = n_n3441 & n_n4180;
  assign n1393 = tin_pv1_3_3_ & ~n_n3441;
  assign pv1_3_3_ = n1392 | n1393;
  assign pv13_0_0_ = n_n3061 & n_n3434;
  assign n1396 = n_n4142 & n_n4185;
  assign n1397 = tin_pv11_1_1_ & ~n_n4185;
  assign pv11_1_1_ = n1396 | n1397;
  assign pv8_3_3_ = n_n3146 & n_n3091;
  assign n1400 = n_n3627 & n_n4110;
  assign n1401 = tin_pv4_4_4_ & ~n_n4110;
  assign pv4_4_4_ = n1400 | n1401;
  assign n1403 = n_n4108 & n_n3354;
  assign n1404_1 = tin_pready_0_0_ & ~n_n4108;
  assign pready_0_0_ = n1403 | n1404_1;
  assign n1406 = n_n4282 & n_n4209;
  assign n1407 = tin_pv10_0_0_ & ~n_n4282;
  assign pv10_0_0_ = n1406 | n1407;
  assign pv7_7_7_ = n_n3136 & n_n4077;
  assign pv3_0_0_ = n_n3173 & n_n3828;
  assign n1411 = n_n3514 & n_n3233;
  assign n1412 = tin_pv11_0_0_ & ~n_n3233;
  assign pv11_0_0_ = n1411 | n1412;
  assign n1414_1 = n_n3144 & n_n3952;
  assign n1415 = tin_pv6_1_1_ & ~n_n3144;
  assign pv6_1_1_ = n1414_1 | n1415;
  assign n1417 = n_n3202 & n_n4354;
  assign n1418 = tin_pv2_2_2_ & ~n_n4354;
  assign pv2_2_2_ = n1417 | n1418;
  assign pv9_2_2_ = n_n3736 & n_n3157;
  assign pv5_3_3_ = n_n3321 & n_n4236;
  assign n1422 = n_n3863 & n_n3806;
  assign n1423 = tin_pv1_4_4_ & ~n_n3863;
  assign pv1_4_4_ = n1422 | n1423;
  assign pv8_4_4_ = n_n3344 & n_n3095;
  assign n1426 = n_n3733 & n_n3087;
  assign n1427 = tin_pv4_5_5_ & ~n_n3087;
  assign pv4_5_5_ = n1426 | n1427;
  assign pv7_0_0_ = n_n3161 & n_n3069;
  assign pv3_1_1_ = n_n3048 & n_n3461;
  assign n1431 = n_n3307 & n_n3138;
  assign n1432 = tin_pv6_2_2_ & ~n_n3307;
  assign pv6_2_2_ = n1431 | n1432;
  assign n1434_1 = n_n3465 & n_n3874;
  assign n1435 = tin_pv2_3_3_ & ~n_n3874;
  assign pv2_3_3_ = n1434_1 | n1435;
  assign pv9_3_3_ = n_n3906 & n_n3749;
  assign pv5_4_4_ = n_n3793 & n_n4213;
  assign n1439_1 = n_n3313 & n_n3101;
  assign n1440 = tin_pv1_5_5_ & ~n_n3101;
  assign pv1_5_5_ = n1439_1 | n1440;
  assign pv8_5_5_ = n_n3116 & n_n3331;
  assign n1443 = n_n3774 & n_n3413;
  assign n1444_1 = tin_pv4_6_6_ & ~n_n3774;
  assign pv4_6_6_ = n1443 | n1444_1;
  assign pv7_1_1_ = n_n3415 & n_n3971;
  assign pv3_2_2_ = n_n3190 & n_n3739;
  assign n1448 = n_n3204 & n_n3486;
  assign n1449_1 = tin_pv6_3_3_ & ~n_n3204;
  assign pv6_3_3_ = n1448 | n1449_1;
  assign n1451 = n_n3133 & n_n3643;
  assign n1452 = tin_pv2_4_4_ & ~n_n3643;
  assign pv2_4_4_ = n1451 | n1452;
  assign pv9_4_4_ = n_n3687 & n_n3650;
  assign pv5_5_5_ = n_n3266 & n_n3408;
  assign n1456 = n_n3118 & n_n4018;
  assign n1457 = tin_pv1_6_6_ & ~n_n4018;
  assign pv1_6_6_ = n1456 | n1457;
  assign pv8_6_6_ = n_n3180 & n_n3223;
  assign n1460 = n_n4114 & n_n4166;
  assign n1461 = tin_pv4_7_7_ & ~n_n4114;
  assign pv4_7_7_ = n1460 | n1461;
  assign pv7_2_2_ = n_n3497 & n_n4105;
  assign pv3_3_3_ = n_n3274 & n_n4342;
  assign n1465 = n_n3093 & n_n4065;
  assign n1466 = tin_pv6_4_4_ & ~n_n3093;
  assign pv6_4_4_ = n1465 | n1466;
  assign n1468 = n_n3780 & n_n4059;
  assign n1469_1 = tin_pv2_5_5_ & ~n_n4059;
  assign pv2_5_5_ = n1468 | n1469_1;
  assign pv14_7_7_ = n_n3449 & n_n4241;
  assign pv9_5_5_ = n_n3985 & n_n4290;
  assign pv5_6_6_ = n_n3567 & n_n3237;
  assign n1474_1 = n_n3544 & n_n4199;
  assign n1475 = tin_pv1_7_7_ & ~n_n3544;
  assign pv1_7_7_ = n1474_1 | n1475;
  assign pv15_7_7_ = n_n3079 & n_n3648;
  assign pv8_7_7_ = n_n3525 & n_n3529;
  assign n1479_1 = n_n3517 & n_n3826;
  assign n1480 = tin_pv4_0_0_ & ~n_n3826;
  assign pv4_0_0_ = n1479_1 | n1480;
  assign pv14_6_6_ = n_n3713 & n_n3262;
  assign pv12_7_7_ = n_n3764 & n_n3720;
  assign pv7_3_3_ = n_n3411 & n_n4303;
  assign pv3_4_4_ = n_n3729 & n_n4162;
  assign pv15_6_6_ = n_n4375 & n_n3020;
  assign pv13_7_7_ = n_n3372 & n_n3394;
  assign n1488 = n_n4189 & n_n3348;
  assign n1489_1 = tin_pv6_5_5_ & ~n_n3348;
  assign pv6_5_5_ = n1488 | n1489_1;
  assign n1491 = n_n3120 & n_n3385;
  assign n1492 = tin_pv2_6_6_ & ~n_n3120;
  assign pv2_6_6_ = n1491 | n1492;
  assign pv14_5_5_ = n_n3008 & n_n3663;
  assign pv12_6_6_ = n_n3782 & n_n3896;
  assign n1496 = n_n3225 & n_n3521;
  assign n1497 = tin_pv10_7_7_ & ~n_n3521;
  assign pv10_7_7_ = n1496 | n1497;
  assign pv9_6_6_ = n_n4243 & n_n3239;
  assign pv5_7_7_ = n_n3111 & n_n4005;
  assign n1501 = n_n3551 & n_n4192;
  assign n1502 = tin_pv1_0_0_ & ~n_n3551;
  assign pv1_0_0_ = n1501 | n1502;
  assign pv15_5_5_ = n_n3277 & n_n3674;
  assign pv13_6_6_ = n_n3155 & n_n3797;
  assign n1506 = n_n3376 & n_n3360;
  assign n1507 = tin_pv11_7_7_ & ~n_n3360;
  assign pv11_7_7_ = n1506 | n1507;
  assign pv8_0_0_ = n_n3014 & n_n4320;
  assign n1510 = n_n4089 & n_n3722;
  assign n1511 = tin_pv4_1_1_ & ~n_n4089;
  assign pv4_1_1_ = n1510 | n1511;
  assign pv14_4_4_ = n_n3326 & n_n3089;
  assign pv12_5_5_ = n_n3619 & n_n3337;
  assign n1515 = n_n3570 & n_n3342;
  assign n1516 = tin_pv10_6_6_ & ~n_n3570;
  assign pv10_6_6_ = n1515 | n1516;
  assign pv7_4_4_ = n_n3073 & n_n3053;
  assign pv3_5_5_ = n_n3436 & n_n3142;
  assign pv15_4_4_ = n_n3305 & n_n3667;
  assign pv13_5_5_ = n_n4139 & n_n3777;
  assign n1522 = n_n4279 & n_n3504;
  assign n1523 = tin_pv11_6_6_ & ~n_n3504;
  assign pv11_6_6_ = n1522 | n1523;
  assign n1525 = n_n3429 & n_n3836;
  assign n1526 = tin_pv6_6_6_ & ~n_n3836;
  assign pv6_6_6_ = n1525 | n1526;
  assign n1528 = n_n4131 & n_n3126;
  assign n1529_1 = tin_pv2_7_7_ & ~n_n4131;
  assign pv2_7_7_ = n1528 | n1529_1;
  assign pv14_3_3_ = n_n3396 & n_n3316;
  assign pv12_4_4_ = n_n3231 & n_n3175;
  assign n1533 = n_n3381 & n_n4247;
  assign n1534_1 = tin_pv10_5_5_ & ~n_n3381;
  assign pv10_5_5_ = n1533 | n1534_1;
  assign pv9_7_7_ = n_n3319 & n_n3040;
  assign pv5_0_0_ = n_n3195 & n_n3572;
  assign n1538 = n_n3215 & n_n3183;
  assign n1539_1 = tin_pv1_1_1_ & ~n_n3215;
  assign pv1_1_1_ = n1538 | n1539_1;
  assign pv15_3_3_ = n_n4172 & n_n3051;
  assign pv13_4_4_ = n_n3075 & n_n3758;
  assign n1543 = n_n3081 & n_n3207;
  assign n1544_1 = tin_pv11_5_5_ & ~n_n3081;
  assign pv11_5_5_ = n1543 | n1544_1;
  assign pv8_1_1_ = n_n3938 & n_n3883;
  assign n1547 = n_n4347 & n_n4372;
  assign n1548 = tin_pv4_2_2_ & ~n_n4347;
  assign pv4_2_2_ = n1547 | n1548;
  assign n1550 = ~n_n4160 & ~n_n4159;
  assign n1551 = ~n_n4383 & n1550;
  assign n1552 = ~n_n4182 & n1551;
  assign n1553 = ~n_n4330 & n1552;
  assign n1554_1 = ~n_n4224 & n1553;
  assign n1555 = ~n_n4251 & n1554_1;
  assign n1556 = n_n4251 & ~n1554_1;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = n_n4224 & ~n1553;
  assign n1559_1 = ~n1554_1 & ~n1558;
  assign n1560 = n_n4330 & ~n1552;
  assign n1561 = ~n1553 & ~n1560;
  assign n1562 = n_n4182 & ~n1551;
  assign n1563 = ~n1552 & ~n1562;
  assign n1564_1 = ~n_n4160 & n_n4222;
  assign n1565 = n_n4159 & ~n_n3976;
  assign n1566 = ~n1564_1 & n1565;
  assign n1567 = n_n4160 & ~n_n4222;
  assign n1568 = ~n1550 & ~n1567;
  assign n1569_1 = ~n1566 & n1568;
  assign n1570 = n_n4383 & ~n1550;
  assign n1571 = ~n1551 & ~n1570;
  assign n1572 = ~n1569_1 & ~n1571;
  assign n1573 = ~n_n4383 & n1569_1;
  assign n1574_1 = ~n_n4316 & ~n1573;
  assign n1575 = ~n1572 & ~n1574_1;
  assign n1576 = n1563 & n1575;
  assign n1577 = ~n1563 & ~n1575;
  assign n1578 = n_n4229 & ~n1577;
  assign n1579_1 = ~n1576 & ~n1578;
  assign n1580 = ~n1561 & n1579_1;
  assign n1581 = n1561 & ~n1579_1;
  assign n1582 = ~n_n3916 & ~n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584_1 = n1559_1 & n1583;
  assign n1585 = ~n1559_1 & ~n1583;
  assign n1586 = n_n3898 & ~n1585;
  assign n1587 = ~n1584_1 & ~n1586;
  assign n1588 = ~n1557 & n1587;
  assign n1589_1 = n1557 & ~n1587;
  assign n1590 = ~n_n4145 & ~n1589_1;
  assign n1591 = ~n1588 & ~n1590;
  assign n1592 = ~n_n4270 & ~n_n3841;
  assign n1593 = n_n4270 & n_n3841;
  assign n1594_1 = ~n1592 & ~n1593;
  assign n1595 = ~n1555 & n1594_1;
  assign n1596 = n1555 & ~n1594_1;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = n1591 & ~n1597;
  assign n1599_1 = ~n1591 & n1597;
  assign n1600 = ~n1598 & ~n1599_1;
  assign n1601 = n_n4360 & n1600;
  assign n1602 = ~n_n4360 & ~n1600;
  assign n1603 = ~n1588 & ~n1589_1;
  assign n1604_1 = n_n4145 & ~n1603;
  assign n1605 = ~n_n4145 & n1603;
  assign n1606 = ~n1604_1 & ~n1605;
  assign n1607 = n_n3898 & n1584_1;
  assign n1608 = ~n_n3898 & n1585;
  assign n1609_1 = n1587 & ~n1608;
  assign n1610 = ~n1607 & ~n1609_1;
  assign n1611 = ~n1580 & ~n1581;
  assign n1612 = n_n3916 & ~n1611;
  assign n1613 = ~n_n3916 & n1611;
  assign n1614_1 = ~n1612 & ~n1613;
  assign n1615 = n_n4229 & n1576;
  assign n1616 = ~n_n4229 & n1577;
  assign n1617 = n1579_1 & ~n1616;
  assign n1618 = ~n1615 & ~n1617;
  assign n1619_1 = ~n_n4159 & n_n3976;
  assign n1620 = ~n1565 & ~n1619_1;
  assign n1621 = ~n_n3756 & ~n1620;
  assign n1622 = n_n3743 & ~n1621;
  assign n1623 = ~n1564_1 & ~n1567;
  assign n1624_1 = ~n1565 & ~n1623;
  assign n1625 = n1565 & n1623;
  assign n1626 = ~n1624_1 & ~n1625;
  assign n1627 = ~n_n3743 & n1621;
  assign n1628 = n1626 & ~n1627;
  assign n1629_1 = ~n1622 & ~n1628;
  assign n1630 = ~n1572 & ~n1573;
  assign n1631 = ~n_n4316 & n1630;
  assign n1632 = n_n4316 & ~n1630;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634_1 = ~n_n3946 & ~n1633;
  assign n1635 = ~n1629_1 & ~n1634_1;
  assign n1636 = n_n3946 & n1633;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n_n4258 & ~n1637;
  assign n1639_1 = ~n1618 & ~n1638;
  assign n1640 = ~n_n4258 & n1637;
  assign n1641 = ~n1639_1 & ~n1640;
  assign n1642 = n_n3876 & n1641;
  assign n1643 = ~n1614_1 & ~n1642;
  assign n1644_1 = ~n_n3876 & ~n1641;
  assign n1645 = ~n1643 & ~n1644_1;
  assign n1646 = n_n4362 & n1645;
  assign n1647 = ~n1610 & ~n1646;
  assign n1648 = ~n_n4362 & ~n1645;
  assign n1649_1 = ~n1647 & ~n1648;
  assign n1650 = n_n4299 & n1649_1;
  assign n1651 = ~n1606 & ~n1650;
  assign n1652 = ~n_n4299 & ~n1649_1;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654_1 = ~n1602 & n1653;
  assign n1655 = ~n1601 & ~n1654_1;
  assign n1656 = ~n_n4067 & n1655;
  assign n1657 = ~n_n3833 & n_n4067;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659_1 = ~preset & ~pdn;
  assign n1660 = preset_0_0_ & ~nlc1_2;
  assign n1661 = nlc1_2 & ~n_n4151;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n1659_1 & n1662;
  assign n1664_1 = ~nsr1_2 & n1663;
  assign n1665 = n_n3851 & n_n4026;
  assign n1666 = ~n_n4026 & ~n1655;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = n1664_1 & ~n1667;
  assign n1669_1 = n1658 & n1668;
  assign n1670 = n_n3724 & n1669_1;
  assign n1671 = nsr1_2 & n1662;
  assign n1672 = ~pdn & ~n1671;
  assign n1673 = ~preset & ~n1672;
  assign n1674_1 = n_n4142 & n1673;
  assign n350 = n1670 | n1674_1;
  assign n1676 = ndn3_8 & ~ndn3_9;
  assign n1677 = ~n_n3936 & ~n1676;
  assign n1678 = ~pv11_1_1_ & n1676;
  assign n1679_1 = ~preset & ~n1678;
  assign n355 = ~n1677 & n1679_1;
  assign n1681 = n_n3707 & n_n3709;
  assign n1682 = ~n_n3198 & n1681;
  assign n1683 = nen3_10 & nsr3_17;
  assign n1684_1 = n_n4093 & n1658;
  assign n1685 = ~n1667 & n1684_1;
  assign n1686 = n1683 & n1685;
  assign n1687 = n_n3831 & n1686;
  assign n1688 = ~n_n4067 & n1667;
  assign n1689_1 = ~n_n3709 & ~n1688;
  assign n1690 = n1687 & n1689_1;
  assign n1691 = ~preset & ~n1690;
  assign n1692 = ~n1682 & n1691;
  assign n1693 = n_n3574 & n1692;
  assign n1694_1 = ~preset & n1682;
  assign n1695 = ~n_n3959 & ~n1620;
  assign n1696 = ~n_n3574 & ~n1626;
  assign n1697 = n_n3574 & n1626;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699_1 = n1695 & ~n1698;
  assign n1700 = ~n1695 & n1698;
  assign n1701 = ~n1699_1 & ~n1700;
  assign n1702 = n1694_1 & n1701;
  assign n1703 = ~preset & n_n3743;
  assign n1704_1 = n1690 & n1703;
  assign n1705 = ~n1702 & ~n1704_1;
  assign n360 = n1693 | ~n1705;
  assign n1707 = n_n4157 & n1664_1;
  assign n1708 = n_n3035 & n1707;
  assign n1709_1 = n_n3008 & n1673;
  assign n365 = n1708 | n1709_1;
  assign n1711 = n_n3726 & n1692;
  assign n1712 = n_n3988 & n1610;
  assign n1713 = ~n_n3988 & ~n1610;
  assign n1714_1 = n1695 & ~n1697;
  assign n1715 = ~n1696 & ~n1714_1;
  assign n1716 = ~n_n3995 & ~n1715;
  assign n1717 = n_n3995 & n1715;
  assign n1718 = ~n1633 & ~n1717;
  assign n1719_1 = ~n1716 & ~n1718;
  assign n1720 = n1618 & n1719_1;
  assign n1721 = ~n1618 & ~n1719_1;
  assign n1722 = n_n3818 & ~n1721;
  assign n1723 = ~n1720 & ~n1722;
  assign n1724_1 = ~n_n4040 & n1723;
  assign n1725 = n_n4040 & ~n1723;
  assign n1726 = ~n1614_1 & ~n1725;
  assign n1727 = ~n1724_1 & ~n1726;
  assign n1728 = ~n1713 & n1727;
  assign n1729_1 = ~n1712 & ~n1728;
  assign n1730 = ~n_n4080 & n1729_1;
  assign n1731 = n_n4080 & ~n1729_1;
  assign n1732 = ~n1606 & ~n1731;
  assign n1733 = ~n1730 & ~n1732;
  assign n1734_1 = ~n_n3726 & n1733;
  assign n1735 = n_n3726 & ~n1733;
  assign n1736 = ~n1734_1 & ~n1735;
  assign n1737 = n1600 & ~n1736;
  assign n1738 = ~n1600 & n1736;
  assign n1739_1 = n1694_1 & ~n1738;
  assign n1740 = ~n1737 & n1739_1;
  assign n1741 = ~preset & n_n4360;
  assign n1742 = n1690 & n1741;
  assign n1743 = ~n1740 & ~n1742;
  assign n370 = n1711 | ~n1743;
  assign n1745 = ~nsr3_17 & nsr3_14;
  assign n1746 = ~n_n4201 & ~n_n3533;
  assign n1747 = ~n_n3968 & ~n_n3922;
  assign n1748 = n1746 & n1747;
  assign n1749_1 = ~n_n3892 & ~n_n4337;
  assign n1750 = ~n_n4349 & ~n_n4071;
  assign n1751 = n1749_1 & n1750;
  assign n1752 = n1748 & n1751;
  assign n1753 = ~n_n3658 & ~n1752;
  assign n1754_1 = n_n4045 & n1753;
  assign n1755 = n1745 & n1754_1;
  assign n1756 = ~n_n3604 & ~n1755;
  assign n375 = ~preset & ~n1756;
  assign n1758 = ~n_n3144 & ~n1672;
  assign n380 = ~preset & ~n1758;
  assign n1760 = ~n_n3782 & ~n1672;
  assign n385 = ~preset & ~n1760;
  assign n1762 = ~n_n3067 & ~n1672;
  assign n390 = ~preset & ~n1762;
  assign n1764_1 = ndn3_7 & ~ndn3_8;
  assign n1765 = ~preset & n_n4258;
  assign n1766 = ~n1764_1 & n1765;
  assign n1767 = ~preset & n1764_1;
  assign n1768 = pv10_3_3_ & n1767;
  assign n395 = n1766 | n1768;
  assign n1770 = n_n4360 & n1664_1;
  assign n1771 = n_n3225 & n1673;
  assign n400 = n1770 | n1771;
  assign n1773 = ~n_n3180 & ~n1672;
  assign n405 = ~preset & ~n1773;
  assign n1775 = ~n_n3274 & ~n1672;
  assign n410 = ~preset & ~n1775;
  assign n1777 = n_n4057 & n_n4056;
  assign n1778 = ~n_n3557 & n1777;
  assign n1779_1 = n_n3604 & n_n3658;
  assign n1780 = ~n1753 & ~n1779_1;
  assign n1781 = n_n4045 & ~n1780;
  assign n1782 = n1745 & n1781;
  assign n1783 = ~n_n4056 & n1782;
  assign n1784_1 = ~n1778 & ~n1783;
  assign n1785 = ~preset & n1784_1;
  assign n1786 = n_n3475 & n1785;
  assign n1787 = ~preset & n1778;
  assign n1788 = ~n_n4222 & ~n_n4125;
  assign n1789_1 = n_n4222 & n_n4125;
  assign n1790 = n_n3934 & n_n3976;
  assign n1791 = ~n1789_1 & ~n1790;
  assign n1792 = ~n1788 & ~n1791;
  assign n1793 = ~n_n3901 & ~n1792;
  assign n1794_1 = n_n3901 & n1792;
  assign n1795 = ~n_n4316 & ~n1794_1;
  assign n1796 = ~n1793 & ~n1795;
  assign n1797 = ~n_n3769 & ~n1796;
  assign n1798 = n_n3769 & n1796;
  assign n1799_1 = ~n_n4229 & ~n1798;
  assign n1800 = ~n1797 & ~n1799_1;
  assign n1801 = n_n4047 & n1800;
  assign n1802 = ~n_n4047 & ~n1800;
  assign n1803 = n_n3916 & ~n1802;
  assign n1804_1 = ~n1801 & ~n1803;
  assign n1805 = n_n3898 & ~n1804_1;
  assign n1806 = ~n_n3898 & n1804_1;
  assign n1807 = n_n4366 & ~n1806;
  assign n1808 = ~n1805 & ~n1807;
  assign n1809_1 = ~n_n4145 & n1808;
  assign n1810 = n_n4145 & ~n1808;
  assign n1811 = ~n1809_1 & ~n1810;
  assign n1812 = n_n3475 & ~n1811;
  assign n1813 = ~n_n3475 & n1811;
  assign n1814_1 = ~n1812 & ~n1813;
  assign n1815 = n1787 & ~n1814_1;
  assign n415 = n1786 | n1815;
  assign n1817 = n_n3458 & n1664_1;
  assign n1818 = n_n3687 & n1673;
  assign n420 = n1817 | n1818;
  assign n1820 = ~n_n3381 & ~n1672;
  assign n425 = ~preset & ~n1820;
  assign n1822 = n_n3688 & n1664_1;
  assign n1823 = n_n3624 & n1822;
  assign n1824_1 = n_n3098 & n1673;
  assign n430 = n1823 | n1824_1;
  assign n1826 = pdn & ~ndn1_34;
  assign n1827 = ~n_n4108 & ~n1826;
  assign n1828 = ~n1672 & n1827;
  assign n435 = ~preset & ~n1828;
  assign n1830 = n1664_1 & ~n1780;
  assign n1831 = n_n3901 & n1830;
  assign n1832 = n_n3497 & n1673;
  assign n440 = n1831 | n1832;
  assign n1834_1 = ~n1614_1 & n1664_1;
  assign n1835 = n_n3793 & n1673;
  assign n445 = n1834_1 | n1835;
  assign n1837 = ~ndn3_10 & nen3_10;
  assign n1838 = ~preset & n1837;
  assign n1839_1 = nrq3_11 & ~ngfdn_3;
  assign n1840 = n_n4316 & n1839_1;
  assign n1841 = ~ndn3_15 & ngfdn_3;
  assign n1842 = n_n4211 & n_n3657;
  assign n1843 = n1841 & n1842;
  assign n1844_1 = n_n3858 & n1837;
  assign n1845 = ~n1843 & ~n1844_1;
  assign n1846 = ~n1840 & n1845;
  assign n1847 = ~n1633 & n1839_1;
  assign n1848 = ~n1780 & n1841;
  assign n1849_1 = n_n3901 & n1848;
  assign n1850 = n_n3978 & n1837;
  assign n1851 = ~n1849_1 & ~n1850;
  assign n1852 = ~n1847 & n1851;
  assign n1853 = n1846 & n1852;
  assign n1854_1 = ~n1846 & ~n1852;
  assign n1855 = ~n1853 & ~n1854_1;
  assign n1856 = n_n4125 & n1848;
  assign n1857 = n_n3328 & n1837;
  assign n1858 = ~n1626 & n1839_1;
  assign n1859_1 = ~n1857 & ~n1858;
  assign n1860 = ~n1856 & n1859_1;
  assign n1861 = n_n3934 & n1848;
  assign n1862 = n_n3931 & n1837;
  assign n1863 = ~n1620 & n1839_1;
  assign n1864_1 = ~n1862 & ~n1863;
  assign n1865 = ~n1861 & n1864_1;
  assign n1866 = n_n3688 & n_n3624;
  assign n1867 = n1841 & n1866;
  assign n1868 = n_n3878 & n1837;
  assign n1869_1 = n_n3976 & n1839_1;
  assign n1870 = ~n1868 & ~n1869_1;
  assign n1871 = ~n1867 & n1870;
  assign n1872 = ~n1865 & ~n1871;
  assign n1873 = n1860 & ~n1872;
  assign n1874_1 = ~n1860 & n1872;
  assign n1875 = n_n3099 & n1841;
  assign n1876 = n_n3936 & n1875;
  assign n1877 = n_n3208 & n1837;
  assign n1878 = n_n4222 & n1839_1;
  assign n1879_1 = ~n1877 & ~n1878;
  assign n1880 = ~n1876 & n1879_1;
  assign n1881 = ~n1874_1 & n1880;
  assign n1882 = ~n1873 & ~n1881;
  assign n1883 = ~n1855 & ~n1882;
  assign n1884_1 = n1855 & n1882;
  assign n1885 = ~n1883 & ~n1884_1;
  assign n1886 = n1838 & n1885;
  assign n1887 = ~preset & ~n1837;
  assign n1888 = n_n4316 & n1887;
  assign n450 = n1886 | n1888;
  assign n1890 = ndn3_6 & ~ndn3_7;
  assign n1891 = ~n_n4349 & ~n1890;
  assign n1892 = ~pv6_0_0_ & n1890;
  assign n1893 = ~preset & ~n1892;
  assign n455 = ~n1891 & n1893;
  assign n1895 = ~n_n3029 & ~n1672;
  assign n460 = ~preset & ~n1895;
  assign n1897 = ~n_n3619 & ~n1672;
  assign n465 = ~preset & ~n1897;
  assign n1899_1 = ~n_n3264 & ~n1672;
  assign n470 = ~preset & ~n1899_1;
  assign n1901 = n_n4288 & n1664_1;
  assign n1902 = ~n1708 & ~n1901;
  assign n1903 = n_n3780 & n1673;
  assign n475 = ~n1902 | n1903;
  assign n1905 = nsr3_3 & ~pready_0_0_;
  assign n1906 = nsr3_3 & ~n1671;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~ndn3_4 & ~n1907;
  assign n1909_1 = ~preset & ~ngfdn_3;
  assign n480 = ~n1908 & n1909_1;
  assign n1911 = ~n_n4114 & ~n1672;
  assign n485 = ~preset & ~n1911;
  assign n1913 = ~n_n3146 & ~n1672;
  assign n490 = ~preset & ~n1913;
  assign n1915 = ~ndn3_4 & n1907;
  assign n1916 = ~pv1_5_5_ & n1915;
  assign n1917 = ~n_n3511 & ~n1915;
  assign n1918 = ~preset & ~n1917;
  assign n495 = ~n1916 & n1918;
  assign n1920 = ~n_n3152 & ~n1672;
  assign n500 = ~preset & ~n1920;
  assign n1922 = ~n_n4067 & n1686;
  assign n1923 = n_n3833 & ~n1922;
  assign n1924_1 = ~n1655 & n1922;
  assign n1925 = ~preset & ~n1924_1;
  assign n505 = n1923 | ~n1925;
  assign n1927 = ~n_n4282 & ~n1672;
  assign n510 = ~preset & ~n1927;
  assign n1929_1 = ~n_n3305 & ~n1672;
  assign n515 = ~preset & ~n1929_1;
  assign n1931 = ~preset & ~n1841;
  assign n1932 = n_n4392 & n1931;
  assign n1933 = ~preset & n1841;
  assign n1934_1 = ~n1873 & ~n1874_1;
  assign n1935 = ~n1880 & ~n1934_1;
  assign n1936 = n1880 & n1934_1;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = n1933 & ~n1937;
  assign n520 = n1932 | n1938;
  assign n1940 = ndn3_5 & ~ndn3_6;
  assign n1941 = ~n_n4224 & ~n1940;
  assign n1942 = ~pv4_5_5_ & n1940;
  assign n1943 = ~preset & ~n1942;
  assign n525 = ~n1941 & n1943;
  assign n1945 = ~n1730 & ~n1731;
  assign n1946 = n1606 & ~n1945;
  assign n1947 = ~n1712 & ~n1713;
  assign n1948 = n1727 & n1947;
  assign n1949_1 = ~n1727 & ~n1947;
  assign n1950 = ~n1948 & ~n1949_1;
  assign n1951 = ~n1724_1 & ~n1725;
  assign n1952 = n1614_1 & ~n1951;
  assign n1953 = ~n1716 & ~n1717;
  assign n1954_1 = n1633 & ~n1953;
  assign n1955 = n1695 & ~n1696;
  assign n1956 = ~n_n3574 & n1620;
  assign n1957 = ~n1697 & ~n1956;
  assign n1958 = ~n1955 & n1957;
  assign n1959_1 = n1953 & ~n1958;
  assign n1960 = ~n1954_1 & ~n1959_1;
  assign n1961 = ~n1618 & n1960;
  assign n1962 = n_n3818 & n1720;
  assign n1963 = ~n_n3818 & n1721;
  assign n1964_1 = n1723 & ~n1963;
  assign n1965 = ~n1962 & ~n1964_1;
  assign n1966 = n1618 & ~n1960;
  assign n1967 = n1965 & ~n1966;
  assign n1968 = ~n1961 & ~n1967;
  assign n1969_1 = n1951 & n1968;
  assign n1970 = ~n1952 & ~n1969_1;
  assign n1971 = ~n1610 & n1970;
  assign n1972 = n1950 & ~n1971;
  assign n1973 = n1610 & ~n1970;
  assign n1974_1 = ~n1972 & ~n1973;
  assign n1975 = n1945 & ~n1974_1;
  assign n1976 = ~n1946 & ~n1975;
  assign n1977 = ~n1736 & n1976;
  assign n1978 = ~n1738 & ~n1977;
  assign n1979_1 = n1682 & ~n1978;
  assign n530 = ~preset & n1979_1;
  assign n1981 = ~n_n3204 & ~n1672;
  assign n535 = ~preset & ~n1981;
  assign n1983 = ~n_n3024 & ~n1672;
  assign n540 = ~preset & ~n1983;
  assign n1985 = ~n_n4139 & ~n1672;
  assign n545 = ~preset & ~n1985;
  assign n550 = ndn3_15 & n1909_1;
  assign n1988 = n_n4074 & n1664_1;
  assign n1989_1 = n_n3578 & n1988;
  assign n1990 = ~n1817 & ~n1989_1;
  assign n1991 = n_n3133 & n1673;
  assign n555 = ~n1990 | n1991;
  assign n2039 = ~preset & n1839_1;
  assign n1994_1 = ~n1614_1 & n1839_1;
  assign n1995 = n_n4047 & n1848;
  assign n1996 = n_n4021 & n1837;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n1994_1 & n1997;
  assign n1999_1 = n_n3916 & n1839_1;
  assign n2000 = n_n3886 & n1837;
  assign n2001 = n_n4074 & n_n3578;
  assign n2002 = n1841 & n2001;
  assign n2003 = ~n2000 & ~n2002;
  assign n2004_1 = ~n1999_1 & n2003;
  assign n2005 = ~n1998 & ~n2004_1;
  assign n2006 = n1998 & n2004_1;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = n_n3085 & n_n3250;
  assign n2009_1 = n1841 & n2008;
  assign n2010 = n_n4229 & n1839_1;
  assign n2011 = n_n4294 & n1837;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n2009_1 & n2012;
  assign n2014_1 = ~n1618 & n1839_1;
  assign n2015 = n_n3769 & n1848;
  assign n2016 = n_n3281 & n1837;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n2014_1 & n2017;
  assign n2019_1 = ~n2013 & ~n2018;
  assign n2020 = n2013 & n2018;
  assign n2021 = ~n1853 & n1882;
  assign n2022 = ~n1854_1 & ~n2021;
  assign n2023 = ~n2020 & ~n2022;
  assign n2024_1 = ~n2019_1 & ~n2023;
  assign n2025 = ~n2007 & ~n2024_1;
  assign n2026 = n2007 & n2024_1;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = n2039 & ~n2027;
  assign n2029_1 = ~preset & ~n1839_1;
  assign n2030 = n_n4074 & n2029_1;
  assign n560 = n2028 | n2030;
  assign n2032 = n_n3743 & n1664_1;
  assign n2033 = n_n3270 & n1673;
  assign n565 = n2032 | n2033;
  assign n2035 = ~pv1_2_2_ & n1915;
  assign n2036 = ~n_n3858 & ~n1915;
  assign n2037 = ~preset & ~n2036;
  assign n570 = ~n2035 & n2037;
  assign n2039_1 = ~n_n3456 & ~n1672;
  assign n575 = ~preset & ~n2039_1;
  assign n2041 = ~n_n3521 & ~n1672;
  assign n580 = ~preset & ~n2041;
  assign n2043 = ~n_n3081 & ~n1672;
  assign n585 = ~preset & ~n2043;
  assign n2045 = n_n4045 & ~n1745;
  assign n2046 = n1780 & ~n2045;
  assign n2047 = ~n_n3493 & n2046;
  assign n2048 = ~n1783 & ~n2047;
  assign n2049_1 = n_n3892 & ~n2048;
  assign n2050 = ~n_n3955 & n_n3954;
  assign n2051 = ~n_n3845 & n2050;
  assign n2052 = ~n_n4029 & n2051;
  assign n2053 = ~n_n3865 & n2052;
  assign n2054_1 = ~n_n4052 & n2053;
  assign n2055 = ~n_n4381 & n2054_1;
  assign n2056 = n_n4381 & ~n2054_1;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = n1778 & ~n2057;
  assign n2059_1 = ~n2049_1 & ~n2058;
  assign n2060 = ~n1781 & ~n2045;
  assign n2061 = ~n_n3493 & n2060;
  assign n2062 = n1784_1 & ~n2061;
  assign n2063 = ~preset & ~n2062;
  assign n2064_1 = ~n2059_1 & n2063;
  assign n2065 = ~n_n3493 & ~n1780;
  assign n2066 = ~n_n4045 & n2065;
  assign n2067 = ~n2062 & ~n2066;
  assign n2068 = ~preset & ~n2067;
  assign n2069_1 = n_n4381 & n2068;
  assign n590 = n2064_1 | n2069_1;
  assign n2071 = n_n3475 & n1830;
  assign n2072 = n_n3670 & n1673;
  assign n595 = n2071 | n2072;
  assign n2074_1 = ~n_n4211 & ~n1676;
  assign n2075 = ~pv11_2_2_ & n1676;
  assign n2076 = ~preset & ~n2075;
  assign n600 = ~n2074_1 & n2076;
  assign n2078 = ~preset & ~n2060;
  assign n605 = n_n3493 & n2078;
  assign n2080 = n1885 & n1933;
  assign n2081 = n_n3495 & n1931;
  assign n610 = n2080 | n2081;
  assign n2083 = n_n3916 & n1887;
  assign n2084_1 = n1838 & ~n2027;
  assign n615 = n2083 | n2084_1;
  assign n2086 = ~n_n3195 & ~n1672;
  assign n620 = ~preset & ~n2086;
  assign n2088 = n_n3242 & n1664_1;
  assign n2089_1 = n_n3525 & n1673;
  assign n625 = n2088 | n2089_1;
  assign n2091 = n_n3916 & n1664_1;
  assign n2092 = n_n3729 & n1673;
  assign n630 = n2091 | n2092;
  assign n2094_1 = ~preset & n_n3876;
  assign n2095 = ~n1764_1 & n2094_1;
  assign n2096 = pv10_4_4_ & n1767;
  assign n635 = n2095 | n2096;
  assign n2098 = ~ndn3_4 & ~ndn3_5;
  assign n640 = n1909_1 & ~n2098;
  assign n2100 = n_n3946 & n1664_1;
  assign n2101 = n_n3549 & n1673;
  assign n645 = n2100 | n2101;
  assign n2103 = ~n_n3489 & ~n1672;
  assign n650 = ~preset & ~n2103;
  assign n2105 = n_n3170 & n2088;
  assign n2106 = n_n3764 & n1673;
  assign n655 = n2105 | n2106;
  assign n2108 = ndn3_4 & ~ndn3_5;
  assign n2109_1 = ~n_n3281 & ~n2108;
  assign n2110 = ~pv2_3_3_ & n2108;
  assign n2111 = ~preset & ~n2110;
  assign n660 = ~n2109_1 & n2111;
  assign n2113 = n_n3707 & ~n1979_1;
  assign n2114_1 = n_n4093 & ~n1683;
  assign n2115 = n1684_1 & ~n1688;
  assign n2116 = ~n2114_1 & ~n2115;
  assign n2117 = ~preset & ~n2116;
  assign n665 = n2113 | ~n2117;
  assign n2119_1 = n_n4159 & n1664_1;
  assign n2120 = n_n3517 & n1673;
  assign n670 = n2119_1 | n2120;
  assign n2122 = ~n_n4160 & ~n1940;
  assign n2123 = ~pv4_1_1_ & n1940;
  assign n2124_1 = ~preset & ~n2123;
  assign n675 = ~n2122 & n2124_1;
  assign n2126 = n_n4222 & n1887;
  assign n2127 = n1838 & ~n1937;
  assign n680 = n2126 | n2127;
  assign n2129_1 = n_n3099 & n1664_1;
  assign n2130 = n_n3936 & n2129_1;
  assign n2131 = n_n3012 & n1673;
  assign n685 = n2130 | n2131;
  assign n2133 = ~n_n4071 & ~n1890;
  assign n2134_1 = ~pv6_5_5_ & n1890;
  assign n2135 = ~preset & ~n2134_1;
  assign n690 = ~n2133 & n2135;
  assign n2137 = ~n_n3372 & ~n1672;
  assign n695 = ~preset & ~n2137;
  assign n2139_1 = n_n3344 & n1673;
  assign n700 = n1988 | n2139_1;
  assign n2141 = n1865 & n1871;
  assign n2142 = ~n1872 & ~n2141;
  assign n2143 = n2039 & n2142;
  assign n2144_1 = n_n3688 & n2029_1;
  assign n705 = n2143 | n2144_1;
  assign n2146 = n_n4233 & n1664_1;
  assign n2147 = ~n2105 & ~n2146;
  assign n2148 = n_n3079 & n1673;
  assign n710 = ~n2147 | n2148;
  assign n2150 = n_n3313 & n1673;
  assign n715 = n1708 | n2150;
  assign n2152 = ~n_n3411 & ~n1672;
  assign n720 = ~preset & ~n2152;
  assign n2154_1 = n_n3231 & n1673;
  assign n725 = n1989_1 | n2154_1;
  assign n2156 = ~n_n3396 & ~n1672;
  assign n730 = ~preset & ~n2156;
  assign n2158 = ~n_n3432 & ~n1672;
  assign n735 = ~preset & ~n2158;
  assign n2160 = ~n_n3606 & ~n1672;
  assign n740 = ~preset & ~n2160;
  assign n2162 = n_n4224 & n1664_1;
  assign n2163 = n_n3733 & n1673;
  assign n745 = n2162 | n2163;
  assign n2165 = ~n_n3556 & ~n1676;
  assign n2166 = ~pv11_6_6_ & n1676;
  assign n2167 = ~preset & ~n2166;
  assign n750 = ~n2165 & n2167;
  assign n2169_1 = n_n4040 & n1692;
  assign n2170 = ~n1614_1 & n1951;
  assign n2171 = ~n1952 & ~n2170;
  assign n2172 = n1694_1 & ~n2171;
  assign n2173 = n1690 & n2094_1;
  assign n2174_1 = ~n2172 & ~n2173;
  assign n755 = n2169_1 | ~n2174_1;
  assign n2176 = ~n_n3120 & ~n1672;
  assign n760 = ~preset & ~n2176;
  assign n2178 = n_n4222 & n1664_1;
  assign n2179_1 = n_n3221 & n1673;
  assign n765 = n2178 | n2179_1;
  assign n2181 = n_n3976 & n1664_1;
  assign n2182 = n_n3173 & n1673;
  assign n770 = n2181 | n2182;
  assign n2184_1 = ~preset & n_n3851;
  assign n2185 = n1683 & n2115;
  assign n2186 = ~preset & n2185;
  assign n2187 = n_n3831 & n1666;
  assign n2188 = n2186 & n2187;
  assign n775 = n2184_1 | n2188;
  assign n2190 = n_n3657 & n1664_1;
  assign n2191 = n_n4211 & n2190;
  assign n2192 = n_n3495 & n1664_1;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194_1 = n_n3113 & n1673;
  assign n780 = ~n2193 | n2194_1;
  assign n2196 = ~n1606 & n1839_1;
  assign n2197 = n_n3475 & n1848;
  assign n2198 = n_n4062 & n1837;
  assign n2199_1 = ~n2197 & ~n2198;
  assign n2200 = ~n2196 & n2199_1;
  assign n2201 = n_n4145 & n1839_1;
  assign n2202 = n_n3556 & n_n4122;
  assign n2203 = n1841 & n2202;
  assign n2204_1 = n_n3919 & n1837;
  assign n2205 = ~n2203 & ~n2204_1;
  assign n2206 = ~n2201 & n2205;
  assign n2207 = ~n2200 & ~n2206;
  assign n2208 = n2200 & n2206;
  assign n2209_1 = ~n1610 & n1839_1;
  assign n2210 = n_n4366 & n1848;
  assign n2211 = n_n3854 & n1837;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2209_1 & n2212;
  assign n2214_1 = n_n3511 & n1837;
  assign n2215 = n_n3898 & n1839_1;
  assign n2216 = n_n3035 & n_n4157;
  assign n2217 = n1841 & n2216;
  assign n2218 = ~n2215 & ~n2217;
  assign n2219_1 = ~n2214_1 & n2218;
  assign n2220 = n2213 & n2219_1;
  assign n2221 = ~n2213 & ~n2219_1;
  assign n2222 = ~n2005 & n2024_1;
  assign n2223 = ~n2006 & ~n2222;
  assign n2224_1 = ~n2221 & ~n2223;
  assign n2225 = ~n2220 & ~n2224_1;
  assign n2226 = ~n2208 & n2225;
  assign n2227 = ~n2207 & ~n2226;
  assign n2228 = ~n1600 & n1839_1;
  assign n2229_1 = n_n4324 & n1848;
  assign n2230 = n_n3451 & n1837;
  assign n2231 = ~n2229_1 & ~n2230;
  assign n2232 = ~n2228 & n2231;
  assign n2233 = n_n3242 & n_n3170;
  assign n2234_1 = n1841 & n2233;
  assign n2235 = n_n3841 & n1839_1;
  assign n2236 = n_n3259 & n1837;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n2234_1 & n2237;
  assign n2239_1 = ~n2232 & n2238;
  assign n2240 = n2232 & ~n2238;
  assign n2241 = ~n2239_1 & ~n2240;
  assign n2242 = n2227 & n2241;
  assign n2243 = ~n2227 & ~n2241;
  assign n2244_1 = ~n2242 & ~n2243;
  assign n2245 = n2039 & n2244_1;
  assign n2246 = n_n3242 & n2029_1;
  assign n785 = n2245 | n2246;
  assign n2248 = n_n4122 & n1664_1;
  assign n2249_1 = n_n3556 & n2248;
  assign n2250 = n_n3118 & n1673;
  assign n790 = n2249_1 | n2250;
  assign n2252 = n_n3483 & n1669_1;
  assign n2253 = n_n3376 & n1673;
  assign n795 = n2252 | n2253;
  assign n2255 = ~n_n4089 & ~n1672;
  assign n800 = ~preset & ~n2255;
  assign n2257 = n_n4392 & n1664_1;
  assign n2258 = n_n3044 & n1673;
  assign n805 = n2257 | n2258;
  assign n2260 = n_n4330 & n1664_1;
  assign n2261 = n_n3627 & n1673;
  assign n810 = n2260 | n2261;
  assign n2263 = ~n_n3035 & ~n1676;
  assign n2264_1 = ~pv11_5_5_ & n1676;
  assign n2265 = ~preset & ~n2264_1;
  assign n815 = ~n2263 & n2265;
  assign n2267 = ~n1600 & n1664_1;
  assign n2268 = n_n3111 & n1673;
  assign n820 = n2267 | n2268;
  assign n2270 = ~n_n3321 & ~n1672;
  assign n825 = ~preset & ~n2270;
  assign n2272 = ~n_n3443 & ~n1672;
  assign n830 = ~preset & ~n2272;
  assign n2274 = ~n_n3215 & ~n1672;
  assign n835 = ~preset & ~n2274;
  assign n2276 = ~ndn3_10 & ~nen3_10;
  assign n840 = n1909_1 & ~n2276;
  assign n2278 = n_n4351 & n1664_1;
  assign n2279 = n_n3085 & n1664_1;
  assign n2280 = n_n3250 & n2279;
  assign n2281 = ~n2278 & ~n2280;
  assign n2282 = n_n4172 & n1673;
  assign n845 = ~n2281 | n2282;
  assign n2284 = ~preset_0_0_ & nsr1_2;
  assign n2285 = ~nlc1_2 & ~n2284;
  assign n850 = n1659_1 & ~n2285;
  assign n2287 = ~n_n3590 & ~n1672;
  assign n855 = ~preset & ~n2287;
  assign n2289 = ~n_n4110 & ~n1672;
  assign n860 = ~preset & ~n2289;
  assign n2291 = n1671 & n1905;
  assign n2292 = ~nlc3_3 & ~n2291;
  assign n865 = n1659_1 & ~n2292;
  assign n2294 = n_n3576 & n1673;
  assign n870 = n2191 | n2294;
  assign n2296 = ~n_n4129 & ~n1672;
  assign n875 = ~preset & ~n2296;
  assign n2298 = n_n4071 & n1664_1;
  assign n2299 = n_n4189 & n1673;
  assign n880 = n2298 | n2299;
  assign n2301 = ~n1633 & n1664_1;
  assign n2302 = n_n4286 & n1673;
  assign n885 = n2301 | n2302;
  assign n2304 = ~n_n4383 & ~n1940;
  assign n2305 = ~pv4_2_2_ & n1940;
  assign n2306 = ~preset & ~n2305;
  assign n890 = ~n2304 & n2306;
  assign n895 = ~preset & n1672;
  assign n2309 = ~n_n3567 & ~n1672;
  assign n899 = ~preset & ~n2309;
  assign n2311 = ~n_n3892 & ~n1890;
  assign n2312 = ~pv6_6_6_ & n1890;
  assign n2313 = ~preset & ~n2312;
  assign n904 = ~n2311 & n2313;
  assign n2315 = ~n_n3075 & ~n1672;
  assign n909 = ~preset & ~n2315;
  assign n2317 = ~preset & n_n3354;
  assign n2318 = ~n1826 & n2317;
  assign n914 = n895 | n2318;
  assign n2320 = n_n3465 & n1673;
  assign n919 = ~n2281 | n2320;
  assign n2322 = ~ndn3_5 & ~ndn3_6;
  assign n924 = n1909_1 & ~n2322;
  assign n2324 = ~n_n3617 & ~n1672;
  assign n929 = ~preset & ~n2324;
  assign n2326 = ~n_n4162 & ~n1672;
  assign n934 = ~preset & ~n2326;
  assign n2328 = n_n4012 & n1669_1;
  assign n2329 = n_n3207 & n1673;
  assign n939 = n2328 | n2329;
  assign n2331 = ~n_n4120 & ~n1672;
  assign n944 = ~preset & ~n2331;
  assign n2333 = ~n_n3065 & ~n1672;
  assign n949 = ~preset & ~n2333;
  assign n2335 = ~n_n4005 & ~n1672;
  assign n954 = ~preset & ~n2335;
  assign n2337 = ~n_n3266 & ~n1672;
  assign n959 = ~preset & ~n2337;
  assign n2339 = ~n_n4337 & ~n1890;
  assign n2340 = ~pv6_7_7_ & n1890;
  assign n2341 = ~preset & ~n2340;
  assign n964 = ~n2339 & n2341;
  assign n2343 = ~n_n3600 & ~n1672;
  assign n969 = ~preset & ~n2343;
  assign n2345 = ~n_n3415 & ~n1672;
  assign n974 = ~preset & ~n2345;
  assign n2347 = n_n4095 & n1664_1;
  assign n2348 = n_n4243 & n1673;
  assign n979 = n2347 | n2348;
  assign n2350 = ~n_n3872 & ~n1672;
  assign n984 = ~preset & ~n2350;
  assign n2352 = ~n_n3648 & ~n1672;
  assign n989 = ~preset & ~n2352;
  assign n2354 = n_n3358 & n1673;
  assign n994 = n2191 | n2354;
  assign n2356 = ~n_n3350 & ~n1672;
  assign n999 = ~preset & ~n2356;
  assign n2358 = ~ndn3_6 & ~ndn3_7;
  assign n1004 = n1909_1 & ~n2358;
  assign n2360 = ~n_n3116 & ~n1672;
  assign n1009 = ~preset & ~n2360;
  assign n2362 = n_n3766 & n1669_1;
  assign n2363 = n_n3583 & n1673;
  assign n1014 = n2362 | n2363;
  assign n2365 = n_n3906 & n1673;
  assign n1019 = n2278 | n2365;
  assign n2367 = ~n_n4131 & ~n1672;
  assign n1024 = ~preset & ~n2367;
  assign n2369 = n_n3316 & n1673;
  assign n1029 = n2280 | n2369;
  assign n2371 = n_n3061 & n1673;
  assign n1034 = n2181 | n2371;
  assign n2373 = n_n3048 & n1673;
  assign n1039 = n2178 | n2373;
  assign n2375 = ~pv1_4_4_ & n1915;
  assign n2376 = ~n_n3886 & ~n1915;
  assign n2377 = ~preset & ~n2376;
  assign n1044 = ~n2375 & n2377;
  assign n2379 = ~pv1_6_6_ & n1915;
  assign n2380 = ~n_n3919 & ~n1915;
  assign n2381 = ~preset & ~n2380;
  assign n1049 = ~n2379 & n2381;
  assign n2383 = n_n3608 & n1664_1;
  assign n2384 = n_n3128 & n1673;
  assign n1054 = n2383 | n2384;
  assign n2386 = n_n3995 & n1692;
  assign n2387 = ~preset & n_n3946;
  assign n2388 = n1690 & n2387;
  assign n2389 = ~n1633 & n1953;
  assign n2390 = ~n1954_1 & ~n2389;
  assign n2391 = n1694_1 & ~n2390;
  assign n2392 = ~n2388 & ~n2391;
  assign n1059 = n2386 | ~n2392;
  assign n2394 = ~n_n4213 & ~n1672;
  assign n1064 = ~preset & ~n2394;
  assign n2396 = n_n3761 & n1673;
  assign n1069 = n1823 | n2396;
  assign n2398 = ~ndn3_7 & ~ndn3_8;
  assign n1074 = n1909_1 & ~n2398;
  assign n2400 = ~n_n3252 & ~n1672;
  assign n1079 = ~preset & ~n2400;
  assign n2402 = n_n4366 & n1785;
  assign n2403 = ~n1805 & n1807;
  assign n2404 = ~n1805 & ~n1806;
  assign n2405 = ~n_n4366 & ~n2404;
  assign n2406 = n1787 & ~n2405;
  assign n2407 = ~n2403 & n2406;
  assign n1084 = n2402 | n2407;
  assign n2409 = ~n_n3328 & ~n2108;
  assign n2410 = ~pv2_1_1_ & n2108;
  assign n2411 = ~preset & ~n2410;
  assign n1089 = ~n2409 & n2411;
  assign n2413 = n_n3988 & n1692;
  assign n2414 = ~preset & n_n4362;
  assign n2415 = n1690 & n2414;
  assign n2416 = n1694_1 & n1950;
  assign n2417 = ~n2415 & ~n2416;
  assign n1094 = n2413 | ~n2417;
  assign n2419 = ~n_n3348 & ~n1672;
  assign n1099 = ~preset & ~n2419;
  assign n2421 = ~n_n3544 & ~n1672;
  assign n1104 = ~preset & ~n2421;
  assign n2423 = ~n_n3101 & ~n1672;
  assign n1109 = ~preset & ~n2423;
  assign n2425 = n_n4334 & n1669_1;
  assign n2426 = n_n4279 & n1673;
  assign n1114 = n2425 | n2426;
  assign n2428 = n_n3896 & n1673;
  assign n1119 = n2249_1 | n2428;
  assign n2430 = n_n3736 & n1673;
  assign n1124 = n2192 | n2430;
  assign n2432 = ~n_n4251 & ~n1940;
  assign n2433 = ~pv4_6_6_ & n1940;
  assign n2434 = ~preset & ~n2433;
  assign n1129 = ~n2432 & n2434;
  assign n2436 = ~n_n3650 & ~n1672;
  assign n1134 = ~preset & ~n2436;
  assign n2438 = ~n_n3307 & ~n1672;
  assign n1139 = ~preset & ~n2438;
  assign n2440 = ~pv1_3_3_ & n1915;
  assign n2441 = ~n_n4294 & ~n1915;
  assign n2442 = ~preset & ~n2441;
  assign n1144 = ~n2440 & n2442;
  assign n2444 = n_n3724 & n_n3814;
  assign n2445 = n_n4227 & n2444;
  assign n2446 = n_n3766 & n2445;
  assign n2447 = n_n4275 & n2446;
  assign n2448 = n_n4012 & n1694_1;
  assign n2449 = n2447 & n2448;
  assign n2450 = ~n_n4334 & ~n2449;
  assign n2451 = ~n_n4012 & n1694_1;
  assign n2452 = ~n1691 & ~n1694_1;
  assign n2453 = n1682 & n2447;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = n_n4334 & ~n2454;
  assign n2456 = ~n2451 & n2455;
  assign n1149 = ~n2450 & ~n2456;
  assign n2458 = n_n4201 & ~n2048;
  assign n2459 = n1778 & n2050;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = n2063 & ~n2460;
  assign n2462 = ~n_n3954 & n1778;
  assign n2463 = n2067 & ~n2462;
  assign n2464 = ~preset & n_n3955;
  assign n2465 = ~n2463 & n2464;
  assign n1154 = n2461 | n2465;
  assign n2467 = ~n_n4164 & ~n1672;
  assign n1159 = ~preset & ~n2467;
  assign n2469 = n_n4145 & n1664_1;
  assign n2470 = n_n3155 & n1673;
  assign n1164 = n2469 | n2470;
  assign n2472 = ~n_n3749 & ~n1672;
  assign n1169 = ~preset & ~n2472;
  assign n2474 = n1933 & n2244_1;
  assign n2475 = n_n4233 & n1931;
  assign n1174 = n2474 | n2475;
  assign n2477 = ~n_n4347 & ~n1672;
  assign n1179 = ~preset & ~n2477;
  assign n2479 = ~n_n3826 & ~n1672;
  assign n1184 = ~preset & ~n2479;
  assign n2481 = ~n_n3360 & ~n1672;
  assign n1189 = ~preset & ~n2481;
  assign n2483 = n_n3458 & n1931;
  assign n2484 = n1933 & ~n2027;
  assign n1194 = n2483 | n2484;
  assign n2486 = ~n_n3093 & ~n1672;
  assign n1199 = ~preset & ~n2486;
  assign n2488 = ~n_n3157 & ~n1672;
  assign n1204 = ~preset & ~n2488;
  assign n2490 = n_n4349 & n1664_1;
  assign n2491 = n_n3506 & n1673;
  assign n1209 = n2490 | n2491;
  assign n2493 = ~n_n3161 & ~n1672;
  assign n1214 = ~preset & ~n2493;
  assign n2495 = n_n3319 & n1673;
  assign n1219 = n2146 | n2495;
  assign n2497 = n_n3892 & n1664_1;
  assign n2498 = n_n3429 & n1673;
  assign n1224 = n2497 | n2498;
  assign n2500 = n_n4125 & n1830;
  assign n2501 = n_n3971 & n1673;
  assign n1229 = n2500 | n2501;
  assign n2503 = n_n3449 & n1673;
  assign n1234 = n2105 | n2503;
  assign n2505 = ~n_n4270 & ~n1940;
  assign n2506 = ~pv4_7_7_ & n1940;
  assign n2507 = ~preset & ~n2506;
  assign n1239 = ~n2505 & n2507;
  assign n2509 = ~n2220 & ~n2221;
  assign n2510 = n2223 & ~n2509;
  assign n2511 = ~n2223 & n2509;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = n1933 & ~n2512;
  assign n2514 = n_n4288 & n1931;
  assign n1244 = n2513 | n2514;
  assign n2516 = n_n3183 & n1673;
  assign n1249 = n2130 | n2516;
  assign n2518 = ~n_n3130 & ~n1672;
  assign n1254 = ~preset & ~n2518;
  assign n2520 = n_n4047 & n1785;
  assign n2521 = n_n3916 & n1801;
  assign n2522 = ~n_n3916 & n1802;
  assign n2523 = n1804_1 & ~n2522;
  assign n2524 = ~n2521 & ~n2523;
  assign n2525 = n1787 & ~n2524;
  assign n1264 = n2520 | n2525;
  assign n2527 = ~n_n3978 & ~n2108;
  assign n2528 = ~pv2_2_2_ & n2108;
  assign n2529 = ~preset & ~n2528;
  assign n1269 = ~n2527 & n2529;
  assign n2531 = ~n_n3239 & ~n1672;
  assign n1274 = ~preset & ~n2531;
  assign n2533 = ~n2207 & ~n2208;
  assign n2534 = ~n2225 & ~n2533;
  assign n2535 = n2225 & n2533;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = n1838 & n2536;
  assign n2538 = n_n4145 & n1887;
  assign n1279 = n2537 | n2538;
  assign n2540 = ~n_n3890 & ~n1672;
  assign n1284 = ~preset & ~n2540;
  assign n2542 = ~n1823 & ~n2383;
  assign n2543 = n_n4003 & n1673;
  assign n1289 = ~n2542 | n2543;
  assign n2545 = n_n3091 & n1673;
  assign n1294 = n2279 | n2545;
  assign n2547 = n_n3985 & n1673;
  assign n1299 = n1901 | n2547;
  assign n2549 = ~n_n3326 & ~n1672;
  assign n1304 = ~preset & ~n2549;
  assign n2551 = n1778 & n2054_1;
  assign n2552 = n1778 & ~n2053;
  assign n2553 = ~n2066 & ~n2552;
  assign n2554 = n_n4052 & ~n2553;
  assign n2555 = n_n4071 & ~n2048;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2551 & n2556;
  assign n2558 = n2063 & ~n2557;
  assign n2559 = n1785 & ~n2061;
  assign n2560 = n_n4052 & n2559;
  assign n1309 = n2558 | n2560;
  assign n1314 = nsr4_2 | ~n1659_1;
  assign n2563 = n_n4099 & n2559;
  assign n2564 = ~n_n4099 & n2551;
  assign n2565 = ~n_n4381 & n2564;
  assign n2566 = n1778 & ~n2055;
  assign n2567 = ~n2066 & ~n2566;
  assign n2568 = n_n4099 & ~n2567;
  assign n2569 = n_n4337 & ~n2048;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2565 & n2570;
  assign n2572 = n2063 & ~n2571;
  assign n1319 = n2563 | n2572;
  assign n2574 = ~n_n4375 & ~n1672;
  assign n1324 = ~preset & ~n2574;
  assign n2576 = ~n_n4067 & ~n1686;
  assign n1329 = n2117 & ~n2576;
  assign n2578 = ~n_n4290 & ~n1672;
  assign n1334 = ~preset & ~n2578;
  assign n2580 = n1838 & ~n2512;
  assign n2581 = n_n3898 & n1887;
  assign n1339 = n2580 | n2581;
  assign n2583 = n2039 & n2536;
  assign n2584 = n_n4122 & n2029_1;
  assign n1344 = n2583 | n2584;
  assign n2586 = ~n_n3774 & ~n1672;
  assign n1349 = ~preset & ~n2586;
  assign n2588 = ~n_n3014 & ~n1672;
  assign n1354 = ~preset & ~n2588;
  assign n2590 = ~n_n4241 & ~n1672;
  assign n1359 = ~preset & ~n2590;
  assign n2592 = n_n4201 & n1664_1;
  assign n2593 = n_n3952 & n1673;
  assign n1364 = n2592 | n2593;
  assign n2595 = ~n1606 & n1664_1;
  assign n2596 = n_n3237 & n1673;
  assign n1369 = n2595 | n2596;
  assign n2598 = ~n_n3968 & ~n1890;
  assign n2599 = ~pv6_2_2_ & n1890;
  assign n2600 = ~preset & ~n2599;
  assign n1374 = ~n2598 & n2600;
  assign n2602 = ~n_n3922 & ~n1890;
  assign n2603 = ~pv6_4_4_ & n1890;
  assign n2604 = ~preset & ~n2603;
  assign n1379 = ~n2602 & n2604;
  assign n2606 = ~n_n3551 & ~n1672;
  assign n1384 = ~preset & ~n2606;
  assign n2608 = ~n_n3379 & ~n1672;
  assign n1389 = ~preset & ~n2608;
  assign n2610 = n1694_1 & n2446;
  assign n2611 = ~n_n4275 & ~n2610;
  assign n2612 = ~n_n3814 & n1694_1;
  assign n2613 = ~n1692 & ~n2612;
  assign n2614 = ~n_n3724 & n1694_1;
  assign n2615 = n2613 & ~n2614;
  assign n2616 = ~n_n4227 & n1694_1;
  assign n2617 = n2615 & ~n2616;
  assign n2618 = ~n_n3766 & n1694_1;
  assign n2619 = n_n4275 & ~n2618;
  assign n2620 = n2617 & n2619;
  assign n1394 = ~n2611 & ~n2620;
  assign n2622 = ~n_n3570 & ~n1672;
  assign n1399 = ~preset & ~n2622;
  assign n2624 = ~n_n3854 & ~n2108;
  assign n2625 = ~pv2_5_5_ & n2108;
  assign n2626 = ~preset & ~n2625;
  assign n1404 = ~n2624 & n2626;
  assign n2628 = ~n_n3845 & ~n_n3865;
  assign n2629 = ~n_n3955 & ~n_n4099;
  assign n2630 = n2628 & n2629;
  assign n2631 = ~n_n4052 & n2462;
  assign n2632 = n_n4029 & ~n2051;
  assign n2633 = ~n2052 & ~n2632;
  assign n2634 = n2631 & n2633;
  assign n2635 = n2630 & n2634;
  assign n2636 = n2057 & n2635;
  assign n2637 = n_n4056 & n2636;
  assign n2638 = n_n4057 & ~n2637;
  assign n2639 = ~preset & ~n2638;
  assign n1409 = n2060 | ~n2639;
  assign n2641 = ~n_n3451 & ~n2108;
  assign n2642 = ~pv2_7_7_ & n2108;
  assign n2643 = ~preset & ~n2642;
  assign n1414 = ~n2641 & n2643;
  assign n2645 = ~n_n4037 & ~n1672;
  assign n1419 = ~preset & ~n2645;
  assign n2647 = ~n1610 & n1664_1;
  assign n2648 = n_n3408 & n1673;
  assign n1424 = n2647 | n2648;
  assign n2650 = n_n4229 & n1887;
  assign n2651 = ~n2019_1 & ~n2020;
  assign n2652 = n2022 & ~n2651;
  assign n2653 = ~n2022 & n2651;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = n1838 & n2654;
  assign n1429 = n2650 | n2655;
  assign n2657 = ~n_n4201 & ~n1890;
  assign n2658 = ~pv6_1_1_ & n1890;
  assign n2659 = ~preset & ~n2658;
  assign n1434 = ~n2657 & n2659;
  assign n2661 = ~n_n3339 & ~n1672;
  assign n1439 = ~preset & ~n2661;
  assign n2663 = ~n1764_1 & n2414;
  assign n2664 = pv10_5_5_ & n1767;
  assign n1444 = n2663 | n2664;
  assign n2666 = n_n3483 & ~n2452;
  assign n2667 = ~n2456 & n2666;
  assign n2668 = ~n_n3483 & n2449;
  assign n2669 = n_n4334 & n2668;
  assign n1449 = n2667 | n2669;
  assign n1454 = ~preset & n2636;
  assign n2672 = ~n_n4185 & ~n1672;
  assign n1459 = ~preset & ~n2672;
  assign n2674 = n_n3934 & n1830;
  assign n2675 = n_n3069 & n1673;
  assign n1464 = n2674 | n2675;
  assign n2677 = ~n_n3643 & ~n1672;
  assign n1469 = ~preset & ~n2677;
  assign n2679 = n_n4229 & n1664_1;
  assign n2680 = n_n3404 & n1673;
  assign n1474 = n2679 | n2680;
  assign n2682 = n_n3057 & n1673;
  assign n1479 = n2469 | n2682;
  assign n2684 = ~n2249_1 & ~n2347;
  assign n2685 = n_n3020 & n1673;
  assign n1484 = ~n2684 | n2685;
  assign n2687 = ~n_n3828 & ~n1672;
  assign n1489 = ~preset & ~n2687;
  assign n2689 = n_n3631 & n1673;
  assign n1494 = n2280 | n2689;
  assign n2691 = n_n3968 & n1664_1;
  assign n2692 = n_n3138 & n1673;
  assign n1499 = n2691 | n2692;
  assign n2694 = ~ngfdn_3 & n1671;
  assign n1504 = ~n1659_1 | n2694;
  assign n2696 = n_n3922 & n1664_1;
  assign n2697 = n_n4065 & n1673;
  assign n1509 = n2696 | n2697;
  assign n2699 = n_n4366 & n1830;
  assign n2700 = n_n3679 & n1673;
  assign n1514 = n2699 | n2700;
  assign n2702 = ~n1626 & n1664_1;
  assign n2703 = n_n3287 & n1673;
  assign n1519 = n2702 | n2703;
  assign n2705 = n_n4351 & n1931;
  assign n2706 = n1933 & n2654;
  assign n1524 = n2705 | n2706;
  assign n2708 = ~n_n4059 & ~n1672;
  assign n1529 = ~preset & ~n2708;
  assign n2710 = n_n3898 & n1664_1;
  assign n2711 = n_n3436 & n1673;
  assign n1534 = n2710 | n2711;
  assign n2713 = ~nen3_10 & ~ndn3_9;
  assign n1539 = n1909_1 & ~n2713;
  assign n2715 = ~n_n3461 & ~n1672;
  assign n1544 = ~preset & ~n2715;
  assign n2717 = n2447 & n2451;
  assign n2718 = n_n4012 & n2454;
  assign n1549 = n2717 | n2718;
  assign n2720 = ~n_n3051 & ~n1672;
  assign n1554 = ~preset & ~n2720;
  assign n2722 = n_n4047 & n1830;
  assign n2723 = n_n3073 & n1673;
  assign n1559 = n2722 | n2723;
  assign n2725 = n_n3777 & n1673;
  assign n1564 = n2710 | n2725;
  assign n2727 = n_n3709 & ~n1979_1;
  assign n2728 = ~n1690 & ~n2727;
  assign n2729 = n_n3707 & ~n2728;
  assign n1569 = ~preset & n2729;
  assign n2731 = ~n1764_1 & n2387;
  assign n2732 = pv10_2_2_ & n1767;
  assign n1574 = n2731 | n2732;
  assign n2734 = n2039 & n2654;
  assign n2735 = n_n3085 & n2029_1;
  assign n1579 = n2734 | n2735;
  assign n2737 = ~pv1_7_7_ & n1915;
  assign n2738 = ~n_n3259 & ~n1915;
  assign n2739 = ~preset & ~n2738;
  assign n1584 = ~n2737 & n2739;
  assign n2741 = ~n_n3504 & ~n1672;
  assign n1589 = ~preset & ~n2741;
  assign n1594 = ~n1782 | ~n2639;
  assign n2744 = ~n_n3954 & n2068;
  assign n2745 = n_n3954 & n1778;
  assign n2746 = n_n4349 & ~n2048;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n2063 & ~n2747;
  assign n1599 = ~n2744 & ~n2748;
  assign n2750 = n_n4324 & n1830;
  assign n2751 = n_n3136 & n1673;
  assign n1604 = n2750 | n2751;
  assign n2753 = n_n4383 & n1664_1;
  assign n2754 = n_n4372 & n1673;
  assign n1609 = n2753 | n2754;
  assign n2756 = ~n1618 & n1664_1;
  assign n2757 = n_n4236 & n1673;
  assign n1614 = n2756 | n2757;
  assign n2759 = ~n_n3040 & ~n1672;
  assign n1619 = ~preset & ~n2759;
  assign n2761 = ~n_n3874 & ~n1672;
  assign n1624 = ~preset & ~n2761;
  assign n2763 = ~n_n3999 & ~n1672;
  assign n1629 = ~preset & ~n2763;
  assign n2765 = n_n3223 & n1673;
  assign n1634 = n2248 | n2765;
  assign n1639 = ndn1_34 & n1659_1;
  assign n2768 = n1703 & ~n1764_1;
  assign n2769 = pv10_1_1_ & n1767;
  assign n1644 = n2768 | n2769;
  assign n2771 = n1885 & n2039;
  assign n2772 = n_n3657 & n2029_1;
  assign n1649 = n2771 | n2772;
  assign n2774 = n_n4258 & n1664_1;
  assign n2775 = n_n3213 & n1673;
  assign n1654 = n2774 | n2775;
  assign n2777 = ~n_n3095 & ~n1672;
  assign n1659 = ~preset & ~n2777;
  assign n2779 = ~n_n3663 & ~n1672;
  assign n1664 = ~preset & ~n2779;
  assign n2781 = n_n3724 & ~n2613;
  assign n2782 = n_n3814 & n2614;
  assign n1669 = n2781 | n2782;
  assign n2784 = ~n_n3038 & ~n1672;
  assign n1674 = ~preset & ~n2784;
  assign n2786 = n_n4337 & n1664_1;
  assign n2787 = n_n3370 & n1673;
  assign n1679 = n2786 | n2787;
  assign n2789 = ~n_n3624 & ~n1676;
  assign n2790 = ~pv11_0_0_ & n1676;
  assign n2791 = ~preset & ~n2790;
  assign n1684 = ~n2789 & n2791;
  assign n2793 = ~n_n3578 & ~n1676;
  assign n2794 = ~pv11_4_4_ & n1676;
  assign n2795 = ~preset & ~n2794;
  assign n1689 = ~n2793 & n2795;
  assign n2797 = n_n3713 & n1673;
  assign n1694 = n2249_1 | n2797;
  assign n2799 = n_n3089 & n1673;
  assign n1699 = n1989_1 | n2799;
  assign n2801 = ~n_n3211 & ~n1672;
  assign n1704 = ~preset & ~n2801;
  assign n2803 = ~n_n3367 & ~n1672;
  assign n1709 = ~preset & ~n2803;
  assign n2805 = ~n_n3434 & ~n1672;
  assign n1714 = ~preset & ~n2805;
  assign n2807 = n_n3126 & n1673;
  assign n1719 = ~n2147 | n2807;
  assign n2809 = n_n4192 & n1673;
  assign n1724 = n1823 | n2809;
  assign n2811 = n_n3876 & n1664_1;
  assign n2812 = n_n4136 & n1673;
  assign n1729 = n2811 | n2812;
  assign n2814 = ~n_n3053 & ~n1672;
  assign n1734 = ~preset & ~n2814;
  assign n2816 = ~n_n3938 & ~n1672;
  assign n1739 = ~preset & ~n2816;
  assign n2818 = n_n3769 & n1785;
  assign n2819 = n_n4229 & n1798;
  assign n2820 = n1800 & ~n2819;
  assign n2821 = ~n_n4229 & n1797;
  assign n2822 = n1787 & ~n2821;
  assign n2823 = ~n2820 & n2822;
  assign n1744 = n2818 | n2823;
  assign n2825 = n_n4390 & n1673;
  assign n1749 = n2130 | n2825;
  assign n2827 = nen3_10 & ~n2115;
  assign n2828 = nsr3_17 & ~n2827;
  assign n1754 = ~n1659_1 | n2828;
  assign n2830 = ~n_n3903 & ~n1672;
  assign n1759 = ~preset & ~n2830;
  assign n2832 = ~n_n3658 & ~n1755;
  assign n1764 = n2078 & ~n2832;
  assign n2834 = ~nrq3_11 & nsr3_14;
  assign n1769 = n1909_1 & ~n2834;
  assign n2836 = n_n3818 & n1692;
  assign n2837 = n1690 & n1765;
  assign n2838 = n1694_1 & ~n1965;
  assign n2839 = ~n2837 & ~n2838;
  assign n1774 = n2836 | ~n2839;
  assign n2841 = ~n_n3533 & ~n1890;
  assign n2842 = ~pv6_3_3_ & n1890;
  assign n2843 = ~preset & ~n2842;
  assign n1779 = ~n2841 & n2843;
  assign n2845 = n_n4316 & n1664_1;
  assign n2846 = n_n3463 & n1673;
  assign n1784 = n2845 | n2846;
  assign n2848 = ~n_n3175 & ~n1672;
  assign n1789 = ~preset & ~n2848;
  assign n2850 = n_n3055 & n1673;
  assign n1794 = n2190 | n2850;
  assign n2852 = n_n3202 & n1673;
  assign n1799 = ~n2193 | n2852;
  assign n2854 = n_n3385 & n1673;
  assign n1804 = ~n2684 | n2854;
  assign n2856 = ~n_n4077 & ~n1672;
  assign n1809 = ~preset & ~n2856;
  assign n2858 = ~n_n3142 & ~n1672;
  assign n1814 = ~preset & ~n2858;
  assign n2860 = ~n1793 & ~n1794_1;
  assign n2861 = n_n4316 & ~n2860;
  assign n2862 = ~n1793 & n1795;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = n1787 & ~n2863;
  assign n2865 = n_n3901 & n1785;
  assign n1819 = n2864 | n2865;
  assign n2867 = n_n3976 & n1787;
  assign n2868 = ~n_n3934 & ~n2867;
  assign n2869 = n1787 & ~n1790;
  assign n2870 = ~n1785 & ~n2869;
  assign n1824 = ~n2868 & ~n2870;
  assign n2872 = n_n4227 & n1669_1;
  assign n2873 = n_n3823 & n1673;
  assign n1829 = n2872 | n2873;
  assign n2875 = n_n4160 & n1664_1;
  assign n2876 = n_n3722 & n1673;
  assign n1834 = n2875 | n2876;
  assign n2878 = n_n4182 & n1664_1;
  assign n2879 = n_n4309 & n1673;
  assign n1839 = n2878 | n2879;
  assign n2881 = ~n_n4159 & ~n1940;
  assign n2882 = ~pv4_0_0_ & n1940;
  assign n2883 = ~preset & ~n2882;
  assign n1844 = ~n2881 & n2883;
  assign n2885 = ~n_n4330 & ~n1940;
  assign n2886 = ~pv4_4_4_ & n1940;
  assign n2887 = ~preset & ~n2886;
  assign n1849 = ~n2885 & n2887;
  assign n2889 = ~n_n3836 & ~n1672;
  assign n1854 = ~preset & ~n2889;
  assign n2891 = ~n_n3470 & ~n1672;
  assign n1859 = ~preset & ~n2891;
  assign n2893 = n_n3331 & n1673;
  assign n1864 = n1707 | n2893;
  assign n2895 = n_n3883 & n1673;
  assign n1869 = n2129_1 | n2895;
  assign n2897 = ~preset & n_n4299;
  assign n2898 = ~n1764_1 & n2897;
  assign n2899 = pv10_6_6_ & n1767;
  assign n1874 = n2898 | n2899;
  assign n2901 = n2039 & ~n2512;
  assign n2902 = n_n4157 & n2029_1;
  assign n1879 = n2901 | n2902;
  assign n2904 = ~ndn3_8 & ~ndn3_9;
  assign n1884 = n1909_1 & ~n2904;
  assign n2906 = ~pv1_1_1_ & n1915;
  assign n2907 = ~n_n3208 & ~n1915;
  assign n2908 = ~preset & ~n2907;
  assign n1889 = ~n2906 & n2908;
  assign n2910 = ~n_n3190 & ~n1672;
  assign n1894 = ~preset & ~n2910;
  assign n2912 = n_n4029 & n2068;
  assign n2913 = n_n3533 & ~n2048;
  assign n2914 = n1778 & ~n2633;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n2063 & ~n2915;
  assign n1899 = n2912 | n2916;
  assign n2918 = ~n_n3042 & ~n1672;
  assign n1904 = ~preset & ~n2918;
  assign n2920 = ~nsr3_17 & ~n1781;
  assign n2921 = nsr3_14 & ~n2920;
  assign n1909 = ~n1659_1 | n2921;
  assign n2923 = ~nlc1_2 & n2284;
  assign n2924 = ~preset & ~n2923;
  assign n1914 = n_n4151 | ~n2924;
  assign n2926 = ~n_n3188 & ~n1672;
  assign n1919 = ~preset & ~n2926;
  assign n2928 = n_n3769 & n1830;
  assign n2929 = n_n4303 & n1673;
  assign n1924 = n2928 | n2929;
  assign n2931 = ~n_n3250 & ~n1676;
  assign n2932 = ~pv11_3_3_ & n1676;
  assign n2933 = ~preset & ~n2932;
  assign n1929 = ~n2931 & n2933;
  assign n2935 = ~n_n3170 & ~n1676;
  assign n2936 = ~pv11_7_7_ & n1676;
  assign n2937 = ~preset & ~n2936;
  assign n1934 = ~n2935 & n2937;
  assign n2939 = n_n3758 & n1673;
  assign n1939 = n2091 | n2939;
  assign n2941 = n_n3910 & n1673;
  assign n1944 = ~n2542 | n2941;
  assign n2943 = ~n2130 & ~n2257;
  assign n2944 = n_n3108 & n1673;
  assign n1949 = ~n2943 | n2944;
  assign n2946 = ~n_n3150 & ~n1672;
  assign n1954 = ~preset & ~n2946;
  assign n2948 = n_n4320 & n1673;
  assign n1959 = n1822 | n2948;
  assign n2950 = n1741 & ~n1764_1;
  assign n2951 = pv10_7_7_ & n1767;
  assign n1964 = n2950 | n2951;
  assign n2953 = n_n4362 & n1664_1;
  assign n2954 = n_n4247 & n1673;
  assign n1969 = n2953 | n2954;
  assign n2956 = n_n4199 & n1673;
  assign n1974 = n2105 | n2956;
  assign n2958 = n_n4275 & n1669_1;
  assign n2959 = n_n3966 & n1673;
  assign n1979 = n2958 | n2959;
  assign n2961 = n_n3766 & ~n2617;
  assign n2962 = n2445 & n2618;
  assign n1984 = n2961 | n2962;
  assign n2964 = ~n_n4021 & ~n2108;
  assign n2965 = ~pv2_4_4_ & n2108;
  assign n2966 = ~preset & ~n2965;
  assign n1989 = ~n2964 & n2966;
  assign n2968 = ~n_n4062 & ~n2108;
  assign n2969 = ~pv2_6_6_ & n2108;
  assign n2970 = ~preset & ~n2969;
  assign n1994 = ~n2968 & n2970;
  assign n2972 = n_n3814 & n1669_1;
  assign n2973 = n_n3514 & n1673;
  assign n1999 = n2972 | n2973;
  assign n2975 = ~n1620 & n1664_1;
  assign n2976 = n_n3572 & n1673;
  assign n2004 = n2975 | n2976;
  assign n2978 = n_n4270 & n1664_1;
  assign n2979 = n_n4166 & n1673;
  assign n2009 = n2978 | n2979;
  assign n2981 = n1838 & n2142;
  assign n2982 = n_n3976 & n1887;
  assign n2014 = n2981 | n2982;
  assign n2984 = n_n3841 & n1664_1;
  assign n2985 = n_n3394 & n1673;
  assign n2019 = n2984 | n2985;
  assign n2987 = n1933 & n2536;
  assign n2988 = n_n4095 & n1931;
  assign n2024 = n2987 | n2988;
  assign n2990 = ~n_n3863 & ~n1672;
  assign n2029 = ~preset & ~n2990;
  assign n2992 = ~n_n3720 & ~n1672;
  assign n2034 = ~preset & ~n2992;
  assign n2994 = ~preset & n_n3756;
  assign n2995 = ~n1764_1 & n2994;
  assign n2996 = pv10_0_0_ & n1767;
  assign n2044 = n2995 | n2996;
  assign n2998 = n_n3667 & n1673;
  assign n2049 = ~n1990 | n2998;
  assign n3000 = n_n4299 & n1664_1;
  assign n3001 = n_n3342 & n1673;
  assign n2054 = n3000 | n3001;
  assign n3003 = ~n_n3529 & ~n1672;
  assign n2059 = ~preset & ~n3003;
  assign n3005 = n_n3756 & n1664_1;
  assign n3006 = n_n4209 & n1673;
  assign n2064 = n3005 | n3006;
  assign n3008 = ~n_n3475 & ~n1810;
  assign n3009 = ~n1809_1 & ~n3008;
  assign n3010 = ~n_n3841 & n3009;
  assign n3011 = n_n3841 & ~n3009;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = n1787 & ~n3012;
  assign n3014 = ~n_n4324 & ~n3013;
  assign n3015 = n1787 & n3012;
  assign n3016 = n_n4324 & ~n1785;
  assign n3017 = ~n3015 & n3016;
  assign n2069 = ~n3014 & ~n3017;
  assign n3019 = n_n3337 & n1673;
  assign n2074 = n1708 | n3019;
  assign n3021 = n_n4227 & ~n2615;
  assign n3022 = n2444 & n2616;
  assign n2079 = n3021 | n3022;
  assign n3024 = ~n_n4153 & ~n1672;
  assign n2084 = ~preset & ~n3024;
  assign n3026 = ~n1667 & n2113;
  assign n3027 = n2185 & ~n3026;
  assign n3028 = n_n3831 & ~n3027;
  assign n2089 = ~n2117 | n3028;
  assign n3030 = ~n_n3233 & ~n1672;
  assign n2094 = ~preset & ~n3030;
  assign n3032 = ~nlc3_3 & n2291;
  assign n3033 = ~n_n4263 & ~n3032;
  assign n2099 = ~preset & ~n3033;
  assign n3035 = n_n4251 & n1664_1;
  assign n3036 = n_n3413 & n1673;
  assign n2104 = n3035 | n3036;
  assign n3038 = ~n_n4182 & ~n1940;
  assign n3039 = ~pv4_3_3_ & n1940;
  assign n3040 = ~preset & ~n3039;
  assign n2109 = ~n3038 & n3040;
  assign n3042 = n1838 & n2244_1;
  assign n3043 = n_n3841 & n1887;
  assign n2114 = n3042 | n3043;
  assign n3045 = ~n_n3441 & ~n1672;
  assign n2119 = ~preset & ~n3045;
  assign n3047 = ~n_n4026 & ~n1687;
  assign n2124 = n2117 & ~n3047;
  assign n3049 = n_n4342 & n1673;
  assign n2129 = n2679 | n3049;
  assign n3051 = n_n4102 & n1673;
  assign n2134 = n2984 | n3051;
  assign n3053 = n_n3277 & n1673;
  assign n2139 = ~n1902 | n3053;
  assign n3055 = n_n4180 & n1673;
  assign n2144 = n2280 | n3055;
  assign n3057 = ~pv1_0_0_ & n1915;
  assign n3058 = ~n_n3878 & ~n1915;
  assign n3059 = ~preset & ~n3058;
  assign n2149 = ~n3057 & n3059;
  assign n3061 = ~n_n3931 & ~n2108;
  assign n3062 = ~pv2_0_0_ & n2108;
  assign n3063 = ~preset & ~n3062;
  assign n2154 = ~n3061 & n3063;
  assign n3065 = n_n3845 & n2068;
  assign n3066 = n_n3968 & ~n2048;
  assign n3067 = n_n3845 & ~n2050;
  assign n3068 = ~n2051 & ~n3067;
  assign n3069 = n1778 & ~n3068;
  assign n3070 = ~n3066 & ~n3069;
  assign n3071 = n2063 & ~n3070;
  assign n2159 = n3065 | n3071;
  assign n3073 = n_n3865 & n2068;
  assign n3074 = n_n3922 & ~n2048;
  assign n3075 = n_n3865 & ~n2052;
  assign n3076 = ~n2053 & ~n3075;
  assign n3077 = n1778 & ~n3076;
  assign n3078 = ~n3074 & ~n3077;
  assign n3079 = n2063 & ~n3078;
  assign n2164 = n3073 | n3079;
  assign n3081 = n_n3533 & n1664_1;
  assign n3082 = n_n3486 & n1673;
  assign n2169 = n3081 | n3082;
  assign n3084 = ~n_n4056 & ~n1782;
  assign n3085 = ~preset & ~n3084;
  assign n2174 = n2638 & n3085;
  assign n3087 = ~n_n3674 & ~n1672;
  assign n2179 = ~preset & ~n3087;
  assign n3089 = ~n1620 & n1682;
  assign n3090 = n_n3959 & ~n2452;
  assign n3091 = ~n3089 & n3090;
  assign n3092 = n1690 & n2994;
  assign n3093 = n1694_1 & n1695;
  assign n3094 = ~n3092 & ~n3093;
  assign n2184 = n3091 | ~n3094;
  assign n3096 = n_n3608 & n1931;
  assign n3097 = n1933 & n2142;
  assign n2189 = n3096 | n3097;
  assign n3099 = n_n4080 & n1692;
  assign n3100 = n1690 & n2897;
  assign n3101 = ~n1606 & n1945;
  assign n3102 = ~n1946 & ~n3101;
  assign n3103 = n1694_1 & ~n3102;
  assign n3104 = ~n3100 & ~n3103;
  assign n2194 = n3099 | ~n3104;
  assign n3106 = ~n_n4018 & ~n1672;
  assign n2199 = ~preset & ~n3106;
  assign n3108 = ~n_n4354 & ~n1672;
  assign n2204 = ~preset & ~n3108;
  assign n3110 = ~n_n3797 & ~n1672;
  assign n2209 = ~preset & ~n3110;
  assign n3112 = n_n3739 & n1673;
  assign n2214 = n2845 | n3112;
  assign n3114 = n_n3646 & n1673;
  assign n2219 = ~n2943 | n3114;
  assign n3116 = ~n1937 & n2039;
  assign n3117 = n_n3099 & n2029_1;
  assign n2224 = n3116 | n3117;
  assign n3119 = n_n3537 & n1673;
  assign n2229 = n2191 | n3119;
  assign n3121 = n_n3806 & n1673;
  assign n2234 = n1989_1 | n3121;
  assign n3123 = ~n_n3087 & ~n1672;
  assign n2239 = ~preset & ~n3123;
  assign n3125 = ~n_n4105 & ~n1672;
  assign n2244 = ~preset & ~n3125;
  assign n3127 = ~n_n3262 & ~n1672;
  assign n2249 = ~preset & ~n3127;
  assign n3129 = n_n4125 & n1785;
  assign n3130 = ~n1788 & ~n1789_1;
  assign n3131 = n1790 & n3130;
  assign n3132 = ~n1790 & ~n3130;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n1787 & n3133;
  assign n2254 = n3129 | n3134;
  assign n3136 = n_n3814 & n1692;
  assign n2259 = n2612 | n3136;
  assign n3138 = n_n3831 & ~n1656;
  assign n3139 = n3026 & n3138;
  assign n2264 = ~n2186 | n3139;
  assign n3141 = nsr4_2 & n1905;
  assign n3142 = n1659_1 & ~n3141;
  assign n2269 = n1906 | ~n3142;
  assign n1259 = 1'b0;
  always @ (posedge clock) begin
    n_n4142 <= n350;
    n_n3936 <= n355;
    n_n3574 <= n360;
    n_n3008 <= n365;
    n_n3726 <= n370;
    n_n3604 <= n375;
    n_n3144 <= n380;
    n_n3782 <= n385;
    n_n3067 <= n390;
    n_n4258 <= n395;
    n_n3225 <= n400;
    n_n3180 <= n405;
    n_n3274 <= n410;
    n_n3475 <= n415;
    n_n3687 <= n420;
    n_n3381 <= n425;
    n_n3098 <= n430;
    n_n4108 <= n435;
    n_n3497 <= n440;
    n_n3793 <= n445;
    n_n4316 <= n450;
    n_n4349 <= n455;
    n_n3029 <= n460;
    n_n3619 <= n465;
    n_n3264 <= n470;
    n_n3780 <= n475;
    ndn3_4 <= n480;
    n_n4114 <= n485;
    n_n3146 <= n490;
    n_n3511 <= n495;
    n_n3152 <= n500;
    n_n3833 <= n505;
    n_n4282 <= n510;
    n_n3305 <= n515;
    n_n4392 <= n520;
    n_n4224 <= n525;
    n_n3198 <= n530;
    n_n3204 <= n535;
    n_n3024 <= n540;
    n_n4139 <= n545;
    ndn3_15 <= n550;
    n_n3133 <= n555;
    n_n4074 <= n560;
    n_n3270 <= n565;
    n_n3858 <= n570;
    n_n3456 <= n575;
    n_n3521 <= n580;
    n_n3081 <= n585;
    n_n4381 <= n590;
    n_n3670 <= n595;
    n_n4211 <= n600;
    n_n3493 <= n605;
    n_n3495 <= n610;
    n_n3916 <= n615;
    n_n3195 <= n620;
    n_n3525 <= n625;
    n_n3729 <= n630;
    n_n3876 <= n635;
    ndn3_5 <= n640;
    n_n3549 <= n645;
    n_n3489 <= n650;
    n_n3764 <= n655;
    n_n3281 <= n660;
    n_n3707 <= n665;
    n_n3517 <= n670;
    n_n4160 <= n675;
    n_n4222 <= n680;
    n_n3012 <= n685;
    n_n4071 <= n690;
    n_n3372 <= n695;
    n_n3344 <= n700;
    n_n3688 <= n705;
    n_n3079 <= n710;
    n_n3313 <= n715;
    n_n3411 <= n720;
    n_n3231 <= n725;
    n_n3396 <= n730;
    n_n3432 <= n735;
    n_n3606 <= n740;
    n_n3733 <= n745;
    n_n3556 <= n750;
    n_n4040 <= n755;
    n_n3120 <= n760;
    n_n3221 <= n765;
    n_n3173 <= n770;
    n_n3851 <= n775;
    n_n3113 <= n780;
    n_n3242 <= n785;
    n_n3118 <= n790;
    n_n3376 <= n795;
    n_n4089 <= n800;
    n_n3044 <= n805;
    n_n3627 <= n810;
    n_n3035 <= n815;
    n_n3111 <= n820;
    n_n3321 <= n825;
    n_n3443 <= n830;
    n_n3215 <= n835;
    ndn3_10 <= n840;
    n_n4172 <= n845;
    nlc1_2 <= n850;
    n_n3590 <= n855;
    n_n4110 <= n860;
    nlc3_3 <= n865;
    n_n3576 <= n870;
    n_n4129 <= n875;
    n_n4189 <= n880;
    n_n4286 <= n885;
    n_n4383 <= n890;
    pdn <= n895;
    n_n3567 <= n899;
    n_n3892 <= n904;
    n_n3075 <= n909;
    n_n3354 <= n914;
    n_n3465 <= n919;
    ndn3_6 <= n924;
    n_n3617 <= n929;
    n_n4162 <= n934;
    n_n3207 <= n939;
    n_n4120 <= n944;
    n_n3065 <= n949;
    n_n4005 <= n954;
    n_n3266 <= n959;
    n_n4337 <= n964;
    n_n3600 <= n969;
    n_n3415 <= n974;
    n_n4243 <= n979;
    n_n3872 <= n984;
    n_n3648 <= n989;
    n_n3358 <= n994;
    n_n3350 <= n999;
    ndn3_7 <= n1004;
    n_n3116 <= n1009;
    n_n3583 <= n1014;
    n_n3906 <= n1019;
    n_n4131 <= n1024;
    n_n3316 <= n1029;
    n_n3061 <= n1034;
    n_n3048 <= n1039;
    n_n3886 <= n1044;
    n_n3919 <= n1049;
    n_n3128 <= n1054;
    n_n3995 <= n1059;
    n_n4213 <= n1064;
    n_n3761 <= n1069;
    ndn3_8 <= n1074;
    n_n3252 <= n1079;
    n_n4366 <= n1084;
    n_n3328 <= n1089;
    n_n3988 <= n1094;
    n_n3348 <= n1099;
    n_n3544 <= n1104;
    n_n3101 <= n1109;
    n_n4279 <= n1114;
    n_n3896 <= n1119;
    n_n3736 <= n1124;
    n_n4251 <= n1129;
    n_n3650 <= n1134;
    n_n3307 <= n1139;
    n_n4294 <= n1144;
    n_n4334 <= n1149;
    n_n3955 <= n1154;
    n_n4164 <= n1159;
    n_n3155 <= n1164;
    n_n3749 <= n1169;
    n_n4233 <= n1174;
    n_n4347 <= n1179;
    n_n3826 <= n1184;
    n_n3360 <= n1189;
    n_n3458 <= n1194;
    n_n3093 <= n1199;
    n_n3157 <= n1204;
    n_n3506 <= n1209;
    n_n3161 <= n1214;
    n_n3319 <= n1219;
    n_n3429 <= n1224;
    n_n3971 <= n1229;
    n_n3449 <= n1234;
    n_n4270 <= n1239;
    n_n4288 <= n1244;
    n_n3183 <= n1249;
    n_n3130 <= n1254;
    nlak4_2 <= n1259;
    n_n4047 <= n1264;
    n_n3978 <= n1269;
    n_n3239 <= n1274;
    n_n4145 <= n1279;
    n_n3890 <= n1284;
    n_n4003 <= n1289;
    n_n3091 <= n1294;
    n_n3985 <= n1299;
    n_n3326 <= n1304;
    n_n4052 <= n1309;
    nsr4_2 <= n1314;
    n_n4099 <= n1319;
    n_n4375 <= n1324;
    n_n4067 <= n1329;
    n_n4290 <= n1334;
    n_n3898 <= n1339;
    n_n4122 <= n1344;
    n_n3774 <= n1349;
    n_n3014 <= n1354;
    n_n4241 <= n1359;
    n_n3952 <= n1364;
    n_n3237 <= n1369;
    n_n3968 <= n1374;
    n_n3922 <= n1379;
    n_n3551 <= n1384;
    n_n3379 <= n1389;
    n_n4275 <= n1394;
    n_n3570 <= n1399;
    n_n3854 <= n1404;
    n_n4057 <= n1409;
    n_n3451 <= n1414;
    n_n4037 <= n1419;
    n_n3408 <= n1424;
    n_n4229 <= n1429;
    n_n4201 <= n1434;
    n_n3339 <= n1439;
    n_n4362 <= n1444;
    n_n3483 <= n1449;
    n_n3557 <= n1454;
    n_n4185 <= n1459;
    n_n3069 <= n1464;
    n_n3643 <= n1469;
    n_n3404 <= n1474;
    n_n3057 <= n1479;
    n_n3020 <= n1484;
    n_n3828 <= n1489;
    n_n3631 <= n1494;
    n_n3138 <= n1499;
    nsr1_2 <= n1504;
    n_n4065 <= n1509;
    n_n3679 <= n1514;
    n_n3287 <= n1519;
    n_n4351 <= n1524;
    n_n4059 <= n1529;
    n_n3436 <= n1534;
    nen3_10 <= n1539;
    n_n3461 <= n1544;
    n_n4012 <= n1549;
    n_n3051 <= n1554;
    n_n3073 <= n1559;
    n_n3777 <= n1564;
    n_n3709 <= n1569;
    n_n3946 <= n1574;
    n_n3085 <= n1579;
    n_n3259 <= n1584;
    n_n3504 <= n1589;
    n_n4045 <= n1594;
    n_n3954 <= n1599;
    n_n3136 <= n1604;
    n_n4372 <= n1609;
    n_n4236 <= n1614;
    n_n3040 <= n1619;
    n_n3874 <= n1624;
    n_n3999 <= n1629;
    n_n3223 <= n1634;
    ndn1_34 <= n1639;
    n_n3743 <= n1644;
    n_n3657 <= n1649;
    n_n3213 <= n1654;
    n_n3095 <= n1659;
    n_n3663 <= n1664;
    n_n3724 <= n1669;
    n_n3038 <= n1674;
    n_n3370 <= n1679;
    n_n3624 <= n1684;
    n_n3578 <= n1689;
    n_n3713 <= n1694;
    n_n3089 <= n1699;
    n_n3211 <= n1704;
    n_n3367 <= n1709;
    n_n3434 <= n1714;
    n_n3126 <= n1719;
    n_n4192 <= n1724;
    n_n4136 <= n1729;
    n_n3053 <= n1734;
    n_n3938 <= n1739;
    n_n3769 <= n1744;
    n_n4390 <= n1749;
    nsr3_17 <= n1754;
    n_n3903 <= n1759;
    n_n3658 <= n1764;
    nrq3_11 <= n1769;
    n_n3818 <= n1774;
    n_n3533 <= n1779;
    n_n3463 <= n1784;
    n_n3175 <= n1789;
    n_n3055 <= n1794;
    n_n3202 <= n1799;
    n_n3385 <= n1804;
    n_n4077 <= n1809;
    n_n3142 <= n1814;
    n_n3901 <= n1819;
    n_n3934 <= n1824;
    n_n3823 <= n1829;
    n_n3722 <= n1834;
    n_n4309 <= n1839;
    n_n4159 <= n1844;
    n_n4330 <= n1849;
    n_n3836 <= n1854;
    n_n3470 <= n1859;
    n_n3331 <= n1864;
    n_n3883 <= n1869;
    n_n4299 <= n1874;
    n_n4157 <= n1879;
    ndn3_9 <= n1884;
    n_n3208 <= n1889;
    n_n3190 <= n1894;
    n_n4029 <= n1899;
    n_n3042 <= n1904;
    nsr3_14 <= n1909;
    n_n4151 <= n1914;
    n_n3188 <= n1919;
    n_n4303 <= n1924;
    n_n3250 <= n1929;
    n_n3170 <= n1934;
    n_n3758 <= n1939;
    n_n3910 <= n1944;
    n_n3108 <= n1949;
    n_n3150 <= n1954;
    n_n4320 <= n1959;
    n_n4360 <= n1964;
    n_n4247 <= n1969;
    n_n4199 <= n1974;
    n_n3966 <= n1979;
    n_n3766 <= n1984;
    n_n4021 <= n1989;
    n_n4062 <= n1994;
    n_n3514 <= n1999;
    n_n3572 <= n2004;
    n_n4166 <= n2009;
    n_n3976 <= n2014;
    n_n3394 <= n2019;
    n_n4095 <= n2024;
    n_n3863 <= n2029;
    n_n3720 <= n2034;
    ngfdn_3 <= n2039;
    n_n3756 <= n2044;
    n_n3667 <= n2049;
    n_n3342 <= n2054;
    n_n3529 <= n2059;
    n_n4209 <= n2064;
    n_n4324 <= n2069;
    n_n3337 <= n2074;
    n_n4227 <= n2079;
    n_n4153 <= n2084;
    n_n3831 <= n2089;
    n_n3233 <= n2094;
    n_n4263 <= n2099;
    n_n3413 <= n2104;
    n_n4182 <= n2109;
    n_n3841 <= n2114;
    n_n3441 <= n2119;
    n_n4026 <= n2124;
    n_n4342 <= n2129;
    n_n4102 <= n2134;
    n_n3277 <= n2139;
    n_n4180 <= n2144;
    n_n3878 <= n2149;
    n_n3931 <= n2154;
    n_n3845 <= n2159;
    n_n3865 <= n2164;
    n_n3486 <= n2169;
    n_n4056 <= n2174;
    n_n3674 <= n2179;
    n_n3959 <= n2184;
    n_n3608 <= n2189;
    n_n4080 <= n2194;
    n_n4018 <= n2199;
    n_n4354 <= n2204;
    n_n3797 <= n2209;
    n_n3739 <= n2214;
    n_n3646 <= n2219;
    n_n3099 <= n2224;
    n_n3537 <= n2229;
    n_n3806 <= n2234;
    n_n3087 <= n2239;
    n_n4105 <= n2244;
    n_n3262 <= n2249;
    n_n4125 <= n2254;
    n_n3814 <= n2259;
    n_n4093 <= n2264;
    nsr3_3 <= n2269;
  end
endmodule


