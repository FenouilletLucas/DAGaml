// Benchmark "i6" written by ABC on Tue May 16 16:07:50 2017

module i6 ( 
    \V32(30) , \V138(3) , \V138(2) , \V138(4) , \V138(0) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(4) , \V32(5) , \V131(27) , \V32(6) ,
    \V131(26) , \V32(7) , \V131(29) , \V32(8) , \V131(28) , \V32(9) ,
    \V96(0) , \V96(1) , \V131(21) , \V96(2) , \V131(20) , \V96(3) ,
    \V131(23) , \V96(4) , \V96(13) , \V131(22) , \V96(5) , \V96(12) ,
    \V131(25) , \V96(6) , \V97(0) , \V96(15) , \V131(24) , \V96(7) ,
    \V96(14) , \V131(17) , \V96(8) , \V131(16) , \V96(9) , \V131(19) ,
    \V96(11) , \V131(18) , \V96(10) , \V98(0) , \V96(17) , \V96(16) ,
    \V131(11) , \V96(19) , \V131(10) , \V99(0) , \V96(18) , \V131(13) ,
    \V96(23) , \V131(12) , \V96(22) , \V131(15) , \V64(13) , \V96(25) ,
    \V131(14) , \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V96(21) ,
    \V96(20) , \V64(11) , \V64(10) , \V96(27) , \V96(26) , \V64(17) ,
    \V96(29) , \V64(16) , \V96(28) , \V131(3) , \V64(19) , \V131(2) ,
    \V64(18) , \V131(5) , \V64(23) , \V131(4) , \V64(22) , \V32(13) ,
    \V64(25) , \V32(12) , \V64(24) , \V32(15) , \V131(1) , \V32(14) ,
    \V96(31) , \V131(0) , \V96(30) , \V64(21) , \V64(20) , \V32(11) ,
    \V32(10) , \V131(7) , \V131(6) , \V131(9) , \V131(31) , \V64(27) ,
    \V131(8) , \V131(30) , \V64(26) , \V32(17) , \V64(29) , \V32(16) ,
    \V64(28) , \V32(19) , \V32(18) , \V133(1) , \V32(23) , \V133(0) ,
    \V64(0) , \V32(22) , \V64(1) , \V32(25) , \V64(2) , \V32(24) ,
    \V64(3) , \V64(4) , \V64(31) , \V64(5) , \V64(30) , \V32(21) ,
    \V64(6) , \V134(0) , \V32(20) , \V64(7) , \V64(8) , \V64(9) ,
    \V32(27) , \V32(26) , \V32(29) , \V32(28) , \V32(31) ,
    \V198(7) , \V198(6) , \V198(9) , \V198(8) , \V166(3) , \V166(2) ,
    \V166(5) , \V166(4) , \V166(1) , \V166(0) , \V166(7) , \V166(6) ,
    \V166(9) , \V198(27) , \V166(8) , \V205(3) , \V198(26) , \V205(2) ,
    \V198(29) , \V205(5) , \V198(28) , \V205(4) , \V205(1) , \V205(0) ,
    \V198(21) , \V198(20) , \V198(23) , \V198(22) , \V205(6) , \V198(25) ,
    \V198(24) , \V198(17) , \V198(16) , \V166(27) , \V198(19) , \V166(26) ,
    \V198(18) , \V198(11) , \V198(10) , \V166(21) , \V198(13) , \V166(20) ,
    \V198(12) , \V166(23) , \V198(15) , \V166(22) , \V198(14) , \V166(25) ,
    \V166(24) , \V166(17) , \V166(16) , \V166(19) , \V166(18) , \V166(11) ,
    \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) , \V198(3) ,
    \V198(2) , \V198(5) , \V198(4) , \V198(31) , \V198(30) , \V198(1) ,
    \V198(0)   );
  input  \V32(30) , \V138(3) , \V138(2) , \V138(4) , \V138(0) , \V32(0) ,
    \V32(1) , \V32(2) , \V32(3) , \V32(4) , \V32(5) , \V131(27) , \V32(6) ,
    \V131(26) , \V32(7) , \V131(29) , \V32(8) , \V131(28) , \V32(9) ,
    \V96(0) , \V96(1) , \V131(21) , \V96(2) , \V131(20) , \V96(3) ,
    \V131(23) , \V96(4) , \V96(13) , \V131(22) , \V96(5) , \V96(12) ,
    \V131(25) , \V96(6) , \V97(0) , \V96(15) , \V131(24) , \V96(7) ,
    \V96(14) , \V131(17) , \V96(8) , \V131(16) , \V96(9) , \V131(19) ,
    \V96(11) , \V131(18) , \V96(10) , \V98(0) , \V96(17) , \V96(16) ,
    \V131(11) , \V96(19) , \V131(10) , \V99(0) , \V96(18) , \V131(13) ,
    \V96(23) , \V131(12) , \V96(22) , \V131(15) , \V64(13) , \V96(25) ,
    \V131(14) , \V64(12) , \V96(24) , \V64(15) , \V64(14) , \V96(21) ,
    \V96(20) , \V64(11) , \V64(10) , \V96(27) , \V96(26) , \V64(17) ,
    \V96(29) , \V64(16) , \V96(28) , \V131(3) , \V64(19) , \V131(2) ,
    \V64(18) , \V131(5) , \V64(23) , \V131(4) , \V64(22) , \V32(13) ,
    \V64(25) , \V32(12) , \V64(24) , \V32(15) , \V131(1) , \V32(14) ,
    \V96(31) , \V131(0) , \V96(30) , \V64(21) , \V64(20) , \V32(11) ,
    \V32(10) , \V131(7) , \V131(6) , \V131(9) , \V131(31) , \V64(27) ,
    \V131(8) , \V131(30) , \V64(26) , \V32(17) , \V64(29) , \V32(16) ,
    \V64(28) , \V32(19) , \V32(18) , \V133(1) , \V32(23) , \V133(0) ,
    \V64(0) , \V32(22) , \V64(1) , \V32(25) , \V64(2) , \V32(24) ,
    \V64(3) , \V64(4) , \V64(31) , \V64(5) , \V64(30) , \V32(21) ,
    \V64(6) , \V134(0) , \V32(20) , \V64(7) , \V64(8) , \V64(9) ,
    \V32(27) , \V32(26) , \V32(29) , \V32(28) , \V32(31) ;
  output \V198(7) , \V198(6) , \V198(9) , \V198(8) , \V166(3) , \V166(2) ,
    \V166(5) , \V166(4) , \V166(1) , \V166(0) , \V166(7) , \V166(6) ,
    \V166(9) , \V198(27) , \V166(8) , \V205(3) , \V198(26) , \V205(2) ,
    \V198(29) , \V205(5) , \V198(28) , \V205(4) , \V205(1) , \V205(0) ,
    \V198(21) , \V198(20) , \V198(23) , \V198(22) , \V205(6) , \V198(25) ,
    \V198(24) , \V198(17) , \V198(16) , \V166(27) , \V198(19) , \V166(26) ,
    \V198(18) , \V198(11) , \V198(10) , \V166(21) , \V198(13) , \V166(20) ,
    \V198(12) , \V166(23) , \V198(15) , \V166(22) , \V198(14) , \V166(25) ,
    \V166(24) , \V166(17) , \V166(16) , \V166(19) , \V166(18) , \V166(11) ,
    \V166(10) , \V166(13) , \V166(12) , \V166(15) , \V166(14) , \V198(3) ,
    \V198(2) , \V198(5) , \V198(4) , \V198(31) , \V198(30) , \V198(1) ,
    \V198(0) ;
  wire n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n218, n219, n220, n221, n222, n224, n225, n226, n227, n228, n230, n231,
    n232, n233, n234, n236, n237, n238, n239, n241, n242, n243, n244, n246,
    n247, n248, n249, n251, n252, n253, n254, n256, n257, n258, n259, n261,
    n262, n263, n264, n266, n267, n268, n269, n271, n272, n273, n274, n276,
    n277, n278, n279, n281, n282, n283, n284, n285, n287, n288, n289, n290,
    n292, n293, n294, n295, n296, n297, n298, n299, n301, n302, n303, n304,
    n305, n307, n308, n309, n310, n311, n313, n314, n315, n316, n317, n319,
    n320, n321, n322, n323, n325, n326, n327, n328, n329, n331, n332, n333,
    n334, n335, n337, n338, n339, n340, n341, n343, n344, n345, n346, n347,
    n349, n350, n351, n352, n353, n355, n356, n357, n358, n359, n361, n362,
    n363, n364, n365, n367, n368, n369, n370, n371, n373, n374, n375, n377,
    n378, n379, n380, n381, n383, n384, n385, n386, n387, n389, n390, n391,
    n392, n393, n395, n396, n397, n398, n399, n401, n402, n403, n404, n406,
    n407, n408, n409, n410, n412, n413, n414, n415, n417, n418, n419, n420,
    n421, n423, n424, n425, n426, n427, n429, n430, n431, n432, n433, n435,
    n436, n437, n438, n440, n441, n442, n443, n444, n446, n447, n448, n449,
    n451, n452, n453, n454, n455, n457, n458, n459, n460, n462, n463, n464,
    n465, n466, n468, n469, n470, n471, n473, n474, n475, n476, n477, n479,
    n480, n481, n482, n484, n485, n486, n487, n489, n490, n491, n492, n494,
    n495, n496, n497, n499, n500, n501, n502, n504, n505, n506, n507, n509,
    n510, n511, n512, n514, n515, n516, n517, n519, n520, n521, n522, n524,
    n525, n526, n527, n529, n530, n531, n532, n534, n535, n536, n537, n539,
    n540, n541, n542, n543, n545, n546, n547, n548, n549, n551, n552, n553,
    n554, n555, n557, n558, n559, n560, n561, n563, n564, n565, n566, n567,
    n569, n570, n571, n572, n573, n575, n576, n577, n578, n579, n581, n582,
    n583, n584, n585;
  assign n206 = ~\V138(2)  & ~\V138(0) ;
  assign n207 = \V138(4)  & n206;
  assign n208 = ~\V138(2)  & \V138(0) ;
  assign n209 = \V138(4)  & n208;
  assign n210 = \V138(2)  & \V138(0) ;
  assign n211 = \V138(2)  & ~\V138(4) ;
  assign n212 = \V96(3)  & n207;
  assign n213 = \V131(3)  & n209;
  assign n214 = ~\V131(3)  & n210;
  assign n215 = ~n211 & ~n214;
  assign n216 = ~n213 & n215;
  assign \V198(7)  = n212 | ~n216;
  assign n218 = \V96(2)  & n207;
  assign n219 = \V131(2)  & n209;
  assign n220 = ~\V131(2)  & n210;
  assign n221 = ~n211 & ~n220;
  assign n222 = ~n219 & n221;
  assign \V198(6)  = n218 | ~n222;
  assign n224 = \V96(5)  & n207;
  assign n225 = \V131(5)  & n209;
  assign n226 = ~\V131(5)  & n210;
  assign n227 = ~n211 & ~n226;
  assign n228 = ~n225 & n227;
  assign \V198(9)  = n224 | ~n228;
  assign n230 = \V96(4)  & n207;
  assign n231 = \V131(4)  & n209;
  assign n232 = ~\V131(4)  & n210;
  assign n233 = ~n211 & ~n232;
  assign n234 = ~n231 & n233;
  assign \V198(8)  = n230 | ~n234;
  assign n236 = ~\V64(3)  & n210;
  assign n237 = \V64(3)  & n208;
  assign n238 = \V32(3)  & n206;
  assign n239 = ~n237 & ~n238;
  assign \V166(3)  = n236 | ~n239;
  assign n241 = ~\V64(2)  & n210;
  assign n242 = \V64(2)  & n208;
  assign n243 = \V32(2)  & n206;
  assign n244 = ~n242 & ~n243;
  assign \V166(2)  = n241 | ~n244;
  assign n246 = ~\V64(5)  & n210;
  assign n247 = \V64(5)  & n208;
  assign n248 = \V32(5)  & n206;
  assign n249 = ~n247 & ~n248;
  assign \V166(5)  = n246 | ~n249;
  assign n251 = ~\V64(4)  & n210;
  assign n252 = \V64(4)  & n208;
  assign n253 = \V32(4)  & n206;
  assign n254 = ~n252 & ~n253;
  assign \V166(4)  = n251 | ~n254;
  assign n256 = ~\V64(1)  & n210;
  assign n257 = \V64(1)  & n208;
  assign n258 = \V32(1)  & n206;
  assign n259 = ~n257 & ~n258;
  assign \V166(1)  = n256 | ~n259;
  assign n261 = ~\V64(0)  & n210;
  assign n262 = \V64(0)  & n208;
  assign n263 = \V32(0)  & n206;
  assign n264 = ~n262 & ~n263;
  assign \V166(0)  = n261 | ~n264;
  assign n266 = ~\V64(7)  & n210;
  assign n267 = \V64(7)  & n208;
  assign n268 = \V32(7)  & n206;
  assign n269 = ~n267 & ~n268;
  assign \V166(7)  = n266 | ~n269;
  assign n271 = ~\V64(6)  & n210;
  assign n272 = \V64(6)  & n208;
  assign n273 = \V32(6)  & n206;
  assign n274 = ~n272 & ~n273;
  assign \V166(6)  = n271 | ~n274;
  assign n276 = ~\V64(9)  & n210;
  assign n277 = \V64(9)  & n208;
  assign n278 = \V32(9)  & n206;
  assign n279 = ~n277 & ~n278;
  assign \V166(9)  = n276 | ~n279;
  assign n281 = \V96(23)  & n207;
  assign n282 = \V131(23)  & n209;
  assign n283 = ~\V131(23)  & n210;
  assign n284 = ~n211 & ~n283;
  assign n285 = ~n282 & n284;
  assign \V198(27)  = n281 | ~n285;
  assign n287 = ~\V64(8)  & n210;
  assign n288 = \V64(8)  & n208;
  assign n289 = \V32(8)  & n206;
  assign n290 = ~n288 & ~n289;
  assign \V166(8)  = n287 | ~n290;
  assign n292 = \V138(3)  & n208;
  assign n293 = \V138(3)  & n206;
  assign n294 = ~\V138(3)  & \V138(2) ;
  assign n295 = \V131(31)  & n292;
  assign n296 = \V96(31)  & n293;
  assign n297 = ~\V131(31)  & n210;
  assign n298 = ~n294 & ~n297;
  assign n299 = ~n296 & n298;
  assign \V205(3)  = n295 | ~n299;
  assign n301 = \V96(22)  & n207;
  assign n302 = \V131(22)  & n209;
  assign n303 = ~\V131(22)  & n210;
  assign n304 = ~n211 & ~n303;
  assign n305 = ~n302 & n304;
  assign \V198(26)  = n301 | ~n305;
  assign n307 = \V131(30)  & n292;
  assign n308 = \V96(30)  & n293;
  assign n309 = ~\V131(30)  & n210;
  assign n310 = ~n294 & ~n309;
  assign n311 = ~n308 & n310;
  assign \V205(2)  = n307 | ~n311;
  assign n313 = \V96(25)  & n207;
  assign n314 = \V131(25)  & n209;
  assign n315 = ~\V131(25)  & n210;
  assign n316 = ~n211 & ~n315;
  assign n317 = ~n314 & n316;
  assign \V198(29)  = n313 | ~n317;
  assign n319 = \V133(1)  & n292;
  assign n320 = \V98(0)  & n293;
  assign n321 = ~\V133(1)  & n210;
  assign n322 = ~n294 & ~n321;
  assign n323 = ~n320 & n322;
  assign \V205(5)  = n319 | ~n323;
  assign n325 = \V96(24)  & n207;
  assign n326 = \V131(24)  & n209;
  assign n327 = ~\V131(24)  & n210;
  assign n328 = ~n211 & ~n327;
  assign n329 = ~n326 & n328;
  assign \V198(28)  = n325 | ~n329;
  assign n331 = \V133(0)  & n292;
  assign n332 = \V97(0)  & n293;
  assign n333 = ~\V133(0)  & n210;
  assign n334 = ~n294 & ~n333;
  assign n335 = ~n332 & n334;
  assign \V205(4)  = n331 | ~n335;
  assign n337 = \V131(29)  & n292;
  assign n338 = \V96(29)  & n293;
  assign n339 = ~\V131(29)  & n210;
  assign n340 = ~n294 & ~n339;
  assign n341 = ~n338 & n340;
  assign \V205(1)  = n337 | ~n341;
  assign n343 = \V131(28)  & n292;
  assign n344 = \V96(28)  & n293;
  assign n345 = ~\V131(28)  & n210;
  assign n346 = ~n294 & ~n345;
  assign n347 = ~n344 & n346;
  assign \V205(0)  = n343 | ~n347;
  assign n349 = \V96(17)  & n207;
  assign n350 = \V131(17)  & n209;
  assign n351 = ~\V131(17)  & n210;
  assign n352 = ~n211 & ~n351;
  assign n353 = ~n350 & n352;
  assign \V198(21)  = n349 | ~n353;
  assign n355 = \V96(16)  & n207;
  assign n356 = \V131(16)  & n209;
  assign n357 = ~\V131(16)  & n210;
  assign n358 = ~n211 & ~n357;
  assign n359 = ~n356 & n358;
  assign \V198(20)  = n355 | ~n359;
  assign n361 = \V96(19)  & n207;
  assign n362 = \V131(19)  & n209;
  assign n363 = ~\V131(19)  & n210;
  assign n364 = ~n211 & ~n363;
  assign n365 = ~n362 & n364;
  assign \V198(23)  = n361 | ~n365;
  assign n367 = \V96(18)  & n207;
  assign n368 = \V131(18)  & n209;
  assign n369 = ~\V131(18)  & n210;
  assign n370 = ~n211 & ~n369;
  assign n371 = ~n368 & n370;
  assign \V198(22)  = n367 | ~n371;
  assign n373 = \V138(3)  & \V138(0) ;
  assign n374 = \V134(0)  & n373;
  assign n375 = \V99(0)  & n293;
  assign \V205(6)  = n374 | n375;
  assign n377 = \V96(21)  & n207;
  assign n378 = \V131(21)  & n209;
  assign n379 = ~\V131(21)  & n210;
  assign n380 = ~n211 & ~n379;
  assign n381 = ~n378 & n380;
  assign \V198(25)  = n377 | ~n381;
  assign n383 = \V96(20)  & n207;
  assign n384 = \V131(20)  & n209;
  assign n385 = ~\V131(20)  & n210;
  assign n386 = ~n211 & ~n385;
  assign n387 = ~n384 & n386;
  assign \V198(24)  = n383 | ~n387;
  assign n389 = \V96(13)  & n207;
  assign n390 = \V131(13)  & n209;
  assign n391 = ~\V131(13)  & n210;
  assign n392 = ~n211 & ~n391;
  assign n393 = ~n390 & n392;
  assign \V198(17)  = n389 | ~n393;
  assign n395 = \V96(12)  & n207;
  assign n396 = \V131(12)  & n209;
  assign n397 = ~\V131(12)  & n210;
  assign n398 = ~n211 & ~n397;
  assign n399 = ~n396 & n398;
  assign \V198(16)  = n395 | ~n399;
  assign n401 = ~\V64(27)  & n210;
  assign n402 = \V64(27)  & n208;
  assign n403 = \V32(27)  & n206;
  assign n404 = ~n402 & ~n403;
  assign \V166(27)  = n401 | ~n404;
  assign n406 = \V96(15)  & n207;
  assign n407 = \V131(15)  & n209;
  assign n408 = ~\V131(15)  & n210;
  assign n409 = ~n211 & ~n408;
  assign n410 = ~n407 & n409;
  assign \V198(19)  = n406 | ~n410;
  assign n412 = ~\V64(26)  & n210;
  assign n413 = \V64(26)  & n208;
  assign n414 = \V32(26)  & n206;
  assign n415 = ~n413 & ~n414;
  assign \V166(26)  = n412 | ~n415;
  assign n417 = \V96(14)  & n207;
  assign n418 = \V131(14)  & n209;
  assign n419 = ~\V131(14)  & n210;
  assign n420 = ~n211 & ~n419;
  assign n421 = ~n418 & n420;
  assign \V198(18)  = n417 | ~n421;
  assign n423 = \V96(7)  & n207;
  assign n424 = \V131(7)  & n209;
  assign n425 = ~\V131(7)  & n210;
  assign n426 = ~n211 & ~n425;
  assign n427 = ~n424 & n426;
  assign \V198(11)  = n423 | ~n427;
  assign n429 = \V96(6)  & n207;
  assign n430 = \V131(6)  & n209;
  assign n431 = ~\V131(6)  & n210;
  assign n432 = ~n211 & ~n431;
  assign n433 = ~n430 & n432;
  assign \V198(10)  = n429 | ~n433;
  assign n435 = ~\V64(21)  & n210;
  assign n436 = \V64(21)  & n208;
  assign n437 = \V32(21)  & n206;
  assign n438 = ~n436 & ~n437;
  assign \V166(21)  = n435 | ~n438;
  assign n440 = \V96(9)  & n207;
  assign n441 = \V131(9)  & n209;
  assign n442 = ~\V131(9)  & n210;
  assign n443 = ~n211 & ~n442;
  assign n444 = ~n441 & n443;
  assign \V198(13)  = n440 | ~n444;
  assign n446 = ~\V64(20)  & n210;
  assign n447 = \V64(20)  & n208;
  assign n448 = \V32(20)  & n206;
  assign n449 = ~n447 & ~n448;
  assign \V166(20)  = n446 | ~n449;
  assign n451 = \V96(8)  & n207;
  assign n452 = \V131(8)  & n209;
  assign n453 = ~\V131(8)  & n210;
  assign n454 = ~n211 & ~n453;
  assign n455 = ~n452 & n454;
  assign \V198(12)  = n451 | ~n455;
  assign n457 = ~\V64(23)  & n210;
  assign n458 = \V64(23)  & n208;
  assign n459 = \V32(23)  & n206;
  assign n460 = ~n458 & ~n459;
  assign \V166(23)  = n457 | ~n460;
  assign n462 = \V96(11)  & n207;
  assign n463 = \V131(11)  & n209;
  assign n464 = ~\V131(11)  & n210;
  assign n465 = ~n211 & ~n464;
  assign n466 = ~n463 & n465;
  assign \V198(15)  = n462 | ~n466;
  assign n468 = ~\V64(22)  & n210;
  assign n469 = \V64(22)  & n208;
  assign n470 = \V32(22)  & n206;
  assign n471 = ~n469 & ~n470;
  assign \V166(22)  = n468 | ~n471;
  assign n473 = \V96(10)  & n207;
  assign n474 = \V131(10)  & n209;
  assign n475 = ~\V131(10)  & n210;
  assign n476 = ~n211 & ~n475;
  assign n477 = ~n474 & n476;
  assign \V198(14)  = n473 | ~n477;
  assign n479 = ~\V64(25)  & n210;
  assign n480 = \V64(25)  & n208;
  assign n481 = \V32(25)  & n206;
  assign n482 = ~n480 & ~n481;
  assign \V166(25)  = n479 | ~n482;
  assign n484 = ~\V64(24)  & n210;
  assign n485 = \V64(24)  & n208;
  assign n486 = \V32(24)  & n206;
  assign n487 = ~n485 & ~n486;
  assign \V166(24)  = n484 | ~n487;
  assign n489 = ~\V64(17)  & n210;
  assign n490 = \V64(17)  & n208;
  assign n491 = \V32(17)  & n206;
  assign n492 = ~n490 & ~n491;
  assign \V166(17)  = n489 | ~n492;
  assign n494 = ~\V64(16)  & n210;
  assign n495 = \V64(16)  & n208;
  assign n496 = \V32(16)  & n206;
  assign n497 = ~n495 & ~n496;
  assign \V166(16)  = n494 | ~n497;
  assign n499 = ~\V64(19)  & n210;
  assign n500 = \V64(19)  & n208;
  assign n501 = \V32(19)  & n206;
  assign n502 = ~n500 & ~n501;
  assign \V166(19)  = n499 | ~n502;
  assign n504 = ~\V64(18)  & n210;
  assign n505 = \V64(18)  & n208;
  assign n506 = \V32(18)  & n206;
  assign n507 = ~n505 & ~n506;
  assign \V166(18)  = n504 | ~n507;
  assign n509 = ~\V64(11)  & n210;
  assign n510 = \V64(11)  & n208;
  assign n511 = \V32(11)  & n206;
  assign n512 = ~n510 & ~n511;
  assign \V166(11)  = n509 | ~n512;
  assign n514 = ~\V64(10)  & n210;
  assign n515 = \V64(10)  & n208;
  assign n516 = \V32(10)  & n206;
  assign n517 = ~n515 & ~n516;
  assign \V166(10)  = n514 | ~n517;
  assign n519 = ~\V64(13)  & n210;
  assign n520 = \V64(13)  & n208;
  assign n521 = \V32(13)  & n206;
  assign n522 = ~n520 & ~n521;
  assign \V166(13)  = n519 | ~n522;
  assign n524 = ~\V64(12)  & n210;
  assign n525 = \V64(12)  & n208;
  assign n526 = \V32(12)  & n206;
  assign n527 = ~n525 & ~n526;
  assign \V166(12)  = n524 | ~n527;
  assign n529 = ~\V64(15)  & n210;
  assign n530 = \V64(15)  & n208;
  assign n531 = \V32(15)  & n206;
  assign n532 = ~n530 & ~n531;
  assign \V166(15)  = n529 | ~n532;
  assign n534 = ~\V64(14)  & n210;
  assign n535 = \V64(14)  & n208;
  assign n536 = \V32(14)  & n206;
  assign n537 = ~n535 & ~n536;
  assign \V166(14)  = n534 | ~n537;
  assign n539 = \V32(31)  & n207;
  assign n540 = \V64(31)  & n209;
  assign n541 = ~\V64(31)  & n210;
  assign n542 = ~n211 & ~n541;
  assign n543 = ~n540 & n542;
  assign \V198(3)  = n539 | ~n543;
  assign n545 = \V32(30)  & n207;
  assign n546 = \V64(30)  & n209;
  assign n547 = ~\V64(30)  & n210;
  assign n548 = ~n211 & ~n547;
  assign n549 = ~n546 & n548;
  assign \V198(2)  = n545 | ~n549;
  assign n551 = \V96(1)  & n207;
  assign n552 = \V131(1)  & n209;
  assign n553 = ~\V131(1)  & n210;
  assign n554 = ~n211 & ~n553;
  assign n555 = ~n552 & n554;
  assign \V198(5)  = n551 | ~n555;
  assign n557 = \V96(0)  & n207;
  assign n558 = \V131(0)  & n209;
  assign n559 = ~\V131(0)  & n210;
  assign n560 = ~n211 & ~n559;
  assign n561 = ~n558 & n560;
  assign \V198(4)  = n557 | ~n561;
  assign n563 = \V96(27)  & n207;
  assign n564 = \V131(27)  & n209;
  assign n565 = ~\V131(27)  & n210;
  assign n566 = ~n211 & ~n565;
  assign n567 = ~n564 & n566;
  assign \V198(31)  = n563 | ~n567;
  assign n569 = \V96(26)  & n207;
  assign n570 = \V131(26)  & n209;
  assign n571 = ~\V131(26)  & n210;
  assign n572 = ~n211 & ~n571;
  assign n573 = ~n570 & n572;
  assign \V198(30)  = n569 | ~n573;
  assign n575 = \V32(29)  & n207;
  assign n576 = \V64(29)  & n209;
  assign n577 = ~\V64(29)  & n210;
  assign n578 = ~n211 & ~n577;
  assign n579 = ~n576 & n578;
  assign \V198(1)  = n575 | ~n579;
  assign n581 = \V32(28)  & n207;
  assign n582 = \V64(28)  & n209;
  assign n583 = ~\V64(28)  & n210;
  assign n584 = ~n211 & ~n583;
  assign n585 = ~n582 & n584;
  assign \V198(0)  = n581 | ~n585;
endmodule


