// Benchmark "dalu" written by ABC on Tue May 16 16:07:48 2017

module dalu ( 
    inA10, inA11, inA12, inA13, inA14, inA15, inB10, inB11, inB12, inB13,
    inB14, inB15, inC10, inC11, inC12, inC13, inC14, inC15, inD10, inD11,
    inD12, inD13, inD14, inD15, inA0, inA1, inA2, inA3, inA4, inA5, inA6,
    inA7, inA8, inA9, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7, inB8,
    inB9, inC0, inC1, inC2, inC3, inC4, inC5, inC6, inC7, inC8, inC9, inD0,
    inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, inD9, sh0, sh1, sh2,
    musel1, musel2, musel3, musel4, opsel0, opsel1, opsel2, opsel3,
    O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15  );
  input  inA10, inA11, inA12, inA13, inA14, inA15, inB10, inB11, inB12,
    inB13, inB14, inB15, inC10, inC11, inC12, inC13, inC14, inC15, inD10,
    inD11, inD12, inD13, inD14, inD15, inA0, inA1, inA2, inA3, inA4, inA5,
    inA6, inA7, inA8, inA9, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7,
    inB8, inB9, inC0, inC1, inC2, inC3, inC4, inC5, inC6, inC7, inC8, inC9,
    inD0, inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, inD9, sh0, sh1,
    sh2, musel1, musel2, musel3, musel4, opsel0, opsel1, opsel2, opsel3;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
  assign n92 = inC0 & musel2;
  assign n93 = inA0 & ~musel2;
  assign n94 = musel1 & n93;
  assign n95 = ~musel1 & n92;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~musel3 & musel4;
  assign n98 = ~n96 & n97;
  assign n99 = inC15 & musel2;
  assign n100 = inA15 & ~musel2;
  assign n101 = musel1 & n100;
  assign n102 = ~musel1 & n99;
  assign n103 = ~n101 & ~n102;
  assign n104 = n97 & ~n103;
  assign n105 = ~n98 & n104;
  assign n106 = n98 & ~n104;
  assign n107 = ~n105 & ~n106;
  assign n108 = n104 & n107;
  assign n109 = ~n104 & ~n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = opsel2 & ~n110;
  assign n112 = ~opsel0 & ~opsel1;
  assign n113 = n111 & n112;
  assign n114 = musel3 & ~musel4;
  assign n115 = inD0 & musel2;
  assign n116 = ~musel1 & musel2;
  assign n117 = musel1 & ~musel2;
  assign n118 = ~n116 & ~n117;
  assign n119 = ~inB0 & ~n115;
  assign n120 = ~inB0 & ~musel1;
  assign n121 = ~n115 & n118;
  assign n122 = ~musel1 & n118;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~n120 & n123;
  assign n125 = ~n119 & n124;
  assign n126 = ~musel1 & ~musel2;
  assign n127 = inD0 & musel4;
  assign n128 = ~musel3 & n127;
  assign n129 = n126 & n128;
  assign n130 = n114 & n125;
  assign n131 = ~n129 & ~n130;
  assign n132 = inD4 & musel2;
  assign n133 = ~inB4 & ~n132;
  assign n134 = ~inB4 & ~musel1;
  assign n135 = n118 & ~n132;
  assign n136 = ~n122 & ~n135;
  assign n137 = ~n134 & n136;
  assign n138 = ~n133 & n137;
  assign n139 = inD4 & musel4;
  assign n140 = ~musel3 & n139;
  assign n141 = n126 & n140;
  assign n142 = n114 & n138;
  assign n143 = ~n141 & ~n142;
  assign n144 = sh2 & ~n143;
  assign n145 = ~sh2 & ~n131;
  assign n146 = ~n144 & ~n145;
  assign n147 = inD2 & musel2;
  assign n148 = ~inB2 & ~n147;
  assign n149 = ~inB2 & ~musel1;
  assign n150 = n118 & ~n147;
  assign n151 = ~n122 & ~n150;
  assign n152 = ~n149 & n151;
  assign n153 = ~n148 & n152;
  assign n154 = inD2 & musel4;
  assign n155 = ~musel3 & n154;
  assign n156 = n126 & n155;
  assign n157 = n114 & n153;
  assign n158 = ~n156 & ~n157;
  assign n159 = inD8 & musel2;
  assign n160 = ~inB8 & ~n159;
  assign n161 = ~inB8 & ~musel1;
  assign n162 = n118 & ~n159;
  assign n163 = ~n122 & ~n162;
  assign n164 = ~n161 & n163;
  assign n165 = ~n160 & n164;
  assign n166 = inD8 & musel4;
  assign n167 = ~musel3 & n166;
  assign n168 = n126 & n167;
  assign n169 = n114 & n165;
  assign n170 = ~n168 & ~n169;
  assign n171 = sh2 & ~n170;
  assign n172 = ~sh2 & ~n158;
  assign n173 = ~n171 & ~n172;
  assign n174 = n146 & n173;
  assign n175 = ~sh1 & n146;
  assign n176 = sh1 & n173;
  assign n177 = ~n175 & ~n176;
  assign n178 = ~n174 & n177;
  assign n179 = inD1 & musel2;
  assign n180 = ~inB1 & ~n179;
  assign n181 = ~inB1 & ~musel1;
  assign n182 = n118 & ~n179;
  assign n183 = ~n122 & ~n182;
  assign n184 = ~n181 & n183;
  assign n185 = ~n180 & n184;
  assign n186 = inD1 & musel4;
  assign n187 = ~musel3 & n186;
  assign n188 = n126 & n187;
  assign n189 = n114 & n185;
  assign n190 = ~n188 & ~n189;
  assign n191 = inD5 & musel2;
  assign n192 = ~inB5 & ~n191;
  assign n193 = ~inB5 & ~musel1;
  assign n194 = n118 & ~n191;
  assign n195 = ~n122 & ~n194;
  assign n196 = ~n193 & n195;
  assign n197 = ~n192 & n196;
  assign n198 = inD5 & musel4;
  assign n199 = ~musel3 & n198;
  assign n200 = n126 & n199;
  assign n201 = n114 & n197;
  assign n202 = ~n200 & ~n201;
  assign n203 = sh2 & ~n202;
  assign n204 = ~sh2 & ~n190;
  assign n205 = ~n203 & ~n204;
  assign n206 = inD3 & musel2;
  assign n207 = ~inB3 & ~n206;
  assign n208 = ~inB3 & ~musel1;
  assign n209 = n118 & ~n206;
  assign n210 = ~n122 & ~n209;
  assign n211 = ~n208 & n210;
  assign n212 = ~n207 & n211;
  assign n213 = inD3 & musel4;
  assign n214 = ~musel3 & n213;
  assign n215 = n126 & n214;
  assign n216 = n114 & n212;
  assign n217 = ~n215 & ~n216;
  assign n218 = sh2 & ~n131;
  assign n219 = ~sh2 & ~n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = n205 & n220;
  assign n222 = ~sh1 & n205;
  assign n223 = sh1 & n220;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~n221 & n224;
  assign n226 = ~sh0 & n178;
  assign n227 = sh0 & n225;
  assign n228 = ~n226 & ~n227;
  assign n229 = n110 & n228;
  assign n230 = ~opsel2 & n110;
  assign n231 = opsel2 & n228;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n229 & n232;
  assign n234 = ~n113 & ~n233;
  assign n235 = n112 & ~n113;
  assign n236 = ~n234 & ~n235;
  assign n237 = opsel0 & opsel1;
  assign n238 = ~n112 & ~n237;
  assign n239 = opsel2 & opsel3;
  assign n240 = ~opsel1 & ~opsel3;
  assign n241 = opsel1 & ~opsel2;
  assign n242 = ~n240 & ~n241;
  assign n243 = ~opsel0 & n242;
  assign n244 = ~n239 & n243;
  assign n245 = ~inA0 & ~n92;
  assign n246 = ~inA0 & ~musel1;
  assign n247 = ~n92 & n118;
  assign n248 = ~n122 & ~n247;
  assign n249 = ~n246 & n248;
  assign n250 = ~n245 & n249;
  assign n251 = n114 & n250;
  assign n252 = inC0 & musel4;
  assign n253 = ~musel3 & n252;
  assign n254 = ~musel2 & n253;
  assign n255 = ~musel1 & n254;
  assign n256 = ~n251 & ~n255;
  assign n257 = ~n244 & ~n256;
  assign n258 = n244 & n256;
  assign n259 = ~n257 & ~n258;
  assign n260 = inB0 & ~musel3;
  assign n261 = musel2 & n260;
  assign n262 = inD0 & musel3;
  assign n263 = ~musel2 & n262;
  assign n264 = ~musel1 & n261;
  assign n265 = ~musel1 & n263;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~inA0 & ~musel2;
  assign n268 = ~inC0 & musel2;
  assign n269 = ~inA0 & ~inC0;
  assign n270 = ~n268 & ~n269;
  assign n271 = ~n267 & n270;
  assign n272 = musel1 & ~musel3;
  assign n273 = n271 & n272;
  assign n274 = n266 & ~n273;
  assign n275 = ~musel4 & ~n274;
  assign n276 = n259 & n275;
  assign n277 = ~n259 & ~n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = opsel2 & ~opsel3;
  assign n280 = opsel1 & n279;
  assign n281 = ~opsel2 & opsel3;
  assign n282 = ~opsel1 & n281;
  assign n283 = ~n280 & ~n282;
  assign n284 = ~opsel0 & ~n283;
  assign n285 = n278 & n284;
  assign n286 = n278 & ~n285;
  assign n287 = n284 & ~n285;
  assign n288 = ~n286 & ~n287;
  assign n289 = n238 & n288;
  assign n290 = n112 & ~n228;
  assign n291 = ~n289 & ~n290;
  assign n292 = n281 & ~n291;
  assign n293 = ~opsel3 & n236;
  assign O0 = n292 | n293;
  assign n295 = n104 & ~n107;
  assign n296 = inC1 & musel2;
  assign n297 = inA1 & ~musel2;
  assign n298 = musel1 & n297;
  assign n299 = ~musel1 & n296;
  assign n300 = ~n298 & ~n299;
  assign n301 = n97 & ~n300;
  assign n302 = n104 & ~n301;
  assign n303 = ~n104 & n301;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~n295 & ~n304;
  assign n306 = n295 & n304;
  assign n307 = ~n305 & ~n306;
  assign n308 = opsel2 & ~n307;
  assign n309 = n112 & n308;
  assign n310 = inD9 & musel2;
  assign n311 = ~inB9 & ~n310;
  assign n312 = ~inB9 & ~musel1;
  assign n313 = n118 & ~n310;
  assign n314 = ~n122 & ~n313;
  assign n315 = ~n312 & n314;
  assign n316 = ~n311 & n315;
  assign n317 = inD9 & musel4;
  assign n318 = ~musel3 & n317;
  assign n319 = n126 & n318;
  assign n320 = n114 & n316;
  assign n321 = ~n319 & ~n320;
  assign n322 = sh2 & ~n321;
  assign n323 = ~n219 & ~n322;
  assign n324 = n205 & n323;
  assign n325 = sh1 & n323;
  assign n326 = ~n222 & ~n325;
  assign n327 = ~n324 & n326;
  assign n328 = inD6 & musel2;
  assign n329 = ~inB6 & ~n328;
  assign n330 = ~inB6 & ~musel1;
  assign n331 = n118 & ~n328;
  assign n332 = ~n122 & ~n331;
  assign n333 = ~n330 & n332;
  assign n334 = ~n329 & n333;
  assign n335 = inD6 & musel4;
  assign n336 = ~musel3 & n335;
  assign n337 = n126 & n336;
  assign n338 = n114 & n334;
  assign n339 = ~n337 & ~n338;
  assign n340 = sh2 & ~n339;
  assign n341 = ~n172 & ~n340;
  assign n342 = sh2 & ~n190;
  assign n343 = ~sh2 & ~n143;
  assign n344 = ~n342 & ~n343;
  assign n345 = n341 & n344;
  assign n346 = ~sh1 & n341;
  assign n347 = sh1 & n344;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n345 & n348;
  assign n350 = ~sh0 & n327;
  assign n351 = sh0 & n349;
  assign n352 = ~n350 & ~n351;
  assign n353 = n307 & n352;
  assign n354 = ~opsel2 & n307;
  assign n355 = opsel2 & n352;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n353 & n356;
  assign n358 = ~n309 & ~n357;
  assign n359 = n112 & ~n309;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~inA1 & ~n296;
  assign n362 = ~inA1 & ~musel1;
  assign n363 = n118 & ~n296;
  assign n364 = ~n122 & ~n363;
  assign n365 = ~n362 & n364;
  assign n366 = ~n361 & n365;
  assign n367 = n114 & n366;
  assign n368 = inC1 & musel4;
  assign n369 = ~musel3 & n368;
  assign n370 = ~musel2 & n369;
  assign n371 = ~musel1 & n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~n244 & ~n372;
  assign n374 = n244 & n372;
  assign n375 = ~n373 & ~n374;
  assign n376 = inB1 & ~musel3;
  assign n377 = musel2 & n376;
  assign n378 = inD1 & musel3;
  assign n379 = ~musel2 & n378;
  assign n380 = ~musel1 & n377;
  assign n381 = ~musel1 & n379;
  assign n382 = ~n380 & ~n381;
  assign n383 = ~inA1 & ~musel2;
  assign n384 = ~inC1 & musel2;
  assign n385 = ~inA1 & ~inC1;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n383 & n386;
  assign n388 = n272 & n387;
  assign n389 = n382 & ~n388;
  assign n390 = ~musel4 & ~n389;
  assign n391 = n375 & n390;
  assign n392 = ~n375 & ~n390;
  assign n393 = ~n391 & ~n392;
  assign n394 = n259 & ~n275;
  assign n395 = n284 & ~n394;
  assign n396 = ~n259 & n275;
  assign n397 = n393 & n395;
  assign n398 = n393 & n396;
  assign n399 = ~n397 & ~n398;
  assign n400 = ~n284 & ~n396;
  assign n401 = ~n394 & ~n400;
  assign n402 = n393 & n399;
  assign n403 = n399 & n401;
  assign n404 = ~n402 & ~n403;
  assign n405 = n238 & n404;
  assign n406 = n112 & ~n352;
  assign n407 = ~n405 & ~n406;
  assign n408 = n281 & ~n407;
  assign n409 = ~opsel3 & n360;
  assign O1 = n408 | n409;
  assign n411 = n104 & ~n304;
  assign n412 = ~n107 & n411;
  assign n413 = inC2 & musel2;
  assign n414 = inA2 & ~musel2;
  assign n415 = musel1 & n414;
  assign n416 = ~musel1 & n413;
  assign n417 = ~n415 & ~n416;
  assign n418 = n97 & ~n417;
  assign n419 = n104 & ~n418;
  assign n420 = ~n104 & n418;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n412 & ~n421;
  assign n423 = n412 & n421;
  assign n424 = ~n422 & ~n423;
  assign n425 = opsel2 & ~n424;
  assign n426 = n112 & n425;
  assign n427 = inD10 & musel2;
  assign n428 = ~inB10 & ~n427;
  assign n429 = ~inB10 & ~musel1;
  assign n430 = n118 & ~n427;
  assign n431 = ~n122 & ~n430;
  assign n432 = ~n429 & n431;
  assign n433 = ~n428 & n432;
  assign n434 = inD10 & musel4;
  assign n435 = ~musel3 & n434;
  assign n436 = n126 & n435;
  assign n437 = n114 & n433;
  assign n438 = ~n436 & ~n437;
  assign n439 = sh2 & ~n438;
  assign n440 = ~n343 & ~n439;
  assign n441 = n341 & n440;
  assign n442 = sh1 & n440;
  assign n443 = ~n346 & ~n442;
  assign n444 = ~n441 & n443;
  assign n445 = inD7 & musel2;
  assign n446 = ~inB7 & ~n445;
  assign n447 = ~inB7 & ~musel1;
  assign n448 = n118 & ~n445;
  assign n449 = ~n122 & ~n448;
  assign n450 = ~n447 & n449;
  assign n451 = ~n446 & n450;
  assign n452 = inD7 & musel4;
  assign n453 = ~musel3 & n452;
  assign n454 = n126 & n453;
  assign n455 = n114 & n451;
  assign n456 = ~n454 & ~n455;
  assign n457 = sh2 & ~n456;
  assign n458 = ~n219 & ~n457;
  assign n459 = sh2 & ~n158;
  assign n460 = ~sh2 & ~n202;
  assign n461 = ~n459 & ~n460;
  assign n462 = n458 & n461;
  assign n463 = ~sh1 & n458;
  assign n464 = sh1 & n461;
  assign n465 = ~n463 & ~n464;
  assign n466 = ~n462 & n465;
  assign n467 = ~sh0 & n444;
  assign n468 = sh0 & n466;
  assign n469 = ~n467 & ~n468;
  assign n470 = n424 & n469;
  assign n471 = ~opsel2 & n424;
  assign n472 = opsel2 & n469;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~n470 & n473;
  assign n475 = ~n426 & ~n474;
  assign n476 = n112 & ~n426;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~inA2 & ~n413;
  assign n479 = ~inA2 & ~musel1;
  assign n480 = n118 & ~n413;
  assign n481 = ~n122 & ~n480;
  assign n482 = ~n479 & n481;
  assign n483 = ~n478 & n482;
  assign n484 = n114 & n483;
  assign n485 = inC2 & musel4;
  assign n486 = ~musel3 & n485;
  assign n487 = ~musel2 & n486;
  assign n488 = ~musel1 & n487;
  assign n489 = ~n484 & ~n488;
  assign n490 = ~n244 & ~n489;
  assign n491 = n244 & n489;
  assign n492 = ~n490 & ~n491;
  assign n493 = inB2 & ~musel3;
  assign n494 = musel2 & n493;
  assign n495 = inD2 & musel3;
  assign n496 = ~musel2 & n495;
  assign n497 = ~musel1 & n494;
  assign n498 = ~musel1 & n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~inA2 & ~musel2;
  assign n501 = ~inC2 & musel2;
  assign n502 = ~inA2 & ~inC2;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n500 & n503;
  assign n505 = n272 & n504;
  assign n506 = n499 & ~n505;
  assign n507 = ~musel4 & ~n506;
  assign n508 = n492 & n507;
  assign n509 = ~n492 & ~n507;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n395 & ~n396;
  assign n512 = n375 & ~n390;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n375 & n390;
  assign n515 = n510 & n513;
  assign n516 = n510 & n514;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n394 & n396;
  assign n519 = ~n395 & ~n518;
  assign n520 = ~n514 & n519;
  assign n521 = ~n512 & ~n520;
  assign n522 = n510 & n517;
  assign n523 = n517 & n521;
  assign n524 = ~n522 & ~n523;
  assign n525 = n238 & n524;
  assign n526 = n112 & ~n469;
  assign n527 = ~n525 & ~n526;
  assign n528 = n281 & ~n527;
  assign n529 = ~opsel3 & n477;
  assign O2 = n528 | n529;
  assign n531 = n104 & ~n421;
  assign n532 = ~n304 & n531;
  assign n533 = ~n107 & n532;
  assign n534 = inC3 & musel2;
  assign n535 = inA3 & ~musel2;
  assign n536 = musel1 & n535;
  assign n537 = ~musel1 & n534;
  assign n538 = ~n536 & ~n537;
  assign n539 = n97 & ~n538;
  assign n540 = n104 & ~n539;
  assign n541 = ~n104 & n539;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~n533 & ~n542;
  assign n544 = n533 & n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = opsel2 & ~n545;
  assign n547 = n112 & n546;
  assign n548 = inD11 & musel2;
  assign n549 = ~inB11 & ~n548;
  assign n550 = ~inB11 & ~musel1;
  assign n551 = n118 & ~n548;
  assign n552 = ~n122 & ~n551;
  assign n553 = ~n550 & n552;
  assign n554 = ~n549 & n553;
  assign n555 = inD11 & musel4;
  assign n556 = ~musel3 & n555;
  assign n557 = n126 & n556;
  assign n558 = n114 & n554;
  assign n559 = ~n557 & ~n558;
  assign n560 = sh2 & ~n559;
  assign n561 = ~n460 & ~n560;
  assign n562 = n458 & n561;
  assign n563 = sh1 & n561;
  assign n564 = ~n463 & ~n563;
  assign n565 = ~n562 & n564;
  assign n566 = ~n171 & ~n343;
  assign n567 = sh2 & ~n217;
  assign n568 = ~sh2 & ~n339;
  assign n569 = ~n567 & ~n568;
  assign n570 = n566 & n569;
  assign n571 = ~sh1 & n566;
  assign n572 = sh1 & n569;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n570 & n573;
  assign n575 = ~sh0 & n565;
  assign n576 = sh0 & n574;
  assign n577 = ~n575 & ~n576;
  assign n578 = n545 & n577;
  assign n579 = ~opsel2 & n545;
  assign n580 = opsel2 & n577;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n578 & n581;
  assign n583 = ~n547 & ~n582;
  assign n584 = n112 & ~n547;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~inA3 & ~n534;
  assign n587 = ~inA3 & ~musel1;
  assign n588 = n118 & ~n534;
  assign n589 = ~n122 & ~n588;
  assign n590 = ~n587 & n589;
  assign n591 = ~n586 & n590;
  assign n592 = n114 & n591;
  assign n593 = inC3 & musel4;
  assign n594 = ~musel3 & n593;
  assign n595 = ~musel2 & n594;
  assign n596 = ~musel1 & n595;
  assign n597 = ~n592 & ~n596;
  assign n598 = ~n244 & ~n597;
  assign n599 = n244 & n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = inB3 & ~musel3;
  assign n602 = musel2 & n601;
  assign n603 = inD3 & musel3;
  assign n604 = ~musel2 & n603;
  assign n605 = ~musel1 & n602;
  assign n606 = ~musel1 & n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~inA3 & ~musel2;
  assign n609 = ~inC3 & musel2;
  assign n610 = ~inA3 & ~inC3;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~n608 & n611;
  assign n613 = n272 & n612;
  assign n614 = n607 & ~n613;
  assign n615 = ~musel4 & ~n614;
  assign n616 = n600 & n615;
  assign n617 = ~n600 & ~n615;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n513 & ~n514;
  assign n620 = n492 & ~n507;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n492 & n507;
  assign n623 = n618 & n621;
  assign n624 = n618 & n622;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n521 & ~n622;
  assign n627 = ~n620 & ~n626;
  assign n628 = n625 & n627;
  assign n629 = n618 & n625;
  assign n630 = ~n628 & ~n629;
  assign n631 = n238 & n630;
  assign n632 = n112 & ~n577;
  assign n633 = ~n631 & ~n632;
  assign n634 = n281 & ~n633;
  assign n635 = ~opsel3 & n585;
  assign O3 = n634 | n635;
  assign n637 = ~n421 & ~n542;
  assign n638 = ~n304 & n637;
  assign n639 = ~n107 & n638;
  assign n640 = n104 & n639;
  assign n641 = inC4 & musel2;
  assign n642 = inA4 & ~musel2;
  assign n643 = musel1 & n642;
  assign n644 = ~musel1 & n641;
  assign n645 = ~n643 & ~n644;
  assign n646 = n97 & ~n645;
  assign n647 = n104 & ~n646;
  assign n648 = ~n104 & n646;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n640 & ~n649;
  assign n651 = n640 & n649;
  assign n652 = ~n650 & ~n651;
  assign n653 = opsel2 & ~n652;
  assign n654 = n112 & n653;
  assign n655 = inD12 & musel2;
  assign n656 = ~inB12 & ~n655;
  assign n657 = ~inB12 & ~musel1;
  assign n658 = n118 & ~n655;
  assign n659 = ~n122 & ~n658;
  assign n660 = ~n657 & n659;
  assign n661 = ~n656 & n660;
  assign n662 = inD12 & musel4;
  assign n663 = ~musel3 & n662;
  assign n664 = n126 & n663;
  assign n665 = n114 & n661;
  assign n666 = ~n664 & ~n665;
  assign n667 = sh2 & ~n666;
  assign n668 = ~n568 & ~n667;
  assign n669 = n566 & n668;
  assign n670 = sh1 & n668;
  assign n671 = ~n571 & ~n670;
  assign n672 = ~n669 & n671;
  assign n673 = ~n322 & ~n460;
  assign n674 = ~sh2 & ~n456;
  assign n675 = ~n144 & ~n674;
  assign n676 = n673 & n675;
  assign n677 = ~sh1 & n673;
  assign n678 = sh1 & n675;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n676 & n679;
  assign n681 = ~sh0 & n672;
  assign n682 = sh0 & n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = n652 & n683;
  assign n685 = ~opsel2 & n652;
  assign n686 = opsel2 & n683;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n684 & n687;
  assign n689 = ~n654 & ~n688;
  assign n690 = n112 & ~n654;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~opsel0 & opsel1;
  assign n693 = opsel0 & ~opsel1;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~inA4 & ~n641;
  assign n696 = ~inA4 & ~musel1;
  assign n697 = n118 & ~n641;
  assign n698 = ~n122 & ~n697;
  assign n699 = ~n696 & n698;
  assign n700 = ~n695 & n699;
  assign n701 = n114 & n700;
  assign n702 = inC4 & musel4;
  assign n703 = ~musel3 & n702;
  assign n704 = ~musel2 & n703;
  assign n705 = ~musel1 & n704;
  assign n706 = ~n701 & ~n705;
  assign n707 = ~n244 & ~n706;
  assign n708 = n244 & n706;
  assign n709 = ~n707 & ~n708;
  assign n710 = inB4 & ~musel3;
  assign n711 = musel2 & n710;
  assign n712 = inD4 & musel3;
  assign n713 = ~musel2 & n712;
  assign n714 = ~musel1 & n711;
  assign n715 = ~musel1 & n713;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~inA4 & ~musel2;
  assign n718 = ~inC4 & musel2;
  assign n719 = ~inA4 & ~inC4;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~n717 & n720;
  assign n722 = n272 & n721;
  assign n723 = n716 & ~n722;
  assign n724 = ~musel4 & ~n723;
  assign n725 = n709 & n724;
  assign n726 = ~n709 & ~n724;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n259 & ~n375;
  assign n729 = ~n259 & n390;
  assign n730 = n275 & n390;
  assign n731 = n275 & ~n375;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n729 & n732;
  assign n734 = ~n728 & n733;
  assign n735 = ~n492 & ~n600;
  assign n736 = ~n492 & n615;
  assign n737 = n507 & n615;
  assign n738 = n507 & ~n600;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = ~n735 & n740;
  assign n742 = ~n734 & ~n741;
  assign n743 = ~n396 & ~n514;
  assign n744 = n512 & ~n514;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n492 & n745;
  assign n747 = n507 & n745;
  assign n748 = ~n746 & ~n747;
  assign n749 = n600 & ~n615;
  assign n750 = ~n622 & n748;
  assign n751 = ~n749 & ~n750;
  assign n752 = ~n600 & n615;
  assign n753 = ~n751 & ~n752;
  assign n754 = n284 & n742;
  assign n755 = n753 & ~n754;
  assign n756 = n727 & ~n755;
  assign n757 = ~n727 & n755;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n112 & n694;
  assign n760 = n683 & n694;
  assign n761 = n683 & n758;
  assign n762 = ~n112 & n758;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n760 & n763;
  assign n765 = ~n759 & n764;
  assign n766 = ~opsel3 & n691;
  assign n767 = n281 & n765;
  assign O4 = n766 | n767;
  assign n769 = n640 & ~n649;
  assign n770 = inC5 & musel2;
  assign n771 = inA5 & ~musel2;
  assign n772 = musel1 & n771;
  assign n773 = ~musel1 & n770;
  assign n774 = ~n772 & ~n773;
  assign n775 = n97 & ~n774;
  assign n776 = n104 & ~n775;
  assign n777 = ~n104 & n775;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n769 & ~n778;
  assign n780 = n769 & n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = opsel2 & ~n781;
  assign n783 = n112 & n782;
  assign n784 = inD13 & musel2;
  assign n785 = ~inB13 & ~n784;
  assign n786 = ~inB13 & ~musel1;
  assign n787 = n118 & ~n784;
  assign n788 = ~n122 & ~n787;
  assign n789 = ~n786 & n788;
  assign n790 = ~n785 & n789;
  assign n791 = inD13 & musel4;
  assign n792 = ~musel3 & n791;
  assign n793 = n126 & n792;
  assign n794 = n114 & n790;
  assign n795 = ~n793 & ~n794;
  assign n796 = sh2 & ~n795;
  assign n797 = ~n674 & ~n796;
  assign n798 = n673 & n797;
  assign n799 = sh1 & n797;
  assign n800 = ~n677 & ~n799;
  assign n801 = ~n798 & n800;
  assign n802 = ~n439 & ~n568;
  assign n803 = ~sh2 & ~n170;
  assign n804 = ~n203 & ~n803;
  assign n805 = n802 & n804;
  assign n806 = ~sh1 & n802;
  assign n807 = sh1 & n804;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~n805 & n808;
  assign n810 = ~sh0 & n801;
  assign n811 = sh0 & n809;
  assign n812 = ~n810 & ~n811;
  assign n813 = n781 & n812;
  assign n814 = ~opsel2 & n781;
  assign n815 = opsel2 & n812;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~n813 & n816;
  assign n818 = ~n783 & ~n817;
  assign n819 = n112 & ~n783;
  assign n820 = ~n818 & ~n819;
  assign n821 = ~inA5 & ~n770;
  assign n822 = ~inA5 & ~musel1;
  assign n823 = n118 & ~n770;
  assign n824 = ~n122 & ~n823;
  assign n825 = ~n822 & n824;
  assign n826 = ~n821 & n825;
  assign n827 = n114 & n826;
  assign n828 = inC5 & musel4;
  assign n829 = ~musel3 & n828;
  assign n830 = ~musel2 & n829;
  assign n831 = ~musel1 & n830;
  assign n832 = ~n827 & ~n831;
  assign n833 = ~n244 & ~n832;
  assign n834 = n244 & n832;
  assign n835 = ~n833 & ~n834;
  assign n836 = inB5 & ~musel3;
  assign n837 = musel2 & n836;
  assign n838 = inD5 & musel3;
  assign n839 = ~musel2 & n838;
  assign n840 = ~musel1 & n837;
  assign n841 = ~musel1 & n839;
  assign n842 = ~n840 & ~n841;
  assign n843 = ~inA5 & ~musel2;
  assign n844 = ~inC5 & musel2;
  assign n845 = ~inA5 & ~inC5;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~n843 & n846;
  assign n848 = n272 & n847;
  assign n849 = n842 & ~n848;
  assign n850 = ~musel4 & ~n849;
  assign n851 = n835 & n850;
  assign n852 = ~n835 & ~n850;
  assign n853 = ~n851 & ~n852;
  assign n854 = n709 & ~n724;
  assign n855 = ~n755 & ~n854;
  assign n856 = ~n709 & n724;
  assign n857 = n853 & n855;
  assign n858 = n853 & n856;
  assign n859 = ~n857 & ~n858;
  assign n860 = n755 & ~n856;
  assign n861 = ~n854 & ~n860;
  assign n862 = n853 & n859;
  assign n863 = n859 & n861;
  assign n864 = ~n862 & ~n863;
  assign n865 = n238 & n864;
  assign n866 = n112 & ~n812;
  assign n867 = ~n865 & ~n866;
  assign n868 = n281 & ~n867;
  assign n869 = ~opsel3 & n820;
  assign O5 = n868 | n869;
  assign n871 = n640 & ~n778;
  assign n872 = ~n649 & n871;
  assign n873 = inC6 & musel2;
  assign n874 = inA6 & ~musel2;
  assign n875 = musel1 & n874;
  assign n876 = ~musel1 & n873;
  assign n877 = ~n875 & ~n876;
  assign n878 = n97 & ~n877;
  assign n879 = n104 & ~n878;
  assign n880 = ~n104 & n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n872 & ~n881;
  assign n883 = n872 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = opsel2 & ~n884;
  assign n886 = n112 & n885;
  assign n887 = inD14 & musel2;
  assign n888 = ~inB14 & ~n887;
  assign n889 = ~inB14 & ~musel1;
  assign n890 = n118 & ~n887;
  assign n891 = ~n122 & ~n890;
  assign n892 = ~n889 & n891;
  assign n893 = ~n888 & n892;
  assign n894 = inD14 & musel4;
  assign n895 = ~musel3 & n894;
  assign n896 = n126 & n895;
  assign n897 = n114 & n893;
  assign n898 = ~n896 & ~n897;
  assign n899 = sh2 & ~n898;
  assign n900 = ~n803 & ~n899;
  assign n901 = n802 & n900;
  assign n902 = sh1 & n900;
  assign n903 = ~n806 & ~n902;
  assign n904 = ~n901 & n903;
  assign n905 = ~n560 & ~n674;
  assign n906 = ~sh2 & ~n321;
  assign n907 = ~n340 & ~n906;
  assign n908 = n905 & n907;
  assign n909 = ~sh1 & n905;
  assign n910 = sh1 & n907;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n908 & n911;
  assign n913 = ~sh0 & n904;
  assign n914 = sh0 & n912;
  assign n915 = ~n913 & ~n914;
  assign n916 = n884 & n915;
  assign n917 = ~opsel2 & n884;
  assign n918 = opsel2 & n915;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n916 & n919;
  assign n921 = ~n886 & ~n920;
  assign n922 = n112 & ~n886;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~inA6 & ~n873;
  assign n925 = ~inA6 & ~musel1;
  assign n926 = n118 & ~n873;
  assign n927 = ~n122 & ~n926;
  assign n928 = ~n925 & n927;
  assign n929 = ~n924 & n928;
  assign n930 = n114 & n929;
  assign n931 = inC6 & musel4;
  assign n932 = ~musel3 & n931;
  assign n933 = ~musel2 & n932;
  assign n934 = ~musel1 & n933;
  assign n935 = ~n930 & ~n934;
  assign n936 = ~n244 & ~n935;
  assign n937 = n244 & n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = inB6 & ~musel3;
  assign n940 = musel2 & n939;
  assign n941 = inD6 & musel3;
  assign n942 = ~musel2 & n941;
  assign n943 = ~musel1 & n940;
  assign n944 = ~musel1 & n942;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~inA6 & ~musel2;
  assign n947 = ~inC6 & musel2;
  assign n948 = ~inA6 & ~inC6;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~n946 & n949;
  assign n951 = n272 & n950;
  assign n952 = n945 & ~n951;
  assign n953 = ~musel4 & ~n952;
  assign n954 = n938 & n953;
  assign n955 = ~n938 & ~n953;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n855 & ~n856;
  assign n958 = n835 & ~n850;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n835 & n850;
  assign n961 = n956 & n959;
  assign n962 = n956 & n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n861 & ~n960;
  assign n965 = ~n958 & ~n964;
  assign n966 = n956 & n963;
  assign n967 = n963 & n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = n238 & n968;
  assign n970 = n112 & ~n915;
  assign n971 = ~n969 & ~n970;
  assign n972 = n281 & ~n971;
  assign n973 = ~opsel3 & n923;
  assign O6 = n972 | n973;
  assign n975 = ~n778 & ~n881;
  assign n976 = ~n649 & n975;
  assign n977 = n640 & n976;
  assign n978 = inC7 & musel2;
  assign n979 = inA7 & ~musel2;
  assign n980 = musel1 & n979;
  assign n981 = ~musel1 & n978;
  assign n982 = ~n980 & ~n981;
  assign n983 = n97 & ~n982;
  assign n984 = n104 & ~n983;
  assign n985 = ~n104 & n983;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n977 & ~n986;
  assign n988 = n977 & n986;
  assign n989 = ~n987 & ~n988;
  assign n990 = opsel2 & ~n989;
  assign n991 = n112 & n990;
  assign n992 = inD15 & musel2;
  assign n993 = ~inB15 & ~n992;
  assign n994 = ~inB15 & ~musel1;
  assign n995 = n118 & ~n992;
  assign n996 = ~n122 & ~n995;
  assign n997 = ~n994 & n996;
  assign n998 = ~n993 & n997;
  assign n999 = inD15 & musel4;
  assign n1000 = ~musel3 & n999;
  assign n1001 = n126 & n1000;
  assign n1002 = n114 & n998;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = sh2 & ~n1003;
  assign n1005 = ~n906 & ~n1004;
  assign n1006 = n905 & n1005;
  assign n1007 = sh1 & n1005;
  assign n1008 = ~n909 & ~n1007;
  assign n1009 = ~n1006 & n1008;
  assign n1010 = ~n667 & ~n803;
  assign n1011 = ~sh2 & ~n438;
  assign n1012 = ~n457 & ~n1011;
  assign n1013 = n1010 & n1012;
  assign n1014 = ~sh1 & n1010;
  assign n1015 = sh1 & n1012;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n1013 & n1016;
  assign n1018 = ~sh0 & n1009;
  assign n1019 = sh0 & n1017;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = n989 & n1020;
  assign n1022 = ~opsel2 & n989;
  assign n1023 = opsel2 & n1020;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n1021 & n1024;
  assign n1026 = ~n991 & ~n1025;
  assign n1027 = n112 & ~n991;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~inA7 & ~n978;
  assign n1030 = ~inA7 & ~musel1;
  assign n1031 = n118 & ~n978;
  assign n1032 = ~n122 & ~n1031;
  assign n1033 = ~n1030 & n1032;
  assign n1034 = ~n1029 & n1033;
  assign n1035 = n114 & n1034;
  assign n1036 = inC7 & musel4;
  assign n1037 = ~musel3 & n1036;
  assign n1038 = ~musel2 & n1037;
  assign n1039 = ~musel1 & n1038;
  assign n1040 = ~n1035 & ~n1039;
  assign n1041 = ~n244 & ~n1040;
  assign n1042 = n244 & n1040;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = inB7 & ~musel3;
  assign n1045 = musel2 & n1044;
  assign n1046 = inD7 & musel3;
  assign n1047 = ~musel2 & n1046;
  assign n1048 = ~musel1 & n1045;
  assign n1049 = ~musel1 & n1047;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = ~inA7 & ~musel2;
  assign n1052 = ~inC7 & musel2;
  assign n1053 = ~inA7 & ~inC7;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = ~n1051 & n1054;
  assign n1056 = n272 & n1055;
  assign n1057 = n1050 & ~n1056;
  assign n1058 = ~musel4 & ~n1057;
  assign n1059 = n1043 & n1058;
  assign n1060 = ~n1043 & ~n1058;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n854 & ~n856;
  assign n1063 = ~n860 & ~n1062;
  assign n1064 = ~n958 & n1063;
  assign n1065 = ~n960 & ~n1064;
  assign n1066 = n938 & ~n953;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~n938 & n953;
  assign n1069 = n1061 & n1067;
  assign n1070 = n1061 & n1068;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = n861 & ~n958;
  assign n1073 = ~n958 & n960;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n1068 & n1074;
  assign n1076 = ~n1066 & ~n1075;
  assign n1077 = n1071 & n1076;
  assign n1078 = n1061 & n1071;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = n238 & n1079;
  assign n1081 = n112 & ~n1020;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n281 & ~n1082;
  assign n1084 = ~opsel3 & n1028;
  assign O7 = n1083 | n1084;
  assign n1086 = inC8 & musel2;
  assign n1087 = inA8 & ~musel2;
  assign n1088 = musel1 & n1087;
  assign n1089 = ~musel1 & n1086;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n97 & ~n1090;
  assign n1092 = n104 & ~n1091;
  assign n1093 = ~n104 & n1091;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = inC9 & musel2;
  assign n1096 = inA9 & ~musel2;
  assign n1097 = musel1 & n1096;
  assign n1098 = ~musel1 & n1095;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = n97 & ~n1099;
  assign n1101 = n104 & ~n1100;
  assign n1102 = ~n104 & n1100;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = inC10 & musel2;
  assign n1105 = inA10 & ~musel2;
  assign n1106 = musel1 & n1105;
  assign n1107 = ~musel1 & n1104;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = n97 & ~n1108;
  assign n1110 = n104 & ~n1109;
  assign n1111 = ~n104 & n1109;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = inC11 & musel2;
  assign n1114 = inA11 & ~musel2;
  assign n1115 = musel1 & n1114;
  assign n1116 = ~musel1 & n1113;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = n97 & ~n1117;
  assign n1119 = n104 & ~n1118;
  assign n1120 = ~n104 & n1118;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n1112 & ~n1121;
  assign n1123 = ~n1103 & n1122;
  assign n1124 = ~n1094 & n1123;
  assign n1125 = n639 & n1124;
  assign n1126 = n104 & n1125;
  assign n1127 = n1094 & n1126;
  assign n1128 = ~n1094 & ~n1126;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = opsel2 & ~n1129;
  assign n1131 = n112 & n1130;
  assign n1132 = ~n1004 & ~n1011;
  assign n1133 = n1010 & n1132;
  assign n1134 = sh1 & n1132;
  assign n1135 = ~n1014 & ~n1134;
  assign n1136 = ~n1133 & n1135;
  assign n1137 = ~n796 & ~n906;
  assign n1138 = ~sh2 & ~n559;
  assign n1139 = ~n171 & ~n1138;
  assign n1140 = n1137 & n1139;
  assign n1141 = ~sh1 & n1137;
  assign n1142 = sh1 & n1139;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n1140 & n1143;
  assign n1145 = ~sh0 & n1136;
  assign n1146 = sh0 & n1144;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = n1129 & n1147;
  assign n1149 = ~opsel2 & n1129;
  assign n1150 = opsel2 & n1147;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1148 & n1151;
  assign n1153 = ~n1131 & ~n1152;
  assign n1154 = n112 & ~n1131;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = ~inA8 & ~n1086;
  assign n1157 = ~inA8 & ~musel1;
  assign n1158 = n118 & ~n1086;
  assign n1159 = ~n122 & ~n1158;
  assign n1160 = ~n1157 & n1159;
  assign n1161 = ~n1156 & n1160;
  assign n1162 = n114 & n1161;
  assign n1163 = inC8 & musel4;
  assign n1164 = ~musel3 & n1163;
  assign n1165 = ~musel2 & n1164;
  assign n1166 = ~musel1 & n1165;
  assign n1167 = ~n1162 & ~n1166;
  assign n1168 = ~n244 & ~n1167;
  assign n1169 = n244 & n1167;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = inB8 & ~musel3;
  assign n1172 = musel2 & n1171;
  assign n1173 = inD8 & musel3;
  assign n1174 = ~musel2 & n1173;
  assign n1175 = ~musel1 & n1172;
  assign n1176 = ~musel1 & n1174;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = ~inA8 & ~musel2;
  assign n1179 = ~inC8 & musel2;
  assign n1180 = ~inA8 & ~inC8;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1178 & n1181;
  assign n1183 = n272 & n1182;
  assign n1184 = n1177 & ~n1183;
  assign n1185 = ~musel4 & ~n1184;
  assign n1186 = n1170 & n1185;
  assign n1187 = ~n1170 & ~n1185;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n709 & ~n835;
  assign n1190 = ~n709 & n850;
  assign n1191 = n724 & n850;
  assign n1192 = n724 & ~n835;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1190 & n1193;
  assign n1195 = ~n1189 & n1194;
  assign n1196 = ~n938 & ~n1043;
  assign n1197 = ~n938 & n1058;
  assign n1198 = n953 & n1058;
  assign n1199 = n953 & ~n1043;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1197 & n1200;
  assign n1202 = ~n1196 & n1201;
  assign n1203 = ~n1195 & ~n1202;
  assign n1204 = ~n856 & ~n960;
  assign n1205 = n958 & ~n960;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n938 & n1206;
  assign n1208 = n953 & n1206;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n1043 & ~n1058;
  assign n1211 = ~n1068 & n1209;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = ~n1043 & n1058;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n755 & n1203;
  assign n1216 = n1214 & ~n1215;
  assign n1217 = n1188 & ~n1216;
  assign n1218 = ~n1188 & n1216;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = n694 & n1147;
  assign n1221 = n1147 & n1219;
  assign n1222 = ~n112 & n1219;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1220 & n1223;
  assign n1225 = ~n759 & n1224;
  assign n1226 = ~opsel3 & n1155;
  assign n1227 = n281 & n1225;
  assign O8 = n1226 | n1227;
  assign n1229 = ~n1094 & n1126;
  assign n1230 = ~n1103 & ~n1229;
  assign n1231 = n1103 & n1229;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = opsel2 & ~n1232;
  assign n1234 = n112 & n1233;
  assign n1235 = ~n1004 & ~n1138;
  assign n1236 = n1137 & n1235;
  assign n1237 = sh1 & n1235;
  assign n1238 = ~n1141 & ~n1237;
  assign n1239 = ~n1236 & n1238;
  assign n1240 = ~n899 & ~n1011;
  assign n1241 = ~sh2 & ~n666;
  assign n1242 = ~n322 & ~n1241;
  assign n1243 = n1240 & n1242;
  assign n1244 = ~sh1 & n1240;
  assign n1245 = sh1 & n1242;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~n1243 & n1246;
  assign n1248 = ~sh0 & n1239;
  assign n1249 = sh0 & n1247;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = n1232 & n1250;
  assign n1252 = ~opsel2 & n1232;
  assign n1253 = opsel2 & n1250;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1251 & n1254;
  assign n1256 = ~n1234 & ~n1255;
  assign n1257 = n112 & ~n1234;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~inA9 & ~n1095;
  assign n1260 = ~inA9 & ~musel1;
  assign n1261 = n118 & ~n1095;
  assign n1262 = ~n122 & ~n1261;
  assign n1263 = ~n1260 & n1262;
  assign n1264 = ~n1259 & n1263;
  assign n1265 = n114 & n1264;
  assign n1266 = inC9 & musel4;
  assign n1267 = ~musel3 & n1266;
  assign n1268 = ~musel2 & n1267;
  assign n1269 = ~musel1 & n1268;
  assign n1270 = ~n1265 & ~n1269;
  assign n1271 = ~n244 & ~n1270;
  assign n1272 = n244 & n1270;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = inB9 & ~musel3;
  assign n1275 = musel2 & n1274;
  assign n1276 = inD9 & musel3;
  assign n1277 = ~musel2 & n1276;
  assign n1278 = ~musel1 & n1275;
  assign n1279 = ~musel1 & n1277;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~inA9 & ~musel2;
  assign n1282 = ~inC9 & musel2;
  assign n1283 = ~inA9 & ~inC9;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = ~n1281 & n1284;
  assign n1286 = n272 & n1285;
  assign n1287 = n1280 & ~n1286;
  assign n1288 = ~musel4 & ~n1287;
  assign n1289 = n1273 & n1288;
  assign n1290 = ~n1273 & ~n1288;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = n1170 & ~n1185;
  assign n1293 = ~n1216 & ~n1292;
  assign n1294 = ~n1170 & n1185;
  assign n1295 = n1291 & n1293;
  assign n1296 = n1291 & n1294;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n1216 & ~n1294;
  assign n1299 = ~n1292 & ~n1298;
  assign n1300 = n1291 & n1297;
  assign n1301 = n1297 & n1299;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = n238 & n1302;
  assign n1304 = n112 & ~n1250;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n281 & ~n1305;
  assign n1307 = ~opsel3 & n1258;
  assign O9 = n1306 | n1307;
  assign n1309 = ~n1094 & ~n1103;
  assign n1310 = n1126 & n1309;
  assign n1311 = ~n1112 & ~n1310;
  assign n1312 = n1112 & n1310;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = opsel2 & ~n1313;
  assign n1315 = n112 & n1314;
  assign n1316 = ~n1004 & ~n1241;
  assign n1317 = n1240 & n1316;
  assign n1318 = sh1 & n1316;
  assign n1319 = ~n1244 & ~n1318;
  assign n1320 = ~n1317 & n1319;
  assign n1321 = ~sh2 & ~n795;
  assign n1322 = ~n439 & ~n1321;
  assign n1323 = n1235 & n1322;
  assign n1324 = ~sh1 & n1235;
  assign n1325 = sh1 & n1322;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = ~n1323 & n1326;
  assign n1328 = ~sh0 & n1320;
  assign n1329 = sh0 & n1327;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = n1313 & n1330;
  assign n1332 = ~opsel2 & n1313;
  assign n1333 = opsel2 & n1330;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1331 & n1334;
  assign n1336 = ~n1315 & ~n1335;
  assign n1337 = n112 & ~n1315;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~inA10 & ~n1104;
  assign n1340 = ~inA10 & ~musel1;
  assign n1341 = n118 & ~n1104;
  assign n1342 = ~n122 & ~n1341;
  assign n1343 = ~n1340 & n1342;
  assign n1344 = ~n1339 & n1343;
  assign n1345 = n114 & n1344;
  assign n1346 = inC10 & musel4;
  assign n1347 = ~musel3 & n1346;
  assign n1348 = ~musel2 & n1347;
  assign n1349 = ~musel1 & n1348;
  assign n1350 = ~n1345 & ~n1349;
  assign n1351 = ~n244 & ~n1350;
  assign n1352 = n244 & n1350;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = inB10 & ~musel3;
  assign n1355 = musel2 & n1354;
  assign n1356 = inD10 & musel3;
  assign n1357 = ~musel2 & n1356;
  assign n1358 = ~musel1 & n1355;
  assign n1359 = ~musel1 & n1357;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~inA10 & ~musel2;
  assign n1362 = ~inC10 & musel2;
  assign n1363 = ~inA10 & ~inC10;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1361 & n1364;
  assign n1366 = n272 & n1365;
  assign n1367 = n1360 & ~n1366;
  assign n1368 = ~musel4 & ~n1367;
  assign n1369 = n1353 & n1368;
  assign n1370 = ~n1353 & ~n1368;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1293 & ~n1294;
  assign n1373 = n1273 & ~n1288;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1273 & n1288;
  assign n1376 = n1371 & n1374;
  assign n1377 = n1371 & n1375;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1299 & ~n1375;
  assign n1380 = ~n1373 & ~n1379;
  assign n1381 = n1371 & n1378;
  assign n1382 = n1378 & n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = n238 & n1383;
  assign n1385 = n112 & ~n1330;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = n281 & ~n1386;
  assign n1388 = ~opsel3 & n1338;
  assign O10 = n1387 | n1388;
  assign n1390 = ~n1103 & ~n1112;
  assign n1391 = ~n1094 & n1390;
  assign n1392 = n1126 & n1391;
  assign n1393 = ~n1121 & ~n1392;
  assign n1394 = n1121 & n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = opsel2 & ~n1395;
  assign n1397 = n112 & n1396;
  assign n1398 = sh0 & sh1;
  assign n1399 = ~sh2 & ~n898;
  assign n1400 = ~sh2 & ~n1399;
  assign n1401 = n559 & ~n1399;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = sh1 & ~n795;
  assign n1404 = n559 & ~n1403;
  assign n1405 = sh1 & ~n1403;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = sh0 & ~sh1;
  assign n1408 = ~sh0 & n1406;
  assign n1409 = ~n666 & n1407;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1004 & n1410;
  assign n1412 = n1398 & n1410;
  assign n1413 = sh2 & n1398;
  assign n1414 = sh2 & ~n1004;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~n1412 & n1415;
  assign n1417 = ~n1411 & n1416;
  assign n1418 = n1398 & n1402;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1395 & n1419;
  assign n1421 = ~opsel2 & n1395;
  assign n1422 = opsel2 & n1419;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~n1420 & n1423;
  assign n1425 = ~n1397 & ~n1424;
  assign n1426 = n112 & ~n1397;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~inA11 & ~n1113;
  assign n1429 = ~inA11 & ~musel1;
  assign n1430 = n118 & ~n1113;
  assign n1431 = ~n122 & ~n1430;
  assign n1432 = ~n1429 & n1431;
  assign n1433 = ~n1428 & n1432;
  assign n1434 = n114 & n1433;
  assign n1435 = inC11 & musel4;
  assign n1436 = ~musel3 & n1435;
  assign n1437 = ~musel2 & n1436;
  assign n1438 = ~musel1 & n1437;
  assign n1439 = ~n1434 & ~n1438;
  assign n1440 = ~n244 & ~n1439;
  assign n1441 = n244 & n1439;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = inB11 & ~musel3;
  assign n1444 = musel2 & n1443;
  assign n1445 = inD11 & musel3;
  assign n1446 = ~musel2 & n1445;
  assign n1447 = ~musel1 & n1444;
  assign n1448 = ~musel1 & n1446;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~inA11 & ~musel2;
  assign n1451 = ~inC11 & musel2;
  assign n1452 = ~inA11 & ~inC11;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~n1450 & n1453;
  assign n1455 = n272 & n1454;
  assign n1456 = n1449 & ~n1455;
  assign n1457 = ~musel4 & ~n1456;
  assign n1458 = n1442 & n1457;
  assign n1459 = ~n1442 & ~n1457;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = n1292 & ~n1294;
  assign n1462 = ~n1298 & ~n1461;
  assign n1463 = ~n1373 & n1462;
  assign n1464 = ~n1375 & ~n1463;
  assign n1465 = n1353 & ~n1368;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1353 & n1368;
  assign n1468 = n1460 & n1466;
  assign n1469 = n1460 & n1467;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n1299 & ~n1373;
  assign n1472 = ~n1373 & n1375;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = ~n1467 & n1473;
  assign n1475 = ~n1465 & ~n1474;
  assign n1476 = n1470 & n1475;
  assign n1477 = n1460 & n1470;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = n238 & n1478;
  assign n1480 = n112 & ~n1419;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = n281 & ~n1481;
  assign n1483 = ~opsel3 & n1427;
  assign O11 = n1482 | n1483;
  assign n1485 = ~n881 & ~n986;
  assign n1486 = ~n778 & n1485;
  assign n1487 = ~n649 & n1486;
  assign n1488 = n1124 & n1487;
  assign n1489 = n104 & n1488;
  assign n1490 = n639 & n1489;
  assign n1491 = inC12 & musel2;
  assign n1492 = inA12 & ~musel2;
  assign n1493 = musel1 & n1492;
  assign n1494 = ~musel1 & n1491;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = n97 & ~n1495;
  assign n1497 = n104 & ~n1496;
  assign n1498 = ~n104 & n1496;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1490 & ~n1499;
  assign n1501 = n1490 & n1499;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = opsel2 & ~n1502;
  assign n1504 = n112 & n1503;
  assign n1505 = ~n795 & n1407;
  assign n1506 = ~n1003 & n1398;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = sh1 & ~n898;
  assign n1509 = ~sh1 & ~n666;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = n1507 & n1510;
  assign n1512 = sh0 & n1507;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = n666 & n1398;
  assign n1515 = n1003 & ~n1398;
  assign n1516 = n666 & n1003;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1514 & n1517;
  assign n1519 = ~sh2 & n1513;
  assign n1520 = sh2 & n1518;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = n1502 & n1521;
  assign n1523 = ~opsel2 & n1502;
  assign n1524 = opsel2 & n1521;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1522 & n1525;
  assign n1527 = ~n1504 & ~n1526;
  assign n1528 = n112 & ~n1504;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = inB12 & ~musel3;
  assign n1531 = musel2 & n1530;
  assign n1532 = inD12 & musel3;
  assign n1533 = ~musel2 & n1532;
  assign n1534 = ~musel1 & n1531;
  assign n1535 = ~musel1 & n1533;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~inA12 & ~musel2;
  assign n1538 = ~inC12 & musel2;
  assign n1539 = ~inA12 & ~inC12;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1537 & n1540;
  assign n1542 = n272 & n1541;
  assign n1543 = n1536 & ~n1542;
  assign n1544 = ~musel4 & ~n1543;
  assign n1545 = ~inA12 & ~n1491;
  assign n1546 = ~inA12 & ~musel1;
  assign n1547 = n118 & ~n1491;
  assign n1548 = ~n122 & ~n1547;
  assign n1549 = ~n1546 & n1548;
  assign n1550 = ~n1545 & n1549;
  assign n1551 = n114 & n1550;
  assign n1552 = inC12 & musel4;
  assign n1553 = ~musel3 & n1552;
  assign n1554 = ~musel2 & n1553;
  assign n1555 = ~musel1 & n1554;
  assign n1556 = ~n1551 & ~n1555;
  assign n1557 = ~n244 & ~n1556;
  assign n1558 = n244 & n1556;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = n1544 & n1559;
  assign n1561 = ~n1544 & ~n1559;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = ~n1273 & n1294;
  assign n1564 = n1288 & n1294;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1375 & n1565;
  assign n1567 = ~n1465 & ~n1566;
  assign n1568 = ~n1467 & ~n1567;
  assign n1569 = n1442 & ~n1457;
  assign n1570 = n1442 & n1568;
  assign n1571 = ~n1457 & n1568;
  assign n1572 = n1442 & n1569;
  assign n1573 = ~n1457 & n1569;
  assign n1574 = ~n1572 & ~n1573;
  assign n1575 = ~n1571 & n1574;
  assign n1576 = ~n1570 & n1575;
  assign n1577 = ~n1170 & ~n1273;
  assign n1578 = ~n1170 & n1288;
  assign n1579 = n1185 & n1288;
  assign n1580 = n1185 & ~n1273;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1578 & n1581;
  assign n1583 = ~n1577 & n1582;
  assign n1584 = ~n1353 & ~n1442;
  assign n1585 = ~n1353 & n1457;
  assign n1586 = n1368 & n1457;
  assign n1587 = n1368 & ~n1442;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n1585 & n1588;
  assign n1590 = ~n1584 & n1589;
  assign n1591 = ~n1216 & ~n1590;
  assign n1592 = ~n1583 & n1591;
  assign n1593 = ~n1576 & ~n1592;
  assign n1594 = n1562 & ~n1593;
  assign n1595 = ~n1562 & n1593;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = n694 & n1521;
  assign n1598 = n1521 & n1596;
  assign n1599 = ~n112 & n1596;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = ~n1597 & n1600;
  assign n1602 = ~n759 & n1601;
  assign n1603 = ~opsel3 & n1529;
  assign n1604 = n281 & n1602;
  assign O12 = n1603 | n1604;
  assign n1606 = n1490 & ~n1499;
  assign n1607 = inC13 & musel2;
  assign n1608 = inA13 & ~musel2;
  assign n1609 = musel1 & n1608;
  assign n1610 = ~musel1 & n1607;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = n97 & ~n1611;
  assign n1613 = n104 & ~n1612;
  assign n1614 = ~n104 & n1612;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1606 & ~n1615;
  assign n1617 = n1606 & n1615;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = opsel2 & ~n1618;
  assign n1620 = n112 & n1619;
  assign n1621 = sh0 & sh2;
  assign n1622 = ~sh1 & ~sh2;
  assign n1623 = sh1 & ~n1621;
  assign n1624 = ~sh1 & sh2;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = sh0 & ~n898;
  assign n1627 = ~sh0 & ~n795;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = ~n1622 & n1625;
  assign n1630 = n1003 & ~n1622;
  assign n1631 = n1625 & n1628;
  assign n1632 = n1003 & n1628;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n1630 & n1633;
  assign n1635 = ~n1629 & n1634;
  assign n1636 = n1403 & n1621;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n1618 & n1637;
  assign n1639 = ~opsel2 & n1618;
  assign n1640 = opsel2 & n1637;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~n1638 & n1641;
  assign n1643 = ~n1620 & ~n1642;
  assign n1644 = n112 & ~n1620;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = inB13 & ~musel3;
  assign n1647 = musel2 & n1646;
  assign n1648 = inD13 & musel3;
  assign n1649 = ~musel2 & n1648;
  assign n1650 = ~musel1 & n1647;
  assign n1651 = ~musel1 & n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = ~inA13 & ~musel2;
  assign n1654 = ~inC13 & musel2;
  assign n1655 = ~inA13 & ~inC13;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1653 & n1656;
  assign n1658 = n272 & n1657;
  assign n1659 = n1652 & ~n1658;
  assign n1660 = ~musel4 & ~n1659;
  assign n1661 = ~inA13 & ~n1607;
  assign n1662 = ~inA13 & ~musel1;
  assign n1663 = n118 & ~n1607;
  assign n1664 = ~n122 & ~n1663;
  assign n1665 = ~n1662 & n1664;
  assign n1666 = ~n1661 & n1665;
  assign n1667 = n114 & n1666;
  assign n1668 = inC13 & musel4;
  assign n1669 = ~musel3 & n1668;
  assign n1670 = ~musel2 & n1669;
  assign n1671 = ~musel1 & n1670;
  assign n1672 = ~n1667 & ~n1671;
  assign n1673 = ~n244 & ~n1672;
  assign n1674 = n244 & n1672;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = n1660 & n1675;
  assign n1677 = ~n1660 & ~n1675;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1544 & n1559;
  assign n1680 = ~n1593 & ~n1679;
  assign n1681 = n1544 & ~n1559;
  assign n1682 = n1678 & n1680;
  assign n1683 = n1678 & n1681;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = n1593 & ~n1681;
  assign n1686 = ~n1679 & ~n1685;
  assign n1687 = n1678 & n1684;
  assign n1688 = n1684 & n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = n238 & n1689;
  assign n1691 = n112 & ~n1637;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = n281 & ~n1692;
  assign n1694 = ~opsel3 & n1645;
  assign O13 = n1693 | n1694;
  assign n1696 = n1490 & ~n1615;
  assign n1697 = ~n1499 & n1696;
  assign n1698 = inC14 & musel2;
  assign n1699 = inA14 & ~musel2;
  assign n1700 = musel1 & n1699;
  assign n1701 = ~musel1 & n1698;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = n97 & ~n1702;
  assign n1704 = n104 & ~n1703;
  assign n1705 = ~n104 & n1703;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1697 & ~n1706;
  assign n1708 = n1697 & n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = opsel2 & ~n1709;
  assign n1711 = n112 & n1710;
  assign n1712 = ~sh0 & ~sh2;
  assign n1713 = sh1 & ~sh2;
  assign n1714 = ~n1398 & ~n1713;
  assign n1715 = ~n1712 & n1714;
  assign n1716 = ~n1713 & ~n1715;
  assign n1717 = ~n1003 & ~n1716;
  assign n1718 = ~n898 & n1716;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = n1709 & n1719;
  assign n1721 = ~opsel2 & n1709;
  assign n1722 = opsel2 & n1719;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = ~n1720 & n1723;
  assign n1725 = ~n1711 & ~n1724;
  assign n1726 = n112 & ~n1711;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = inB14 & ~musel3;
  assign n1729 = musel2 & n1728;
  assign n1730 = inD14 & musel3;
  assign n1731 = ~musel2 & n1730;
  assign n1732 = ~musel1 & n1729;
  assign n1733 = ~musel1 & n1731;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~inA14 & ~musel2;
  assign n1736 = ~inC14 & musel2;
  assign n1737 = ~inA14 & ~inC14;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = n272 & n1739;
  assign n1741 = n1734 & ~n1740;
  assign n1742 = ~musel4 & ~n1741;
  assign n1743 = ~inA14 & ~n1698;
  assign n1744 = ~inA14 & ~musel1;
  assign n1745 = n118 & ~n1698;
  assign n1746 = ~n122 & ~n1745;
  assign n1747 = ~n1744 & n1746;
  assign n1748 = ~n1743 & n1747;
  assign n1749 = n114 & n1748;
  assign n1750 = inC14 & musel4;
  assign n1751 = ~musel3 & n1750;
  assign n1752 = ~musel2 & n1751;
  assign n1753 = ~musel1 & n1752;
  assign n1754 = ~n1749 & ~n1753;
  assign n1755 = ~n244 & ~n1754;
  assign n1756 = n244 & n1754;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = n1742 & n1757;
  assign n1759 = ~n1742 & ~n1757;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = ~n1680 & ~n1681;
  assign n1762 = ~n1660 & n1675;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = n1660 & ~n1675;
  assign n1765 = n1760 & n1763;
  assign n1766 = n1760 & n1764;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = ~n1686 & ~n1764;
  assign n1769 = ~n1762 & ~n1768;
  assign n1770 = n1760 & n1767;
  assign n1771 = n1767 & n1769;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = n238 & n1772;
  assign n1774 = n112 & ~n1719;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = n281 & ~n1775;
  assign n1777 = ~opsel3 & n1727;
  assign O14 = n1776 | n1777;
  assign n1779 = ~n1615 & ~n1706;
  assign n1780 = ~n1499 & n1779;
  assign n1781 = n1490 & n1780;
  assign n1782 = opsel2 & n112;
  assign n1783 = n1781 & n1782;
  assign n1784 = opsel2 & ~n1003;
  assign n1785 = ~opsel2 & n1781;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1783 & n1786;
  assign n1788 = n112 & ~n1783;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~inA15 & ~n99;
  assign n1791 = ~inA15 & ~musel1;
  assign n1792 = ~n99 & n118;
  assign n1793 = ~n122 & ~n1792;
  assign n1794 = ~n1791 & n1793;
  assign n1795 = ~n1790 & n1794;
  assign n1796 = n114 & n1795;
  assign n1797 = inC15 & musel4;
  assign n1798 = ~musel3 & n1797;
  assign n1799 = ~musel2 & n1798;
  assign n1800 = ~musel1 & n1799;
  assign n1801 = ~n1796 & ~n1800;
  assign n1802 = ~n244 & ~n1801;
  assign n1803 = n244 & n1801;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = inB15 & ~musel3;
  assign n1806 = musel2 & n1805;
  assign n1807 = inD15 & musel3;
  assign n1808 = ~musel2 & n1807;
  assign n1809 = ~musel1 & n1806;
  assign n1810 = ~musel1 & n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~inA15 & ~musel2;
  assign n1813 = ~inC15 & musel2;
  assign n1814 = ~inA15 & ~inC15;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1812 & n1815;
  assign n1817 = n272 & n1816;
  assign n1818 = n1811 & ~n1817;
  assign n1819 = ~musel4 & ~n1818;
  assign n1820 = ~n1804 & ~n1819;
  assign n1821 = n1804 & n1819;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = n1679 & ~n1681;
  assign n1824 = ~n1685 & ~n1823;
  assign n1825 = ~n1762 & n1824;
  assign n1826 = ~n1764 & ~n1825;
  assign n1827 = ~n1742 & n1757;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = n1742 & ~n1757;
  assign n1830 = n1822 & n1828;
  assign n1831 = n1822 & n1829;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1686 & ~n1762;
  assign n1834 = ~n1762 & n1764;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~n1829 & n1835;
  assign n1837 = ~n1827 & ~n1836;
  assign n1838 = n1832 & n1837;
  assign n1839 = n1822 & n1832;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = n238 & n1840;
  assign n1842 = n112 & ~n1003;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = n281 & ~n1843;
  assign n1845 = ~opsel3 & n1789;
  assign O15 = n1844 | n1845;
endmodule


