// Benchmark "frg2" written by ABC on Tue May 16 16:07:49 2017

module frg2 ( 
    z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r,
    s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4, c0, c1,
    c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2, f3, f4,
    g0, g1, g2, g3, g4, h0, h1, h2, h3, h4, i0, i1, i2, i3, i4, j0, j1, j2,
    j3, j4, k0, k1, k2, k3, k4, l0, l1, l2, l3, l4, m0, m1, m2, m3, m4, n0,
    n1, n2, n3, n4, o0, o1, o2, o3, p0, p1, p2, p3, q0, q1, q2, q3, r1, r2,
    r3, s0, s1, s2, s3, t0, t1, t2, t3, u0, u1, u2, u3, v0, v1, v2, v3, w0,
    w1, w2, w3, x0, x1, x2, x3, y0, y1, y2, y3,
    z4, z5, z6, z7, z8, a5, a6, a7, a8, a9, b5, b6, b7, b8, b9, c5, c6, c7,
    c8, c9, d5, d6, d7, d8, d9, e5, e6, e7, e8, e9, f5, f6, f7, f8, f9, g5,
    g6, g7, g8, g9, h5, h6, h7, h8, h9, i5, i6, i7, i8, i9, j5, j6, j7, j8,
    j9, k5, k6, k7, k8, k9, l5, l6, l7, l8, l9, m5, m6, m7, m8, m9, n5, n6,
    n7, n8, n9, o4, o5, o6, o7, o8, o9, p4, p5, p6, p7, p8, p9, q4, q5, q6,
    q7, q8, q9, r4, r5, r6, r7, r8, r9, s4, s5, s6, s7, s8, s9, t4, t5, t6,
    t7, t8, t9, u4, u5, u6, u7, u8, u9, v4, v5, v6, v7, v8, v9, w4, w5, w6,
    w7, w8, w9, x4, x5, x6, x7, x8, y4, y5, y6, y7, y8  );
  input  z0, z1, z2, z3, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p,
    q, r, s, t, u, v, w, x, y, z, a0, a1, a2, a3, a4, b0, b1, b2, b3, b4,
    c0, c1, c2, c3, c4, d0, d1, d2, d3, d4, e0, e1, e2, e3, e4, f0, f1, f2,
    f3, f4, g0, g1, g2, g3, g4, h0, h1, h2, h3, h4, i0, i1, i2, i3, i4, j0,
    j1, j2, j3, j4, k0, k1, k2, k3, k4, l0, l1, l2, l3, l4, m0, m1, m2, m3,
    m4, n0, n1, n2, n3, n4, o0, o1, o2, o3, p0, p1, p2, p3, q0, q1, q2, q3,
    r1, r2, r3, s0, s1, s2, s3, t0, t1, t2, t3, u0, u1, u2, u3, v0, v1, v2,
    v3, w0, w1, w2, w3, x0, x1, x2, x3, y0, y1, y2, y3;
  output z4, z5, z6, z7, z8, a5, a6, a7, a8, a9, b5, b6, b7, b8, b9, c5, c6,
    c7, c8, c9, d5, d6, d7, d8, d9, e5, e6, e7, e8, e9, f5, f6, f7, f8, f9,
    g5, g6, g7, g8, g9, h5, h6, h7, h8, h9, i5, i6, i7, i8, i9, j5, j6, j7,
    j8, j9, k5, k6, k7, k8, k9, l5, l6, l7, l8, l9, m5, m6, m7, m8, m9, n5,
    n6, n7, n8, n9, o4, o5, o6, o7, o8, o9, p4, p5, p6, p7, p8, p9, q4, q5,
    q6, q7, q8, q9, r4, r5, r6, r7, r8, r9, s4, s5, s6, s7, s8, s9, t4, t5,
    t6, t7, t8, t9, u4, u5, u6, u7, u8, u9, v4, v5, v6, v7, v8, v9, w4, w5,
    w6, w7, w8, w9, x4, x5, x6, x7, x8, y4, y5, y6, y7, y8;
  wire n283, n284, n285, n286, n288, n289, n291, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n356, n357, n358, n359,
    n360, n361, n362, n365, n366, n369, n370, n371, n372, n373, n374, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n386, n387, n390, n391,
    n394, n395, n396, n397, n398, n399, n401, n402, n403, n404, n405, n406,
    n407, n408, n410, n411, n414, n415, n418, n419, n420, n421, n422, n423,
    n425, n426, n427, n428, n430, n431, n435, n436, n437, n438, n439, n440,
    n442, n443, n444, n445, n447, n448, n452, n453, n454, n455, n456, n457,
    n459, n460, n461, n462, n464, n465, n469, n470, n471, n472, n473, n474,
    n476, n477, n478, n479, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n507, n508, n509, n510, n511, n512, n514, n515, n516,
    n517, n519, n520, n521, n522, n524, n525, n526, n527, n528, n529, n531,
    n532, n533, n534, n536, n537, n538, n539, n540, n541, n542, n543, n545,
    n546, n547, n548, n549, n550, n552, n553, n555, n556, n557, n558, n559,
    n560, n562, n563, n564, n565, n566, n567, n569, n570, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n588, n589, n590, n591, n592, n593, n595, n596, n598, n599, n600, n601,
    n602, n603, n604, n607, n608, n609, n610, n611, n612, n614, n615, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n629, n630,
    n631, n632, n633, n635, n636, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n649, n651, n652, n654, n655, n656, n657, n658, n659,
    n661, n662, n664, n665, n666, n667, n668, n672, n673, n674, n675, n676,
    n677, n679, n680, n682, n683, n684, n685, n687, n688, n689, n690, n691,
    n694, n695, n696, n698, n699, n700, n701, n702, n703, n705, n706, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n720, n721,
    n722, n723, n726, n727, n728, n729, n730, n732, n733, n734, n735, n736,
    n737, n739, n740, n742, n743, n744, n745, n746, n747, n748, n749, n751,
    n752, n753, n754, n757, n758, n759, n761, n762, n763, n764, n765, n766,
    n768, n769, n771, n772, n773, n774, n775, n776, n778, n779, n780, n781,
    n783, n784, n786, n787, n788, n790, n791, n792, n793, n794, n795, n797,
    n798, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n813, n814, n815, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n828, n829, n831, n833, n834, n835, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n847, n848, n851, n852, n854, n855, n856,
    n857, n859, n860, n861, n862, n863, n864, n865, n866, n867, n869, n870,
    n872, n873, n875, n876, n878, n879, n880, n881, n882, n883, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n895, n896, n898, n899, n902,
    n903, n904, n905, n906, n907, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n919, n920, n922, n923, n926, n927, n928, n929, n930, n931,
    n933, n934, n935, n936, n937, n938, n939, n940, n942, n943;
  assign n283 = k0 & ~l0;
  assign n284 = ~k0 & l0;
  assign n285 = ~n283 & ~n284;
  assign n286 = m0 & n285;
  assign h5 = m0 & q3;
  assign n288 = i3 & n286;
  assign n289 = ~n285 & h5;
  assign z4 = n288 | n289;
  assign n291 = ~k4 & m1;
  assign z5 = ~j1 | ~n291;
  assign n293 = o0 & ~q0;
  assign n294 = ~k1 & ~l1;
  assign n295 = ~j1 & n294;
  assign n296 = ~i1 & n295;
  assign n297 = ~h1 & n296;
  assign n298 = ~n0 & n297;
  assign n299 = n293 & ~n298;
  assign n300 = z3 & y3;
  assign n301 = ~a4 & ~b4;
  assign n302 = n300 & n301;
  assign n303 = ~c4 & n302;
  assign n304 = ~x3 & n303;
  assign n305 = l4 & ~n304;
  assign n306 = n293 & n298;
  assign n307 = q1 & ~n305;
  assign n308 = n299 & n307;
  assign n309 = r1 & n305;
  assign n310 = n299 & n309;
  assign n311 = g0 & n306;
  assign n312 = ~n310 & ~n311;
  assign z6 = n308 | ~n312;
  assign n314 = ~m0 & n298;
  assign n315 = k0 & ~n285;
  assign n316 = n314 & n315;
  assign n317 = n305 & ~n314;
  assign n318 = ~n305 & ~n314;
  assign n319 = n285 & n314;
  assign n320 = l0 & n314;
  assign n321 = ~n319 & ~n320;
  assign n322 = o & n293;
  assign n323 = n316 & n322;
  assign n324 = r2 & n293;
  assign n325 = n317 & n324;
  assign n326 = q2 & n293;
  assign n327 = n318 & n326;
  assign n328 = g & n293;
  assign n329 = ~n321 & n328;
  assign n330 = ~n327 & ~n329;
  assign n331 = ~n325 & n330;
  assign z7 = n323 | ~n331;
  assign n333 = f4 & ~g4;
  assign n334 = e4 & n333;
  assign n335 = ~h4 & n334;
  assign n336 = j1 & ~n294;
  assign n337 = h1 & ~n296;
  assign n338 = i1 & ~n295;
  assign n339 = k1 & l1;
  assign n340 = ~n297 & ~n335;
  assign n341 = ~n339 & n340;
  assign n342 = ~n338 & n341;
  assign n343 = ~n337 & n342;
  assign n344 = ~n336 & n343;
  assign n345 = i1 & ~y0;
  assign n346 = ~a1 & k1;
  assign n347 = h1 & ~x0;
  assign n348 = ~z0 & j1;
  assign n349 = ~b1 & l1;
  assign n350 = ~n347 & ~n348;
  assign n351 = ~n346 & n350;
  assign n352 = ~n345 & n351;
  assign n353 = ~n349 & n352;
  assign n354 = n293 & ~n353;
  assign w9 = k4 & n354;
  assign n356 = n344 & w9;
  assign n357 = k4 & ~n353;
  assign n358 = n293 & ~n344;
  assign n359 = n293 & ~n357;
  assign n360 = ~n358 & ~n359;
  assign n361 = r3 & n356;
  assign n362 = q3 & ~n360;
  assign z8 = n361 | n362;
  assign i5 = m0 & r3;
  assign n365 = j3 & n286;
  assign n366 = ~n285 & i5;
  assign a5 = n365 | n366;
  assign a6 = ~k1 | ~n291;
  assign n369 = r1 & ~n305;
  assign n370 = n299 & n369;
  assign n371 = s1 & n305;
  assign n372 = n299 & n371;
  assign n373 = f0 & n306;
  assign n374 = ~n372 & ~n373;
  assign a7 = n370 | ~n374;
  assign n376 = p & n293;
  assign n377 = n316 & n376;
  assign n378 = s2 & n293;
  assign n379 = n317 & n378;
  assign n380 = n318 & n324;
  assign n381 = h & n293;
  assign n382 = ~n321 & n381;
  assign n383 = ~n380 & ~n382;
  assign n384 = ~n379 & n383;
  assign a8 = n377 | ~n384;
  assign n386 = s3 & n356;
  assign n387 = r3 & ~n360;
  assign a9 = n386 | n387;
  assign j5 = m0 & s3;
  assign n390 = k3 & n286;
  assign n391 = ~n285 & j5;
  assign b5 = n390 | n391;
  assign b6 = ~l1 | ~n291;
  assign n394 = s1 & ~n305;
  assign n395 = n299 & n394;
  assign n396 = t1 & n305;
  assign n397 = n299 & n396;
  assign n398 = e0 & n306;
  assign n399 = ~n397 & ~n398;
  assign b7 = n395 | ~n399;
  assign n401 = n293 & ~n319;
  assign n402 = n305 & n401;
  assign n403 = ~n305 & n401;
  assign n404 = n293 & n319;
  assign n405 = t2 & n402;
  assign n406 = s2 & n403;
  assign n407 = i & n404;
  assign n408 = ~n406 & ~n407;
  assign b8 = n405 | ~n408;
  assign n410 = t3 & n356;
  assign n411 = s3 & ~n360;
  assign b9 = n410 | n411;
  assign k5 = m0 & t3;
  assign n414 = l3 & n286;
  assign n415 = ~n285 & k5;
  assign c5 = n414 | n415;
  assign c6 = ~h1 | ~l4;
  assign n418 = t1 & ~n305;
  assign n419 = n299 & n418;
  assign n420 = u1 & n305;
  assign n421 = n299 & n420;
  assign n422 = d0 & n306;
  assign n423 = ~n421 & ~n422;
  assign c7 = n419 | ~n423;
  assign n425 = u2 & n402;
  assign n426 = t2 & n403;
  assign n427 = j & n404;
  assign n428 = ~n426 & ~n427;
  assign c8 = n425 | ~n428;
  assign n430 = u3 & n356;
  assign n431 = t3 & ~n360;
  assign c9 = n430 | n431;
  assign d5 = m0 & m3;
  assign d6 = ~i1 | ~l4;
  assign n435 = n306 & ~n314;
  assign n436 = v1 & n293;
  assign n437 = n317 & n436;
  assign n438 = u1 & n293;
  assign n439 = n318 & n438;
  assign n440 = ~n435 & ~n439;
  assign d7 = n437 | ~n440;
  assign n442 = v2 & n402;
  assign n443 = u2 & n403;
  assign n444 = k & n404;
  assign n445 = ~n443 & ~n444;
  assign d8 = n442 | ~n445;
  assign n447 = v3 & n356;
  assign n448 = u3 & ~n360;
  assign d9 = n447 | n448;
  assign e5 = m0 & n3;
  assign e6 = ~j1 | ~l4;
  assign n452 = v1 & ~n305;
  assign n453 = n299 & n452;
  assign n454 = w1 & n305;
  assign n455 = n299 & n454;
  assign n456 = k0 & n306;
  assign n457 = ~n455 & ~n456;
  assign e7 = n453 | ~n457;
  assign n459 = w2 & n402;
  assign n460 = v2 & n403;
  assign n461 = l & n404;
  assign n462 = ~n460 & ~n461;
  assign e8 = n459 | ~n462;
  assign n464 = w3 & n356;
  assign n465 = v3 & ~n360;
  assign e9 = n464 | n465;
  assign f5 = m0 & o3;
  assign f6 = ~k1 | ~l4;
  assign n469 = w1 & ~n305;
  assign n470 = n299 & n469;
  assign n471 = x1 & n305;
  assign n472 = n299 & n471;
  assign n473 = l0 & n306;
  assign n474 = ~n472 & ~n473;
  assign f7 = n470 | ~n474;
  assign n476 = x2 & n402;
  assign n477 = w2 & n403;
  assign n478 = m & n404;
  assign n479 = ~n477 & ~n478;
  assign f8 = n476 | ~n479;
  assign n481 = ~j1 & v0;
  assign n482 = ~i1 & w0;
  assign n483 = ~j1 & n482;
  assign n484 = ~k1 & n483;
  assign n485 = l1 & n484;
  assign n486 = ~i1 & k1;
  assign n487 = ~l1 & n486;
  assign n488 = n481 & n487;
  assign n489 = ~i1 & u0;
  assign n490 = j1 & n489;
  assign n491 = n294 & n490;
  assign n492 = i1 & t0;
  assign n493 = n295 & n492;
  assign n494 = ~n491 & ~n493;
  assign n495 = ~n488 & n494;
  assign n496 = ~n485 & n495;
  assign n497 = ~h1 & n496;
  assign n498 = h1 & ~s0;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n337 & n499;
  assign n501 = w9 & n500;
  assign n502 = ~n335 & n501;
  assign n503 = w3 & ~n360;
  assign f9 = n502 | n503;
  assign g5 = m0 & p3;
  assign g6 = ~l1 | ~l4;
  assign n507 = x1 & ~n305;
  assign n508 = n299 & n507;
  assign n509 = y1 & n305;
  assign n510 = n299 & n509;
  assign n511 = q & n306;
  assign n512 = ~n510 & ~n511;
  assign g7 = n508 | ~n512;
  assign n514 = y2 & n402;
  assign n515 = x2 & n403;
  assign n516 = n & n404;
  assign n517 = ~n515 & ~n516;
  assign g8 = n514 | ~n517;
  assign n519 = x3 & ~n305;
  assign n520 = n299 & n519;
  assign n521 = ~x3 & n305;
  assign n522 = n299 & n521;
  assign g9 = n520 | n522;
  assign n524 = y1 & ~n305;
  assign n525 = n299 & n524;
  assign n526 = z1 & n305;
  assign n527 = n299 & n526;
  assign n528 = r & n306;
  assign n529 = ~n527 & ~n528;
  assign h7 = n525 | ~n529;
  assign n531 = z2 & n402;
  assign n532 = y2 & n403;
  assign n533 = o & n404;
  assign n534 = ~n532 & ~n533;
  assign h8 = n531 | ~n534;
  assign n536 = ~x3 & y3;
  assign n537 = ~n304 & n536;
  assign n538 = n305 & g9;
  assign n539 = ~n537 & n538;
  assign n540 = y3 & ~n537;
  assign n541 = ~n305 & n537;
  assign n542 = n299 & ~n541;
  assign n543 = ~n540 & n542;
  assign h9 = n539 | ~n543;
  assign n545 = z1 & ~n305;
  assign n546 = n299 & n545;
  assign n547 = a2 & n305;
  assign n548 = n299 & n547;
  assign n549 = s & n306;
  assign n550 = ~n548 & ~n549;
  assign i7 = n546 | ~n550;
  assign n552 = z2 & n403;
  assign n553 = p & n404;
  assign i8 = n552 | n553;
  assign n555 = n537 & ~h9;
  assign n556 = ~n300 & n555;
  assign n557 = n300 & ~n305;
  assign n558 = z3 & ~n537;
  assign n559 = n299 & ~n558;
  assign n560 = ~n557 & n559;
  assign i9 = n556 | ~n560;
  assign n562 = a2 & ~n305;
  assign n563 = n299 & n562;
  assign n564 = b2 & n305;
  assign n565 = n299 & n564;
  assign n566 = t & n306;
  assign n567 = ~n565 & ~n566;
  assign j7 = n563 | ~n567;
  assign n569 = b3 & n356;
  assign n570 = a3 & ~n360;
  assign j8 = n569 | n570;
  assign n572 = z3 & ~a4;
  assign n573 = n293 & n537;
  assign n574 = n317 & n573;
  assign n575 = n572 & n574;
  assign n576 = a4 & ~n314;
  assign n577 = n293 & n576;
  assign n578 = ~n300 & n577;
  assign n579 = ~n537 & n576;
  assign n580 = n293 & n579;
  assign n581 = a4 & n293;
  assign n582 = n318 & n581;
  assign n583 = ~n404 & ~n435;
  assign n584 = ~n582 & n583;
  assign n585 = ~n580 & n584;
  assign n586 = ~n578 & n585;
  assign j9 = n575 | ~n586;
  assign n588 = b2 & ~n305;
  assign n589 = n299 & n588;
  assign n590 = c2 & n305;
  assign n591 = n299 & n590;
  assign n592 = u & n306;
  assign n593 = ~n591 & ~n592;
  assign k7 = n589 | ~n593;
  assign n595 = c3 & n356;
  assign n596 = b3 & ~n360;
  assign k8 = n595 | n596;
  assign n598 = b4 & i9;
  assign n599 = n299 & n598;
  assign n600 = b4 & ~i9;
  assign n601 = ~n572 & n600;
  assign n602 = n302 & ~i9;
  assign n603 = ~n435 & ~n602;
  assign n604 = ~n601 & n603;
  assign k9 = n599 | ~n604;
  assign l5 = g1 & ~j4;
  assign n607 = c2 & ~n305;
  assign n608 = n299 & n607;
  assign n609 = d2 & n305;
  assign n610 = n299 & n609;
  assign n611 = v & n306;
  assign n612 = ~n610 & ~n611;
  assign l7 = n608 | ~n612;
  assign n614 = d3 & n356;
  assign n615 = c3 & ~n360;
  assign l8 = n614 | n615;
  assign n617 = c4 & i9;
  assign n618 = ~n435 & n617;
  assign n619 = n293 & n618;
  assign n620 = c4 & ~i9;
  assign n621 = ~n572 & n620;
  assign n622 = b4 & c4;
  assign n623 = ~i9 & n622;
  assign n624 = n293 & n314;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n621 & n625;
  assign l9 = n619 | ~n626;
  assign n628 = d2 & ~n305;
  assign n629 = n299 & n628;
  assign n630 = e2 & n305;
  assign n631 = n299 & n630;
  assign n632 = w & n306;
  assign n633 = ~n631 & ~n632;
  assign m7 = n629 | ~n633;
  assign n635 = e3 & n356;
  assign n636 = d3 & ~n360;
  assign m8 = n635 | n636;
  assign n638 = ~d4 & ~n335;
  assign n639 = ~g1 & n293;
  assign n640 = ~g1 & w9;
  assign n641 = n638 & n640;
  assign n642 = d4 & n639;
  assign n643 = ~n357 & n642;
  assign n644 = d4 & n335;
  assign n645 = n639 & n644;
  assign n646 = ~n306 & ~n645;
  assign n647 = ~n643 & n646;
  assign m9 = n641 | ~n647;
  assign n649 = ~k4 & ~n0;
  assign n5 = ~h1 | ~n649;
  assign n651 = ~f1 & ~i4;
  assign n652 = f1 & i4;
  assign n6 = n651 | n652;
  assign n654 = e2 & ~n305;
  assign n655 = n299 & n654;
  assign n656 = f2 & n305;
  assign n657 = n299 & n656;
  assign n658 = x & n306;
  assign n659 = ~n657 & ~n658;
  assign n7 = n655 | ~n659;
  assign n661 = f3 & n356;
  assign n662 = e3 & ~n360;
  assign n8 = n661 | n662;
  assign n664 = n638 & m9;
  assign n665 = ~n298 & n639;
  assign n666 = ~e4 & n664;
  assign n667 = e4 & ~n664;
  assign n668 = n665 & ~n667;
  assign n9 = n666 | ~n668;
  assign o5 = ~i1 | ~n649;
  assign o6 = x3 & n303;
  assign n672 = f2 & ~n305;
  assign n673 = n299 & n672;
  assign n674 = g2 & n305;
  assign n675 = n299 & n674;
  assign n676 = y & n306;
  assign n677 = ~n675 & ~n676;
  assign o7 = n673 | ~n677;
  assign n679 = g3 & n356;
  assign n680 = f3 & ~n360;
  assign o8 = n679 | n680;
  assign n682 = e4 & ~n9;
  assign n683 = ~f4 & n682;
  assign n684 = f4 & ~n682;
  assign n685 = n665 & ~n684;
  assign o9 = n683 | ~n685;
  assign n687 = m0 & ~n285;
  assign n688 = l3 & n687;
  assign n689 = t3 & ~k5;
  assign n690 = d3 & n286;
  assign n691 = ~n689 & ~n690;
  assign p4 = n688 | ~n691;
  assign p5 = ~j1 | ~n649;
  assign n694 = n4 & ~n335;
  assign n695 = n293 & n353;
  assign n696 = n694 & n695;
  assign p6 = n645 | n696;
  assign n698 = g2 & ~n305;
  assign n699 = n299 & n698;
  assign n700 = h2 & n305;
  assign n701 = n299 & n700;
  assign n702 = z & n306;
  assign n703 = ~n701 & ~n702;
  assign p7 = n699 | ~n703;
  assign n705 = h3 & n356;
  assign n706 = g3 & ~n360;
  assign p8 = n705 | n706;
  assign n708 = g4 & o9;
  assign n709 = n665 & n708;
  assign n710 = ~f4 & g4;
  assign n711 = n665 & n710;
  assign n712 = n285 & m9;
  assign n713 = ~n665 & n712;
  assign n714 = n333 & ~o9;
  assign n715 = n314 & m9;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n713 & n716;
  assign n718 = ~n711 & n717;
  assign p9 = n709 | ~n718;
  assign n720 = k3 & n687;
  assign n721 = s3 & ~j5;
  assign n722 = c3 & n286;
  assign n723 = ~n721 & ~n722;
  assign q4 = n720 | ~n723;
  assign q5 = ~k1 | ~n649;
  assign n726 = ~e1 & n298;
  assign n727 = n293 & n726;
  assign n728 = ~c1 & ~d1;
  assign n729 = h1 & n639;
  assign n730 = n727 & n728;
  assign q6 = n729 | n730;
  assign n732 = h2 & ~n305;
  assign n733 = n299 & n732;
  assign n734 = i2 & n305;
  assign n735 = n299 & n734;
  assign n736 = a0 & n306;
  assign n737 = ~n735 & ~n736;
  assign q7 = n733 | ~n737;
  assign n739 = i3 & n356;
  assign n740 = h3 & ~n360;
  assign q8 = n739 | n740;
  assign n742 = h4 & ~n334;
  assign n743 = n665 & n742;
  assign n744 = h4 & ~w9;
  assign n745 = n665 & n744;
  assign n746 = h4 & ~m9;
  assign n747 = n665 & n746;
  assign n748 = ~n435 & ~n747;
  assign n749 = ~n745 & n748;
  assign q9 = n743 | ~n749;
  assign n751 = j3 & n687;
  assign n752 = r3 & ~i5;
  assign n753 = b3 & n286;
  assign n754 = ~n752 & ~n753;
  assign r4 = n751 | ~n754;
  assign r5 = ~l1 | ~n649;
  assign n757 = c1 & ~d1;
  assign n758 = n727 & n757;
  assign n759 = i1 & n639;
  assign r6 = n758 | n759;
  assign n761 = i2 & ~n305;
  assign n762 = n299 & n761;
  assign n763 = j2 & n305;
  assign n764 = n299 & n763;
  assign n765 = b0 & n306;
  assign n766 = ~n764 & ~n765;
  assign r7 = n762 | ~n766;
  assign n768 = j3 & n356;
  assign n769 = i3 & ~n360;
  assign r8 = n768 | n769;
  assign n771 = ~i4 & n1;
  assign n772 = n305 & n771;
  assign n773 = n293 & n772;
  assign n774 = i4 & ~n1;
  assign n775 = n305 & n774;
  assign n776 = n293 & n775;
  assign r9 = n773 | n776;
  assign n778 = i3 & n687;
  assign n779 = q3 & ~h5;
  assign n780 = a3 & n286;
  assign n781 = ~n779 & ~n780;
  assign s4 = n778 | ~n781;
  assign n783 = n303 & n6;
  assign n784 = n1 & ~n303;
  assign s5 = n783 | n784;
  assign n786 = j1 & n639;
  assign n787 = ~c1 & d1;
  assign n788 = n727 & n787;
  assign s6 = n786 | n788;
  assign n790 = j2 & ~n305;
  assign n791 = n299 & n790;
  assign n792 = k2 & n305;
  assign n793 = n299 & n792;
  assign n794 = c0 & n306;
  assign n795 = ~n793 & ~n794;
  assign s7 = n791 | ~n795;
  assign n797 = k3 & n356;
  assign n798 = j3 & ~n360;
  assign s8 = n797 | n798;
  assign n800 = ~j4 & n500;
  assign n801 = n356 & n800;
  assign n802 = n639 & n801;
  assign n803 = n694 & n802;
  assign n804 = j4 & ~n356;
  assign n805 = n639 & n804;
  assign n806 = j4 & ~n500;
  assign n807 = n639 & n806;
  assign n808 = j4 & ~n4;
  assign n809 = n639 & n808;
  assign n810 = ~n807 & ~n809;
  assign n811 = ~n805 & n810;
  assign s9 = n803 | ~n811;
  assign n813 = k1 & n639;
  assign n814 = c1 & d1;
  assign n815 = n727 & n814;
  assign t6 = n813 | n815;
  assign n817 = i & n293;
  assign n818 = n316 & n817;
  assign n819 = l2 & n293;
  assign n820 = n317 & n819;
  assign n821 = k2 & n293;
  assign n822 = n318 & n821;
  assign n823 = a & n293;
  assign n824 = ~n321 & n823;
  assign n825 = ~n822 & ~n824;
  assign n826 = ~n820 & n825;
  assign t7 = n818 | ~n826;
  assign n828 = l3 & n356;
  assign n829 = k3 & ~n360;
  assign t8 = n828 | n829;
  assign n831 = m1 & n293;
  assign t9 = n303 & n831;
  assign n833 = ~n726 & n728;
  assign n834 = n306 & n833;
  assign n835 = l1 & n639;
  assign u6 = n834 | n835;
  assign n837 = j & n293;
  assign n838 = n316 & n837;
  assign n839 = m2 & n293;
  assign n840 = n317 & n839;
  assign n841 = n318 & n819;
  assign n842 = b & n293;
  assign n843 = ~n321 & n842;
  assign n844 = ~n841 & ~n843;
  assign n845 = ~n840 & n844;
  assign u7 = n838 | ~n845;
  assign n847 = m3 & n356;
  assign n848 = l3 & ~n360;
  assign u8 = n847 | n848;
  assign u9 = ~n304 & n831;
  assign n851 = e3 & n286;
  assign n852 = ~n285 & d5;
  assign v4 = n851 | n852;
  assign n854 = ~p6 & n831;
  assign n855 = ~n0 & p0;
  assign n856 = ~m1 & n855;
  assign n857 = n293 & n856;
  assign v6 = n854 | n857;
  assign n859 = k & n293;
  assign n860 = n316 & n859;
  assign n861 = n2 & n293;
  assign n862 = n317 & n861;
  assign n863 = n318 & n839;
  assign n864 = c & n293;
  assign n865 = ~n321 & n864;
  assign n866 = ~n863 & ~n865;
  assign n867 = ~n862 & n866;
  assign v7 = n860 | ~n867;
  assign n869 = n3 & n356;
  assign n870 = m3 & ~n360;
  assign v8 = n869 | n870;
  assign n872 = n694 & p6;
  assign n873 = ~n353 & p6;
  assign v9 = n872 | n873;
  assign n875 = f3 & n286;
  assign n876 = ~n285 & e5;
  assign w4 = n875 | n876;
  assign n878 = n1 & ~n305;
  assign n879 = n299 & n878;
  assign n880 = o1 & n305;
  assign n881 = n299 & n880;
  assign n882 = j0 & n306;
  assign n883 = ~n881 & ~n882;
  assign w6 = n879 | ~n883;
  assign n885 = l & n293;
  assign n886 = n316 & n885;
  assign n887 = o2 & n293;
  assign n888 = n317 & n887;
  assign n889 = n318 & n861;
  assign n890 = d & n293;
  assign n891 = ~n321 & n890;
  assign n892 = ~n889 & ~n891;
  assign n893 = ~n888 & n892;
  assign w7 = n886 | ~n893;
  assign n895 = o3 & n356;
  assign n896 = n3 & ~n360;
  assign w8 = n895 | n896;
  assign n898 = g3 & n286;
  assign n899 = ~n285 & f5;
  assign x4 = n898 | n899;
  assign x5 = ~h1 | ~n291;
  assign n902 = o1 & ~n305;
  assign n903 = n299 & n902;
  assign n904 = p1 & n305;
  assign n905 = n299 & n904;
  assign n906 = i0 & n306;
  assign n907 = ~n905 & ~n906;
  assign x6 = n903 | ~n907;
  assign n909 = m & n293;
  assign n910 = n316 & n909;
  assign n911 = p2 & n293;
  assign n912 = n317 & n911;
  assign n913 = n318 & n887;
  assign n914 = e & n293;
  assign n915 = ~n321 & n914;
  assign n916 = ~n913 & ~n915;
  assign n917 = ~n912 & n916;
  assign x7 = n910 | ~n917;
  assign n919 = p3 & n356;
  assign n920 = o3 & ~n360;
  assign x8 = n919 | n920;
  assign n922 = h3 & n286;
  assign n923 = ~n285 & g5;
  assign y4 = n922 | n923;
  assign y5 = ~i1 | ~n291;
  assign n926 = p1 & ~n305;
  assign n927 = n299 & n926;
  assign n928 = q1 & n305;
  assign n929 = n299 & n928;
  assign n930 = h0 & n306;
  assign n931 = ~n929 & ~n930;
  assign y6 = n927 | ~n931;
  assign n933 = n & n293;
  assign n934 = n316 & n933;
  assign n935 = n317 & n326;
  assign n936 = n318 & n911;
  assign n937 = f & n293;
  assign n938 = ~n321 & n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~n935 & n939;
  assign y7 = n934 | ~n940;
  assign n942 = q3 & n356;
  assign n943 = p3 & ~n360;
  assign y8 = n942 | n943;
  assign h6 = ~h1;
  assign i6 = ~i1;
  assign j6 = ~j1;
  assign k6 = ~k1;
  assign l6 = ~l1;
  assign o4 = ~g1;
  assign m5 = m4;
  assign m6 = k4;
  assign t4 = u3;
  assign t5 = s5;
  assign u4 = v3;
  assign u5 = s5;
  assign v5 = s5;
  assign w5 = s5;
endmodule


